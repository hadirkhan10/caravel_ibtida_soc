magic
tech sky130A
magscale 1 2
timestamp 1607603059
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 412649 683247 412683 692733
rect 218989 666587 219023 676141
rect 413017 666587 413051 683077
rect 429577 666587 429611 683077
rect 542737 666587 542771 683077
rect 559297 666587 559331 683077
rect 72985 647275 73019 656829
rect 219265 647275 219299 656829
rect 72801 627963 72835 637517
rect 219081 627963 219115 637517
rect 395813 87023 395847 96577
rect 152841 77299 152875 86921
rect 410993 77367 411027 82093
rect 148885 67643 148919 77197
rect 188537 67643 188571 77197
rect 225889 67643 225923 77197
rect 235641 67643 235675 77197
rect 297741 67643 297775 77197
rect 378149 67711 378183 77197
rect 235825 45611 235859 50405
rect 353309 48331 353343 57885
rect 371249 56627 371283 66181
rect 378149 57987 378183 67541
rect 499589 57987 499623 67541
rect 378149 48331 378183 57817
rect 410717 50983 410751 56525
rect 495449 48331 495483 57885
rect 333805 47583 333839 48161
rect 235733 29631 235767 41429
rect 371249 37315 371283 46869
rect 378149 29087 378183 38573
rect 369869 9707 369903 19261
rect 371249 18003 371283 27557
rect 410901 26299 410935 35853
rect 495449 29019 495483 38573
rect 378149 9707 378183 19261
rect 397469 9707 397503 19261
rect 410901 8415 410935 22117
rect 415409 9707 415443 19261
rect 561689 9707 561723 19261
rect 410901 6171 410935 8245
rect 356069 4879 356103 4981
rect 365637 4811 365671 4981
rect 365729 4879 365763 4981
rect 370513 4879 370547 4981
rect 376803 4777 376861 4811
rect 496553 595 496587 9605
rect 547889 3655 547923 3757
rect 500083 3621 500325 3655
rect 558193 3655 558227 3757
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 412649 692733 412683 692767
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 412649 683213 412683 683247
rect 284033 676209 284067 676243
rect 413017 683077 413051 683111
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 413017 666553 413051 666587
rect 429577 683077 429611 683111
rect 429577 666553 429611 666587
rect 542737 683077 542771 683111
rect 542737 666553 542771 666587
rect 559297 683077 559331 683111
rect 559297 666553 559331 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 72801 637517 72835 637551
rect 72801 627929 72835 627963
rect 219081 637517 219115 637551
rect 219081 627929 219115 627963
rect 395813 96577 395847 96611
rect 395813 86989 395847 87023
rect 152841 86921 152875 86955
rect 410993 82093 411027 82127
rect 410993 77333 411027 77367
rect 152841 77265 152875 77299
rect 148885 77197 148919 77231
rect 148885 67609 148919 67643
rect 188537 77197 188571 77231
rect 188537 67609 188571 67643
rect 225889 77197 225923 77231
rect 225889 67609 225923 67643
rect 235641 77197 235675 77231
rect 235641 67609 235675 67643
rect 297741 77197 297775 77231
rect 378149 77197 378183 77231
rect 378149 67677 378183 67711
rect 297741 67609 297775 67643
rect 378149 67541 378183 67575
rect 371249 66181 371283 66215
rect 353309 57885 353343 57919
rect 235825 50405 235859 50439
rect 378149 57953 378183 57987
rect 499589 67541 499623 67575
rect 499589 57953 499623 57987
rect 495449 57885 495483 57919
rect 371249 56593 371283 56627
rect 378149 57817 378183 57851
rect 353309 48297 353343 48331
rect 410717 56525 410751 56559
rect 410717 50949 410751 50983
rect 378149 48297 378183 48331
rect 495449 48297 495483 48331
rect 333805 48161 333839 48195
rect 333805 47549 333839 47583
rect 235825 45577 235859 45611
rect 371249 46869 371283 46903
rect 235733 41429 235767 41463
rect 371249 37281 371283 37315
rect 378149 38573 378183 38607
rect 235733 29597 235767 29631
rect 495449 38573 495483 38607
rect 378149 29053 378183 29087
rect 410901 35853 410935 35887
rect 371249 27557 371283 27591
rect 369869 19261 369903 19295
rect 495449 28985 495483 29019
rect 410901 26265 410935 26299
rect 410901 22117 410935 22151
rect 371249 17969 371283 18003
rect 378149 19261 378183 19295
rect 369869 9673 369903 9707
rect 378149 9673 378183 9707
rect 397469 19261 397503 19295
rect 397469 9673 397503 9707
rect 415409 19261 415443 19295
rect 415409 9673 415443 9707
rect 561689 19261 561723 19295
rect 561689 9673 561723 9707
rect 410901 8381 410935 8415
rect 496553 9605 496587 9639
rect 410901 8245 410935 8279
rect 410901 6137 410935 6171
rect 356069 4981 356103 5015
rect 356069 4845 356103 4879
rect 365637 4981 365671 5015
rect 365729 4981 365763 5015
rect 365729 4845 365763 4879
rect 370513 4981 370547 5015
rect 370513 4845 370547 4879
rect 365637 4777 365671 4811
rect 376769 4777 376803 4811
rect 376861 4777 376895 4811
rect 547889 3757 547923 3791
rect 500049 3621 500083 3655
rect 500325 3621 500359 3655
rect 547889 3621 547923 3655
rect 558193 3757 558227 3791
rect 558193 3621 558227 3655
rect 496553 561 496587 595
<< metal1 >>
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 331214 697552 331220 697604
rect 331272 697592 331278 697604
rect 332502 697592 332508 697604
rect 331272 697564 332508 697592
rect 331272 697552 331278 697564
rect 332502 697552 332508 697564
rect 332560 697552 332566 697604
rect 538858 696940 538864 696992
rect 538916 696980 538922 696992
rect 580166 696980 580172 696992
rect 538916 696952 580172 696980
rect 538916 696940 538922 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 347774 692792 347780 692844
rect 347832 692832 347838 692844
rect 348878 692832 348884 692844
rect 347832 692804 348884 692832
rect 347832 692792 347838 692804
rect 348878 692792 348884 692804
rect 348936 692792 348942 692844
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 542538 692724 542544 692776
rect 542596 692764 542602 692776
rect 542722 692764 542728 692776
rect 542596 692736 542728 692764
rect 542596 692724 542602 692736
rect 542722 692724 542728 692736
rect 542780 692724 542786 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 429194 684428 429200 684480
rect 429252 684468 429258 684480
rect 429838 684468 429844 684480
rect 429252 684440 429844 684468
rect 429252 684428 429258 684440
rect 429838 684428 429844 684440
rect 429896 684428 429902 684480
rect 558914 684428 558920 684480
rect 558972 684468 558978 684480
rect 559650 684468 559656 684480
rect 558972 684440 559656 684468
rect 558972 684428 558978 684440
rect 559650 684428 559656 684440
rect 559708 684428 559714 684480
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 429194 683068 429200 683120
rect 429252 683108 429258 683120
rect 429565 683111 429623 683117
rect 429565 683108 429577 683111
rect 429252 683080 429577 683108
rect 429252 683068 429258 683080
rect 429565 683077 429577 683080
rect 429611 683077 429623 683111
rect 429565 683071 429623 683077
rect 542354 683068 542360 683120
rect 542412 683108 542418 683120
rect 542725 683111 542783 683117
rect 542725 683108 542737 683111
rect 542412 683080 542737 683108
rect 542412 683068 542418 683080
rect 542725 683077 542737 683080
rect 542771 683077 542783 683111
rect 542725 683071 542783 683077
rect 558914 683068 558920 683120
rect 558972 683108 558978 683120
rect 559285 683111 559343 683117
rect 559285 683108 559297 683111
rect 558972 683080 559297 683108
rect 558972 683068 558978 683080
rect 559285 683077 559297 683080
rect 559331 683077 559343 683111
rect 559285 683071 559343 683077
rect 3786 681708 3792 681760
rect 3844 681748 3850 681760
rect 32398 681748 32404 681760
rect 3844 681720 32404 681748
rect 3844 681708 3850 681720
rect 32398 681708 32404 681720
rect 32456 681708 32462 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 347774 673480 347780 673532
rect 347832 673520 347838 673532
rect 347958 673520 347964 673532
rect 347832 673492 347964 673520
rect 347832 673480 347838 673492
rect 347958 673480 347964 673492
rect 348016 673480 348022 673532
rect 364334 673480 364340 673532
rect 364392 673520 364398 673532
rect 364518 673520 364524 673532
rect 364392 673492 364524 673520
rect 364392 673480 364398 673492
rect 364518 673480 364524 673492
rect 364576 673480 364582 673532
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 494054 673480 494060 673532
rect 494112 673520 494118 673532
rect 494238 673520 494244 673532
rect 494112 673492 494244 673520
rect 494112 673480 494118 673492
rect 494238 673480 494244 673492
rect 494296 673480 494302 673532
rect 536098 673480 536104 673532
rect 536156 673520 536162 673532
rect 580166 673520 580172 673532
rect 536156 673492 580172 673520
rect 536156 673480 536162 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 284018 654100 284024 654152
rect 284076 654140 284082 654152
rect 284202 654140 284208 654152
rect 284076 654112 284208 654140
rect 284076 654100 284082 654112
rect 284202 654100 284208 654112
rect 284260 654100 284266 654152
rect 347774 654100 347780 654152
rect 347832 654140 347838 654152
rect 347958 654140 347964 654152
rect 347832 654112 347964 654140
rect 347832 654100 347838 654112
rect 347958 654100 347964 654112
rect 348016 654100 348022 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 10318 652780 10324 652792
rect 3108 652752 10324 652780
rect 3108 652740 3114 652752
rect 10318 652740 10324 652752
rect 10376 652740 10382 652792
rect 529198 650020 529204 650072
rect 529256 650060 529262 650072
rect 580166 650060 580172 650072
rect 529256 650032 580172 650060
rect 529256 650020 529262 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 72786 637548 72792 637560
rect 72747 637520 72792 637548
rect 72786 637508 72792 637520
rect 72844 637508 72850 637560
rect 219066 637548 219072 637560
rect 219027 637520 219072 637548
rect 219066 637508 219072 637520
rect 219124 637508 219130 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 284018 634788 284024 634840
rect 284076 634828 284082 634840
rect 284202 634828 284208 634840
rect 284076 634800 284208 634828
rect 284076 634788 284082 634800
rect 284202 634788 284208 634800
rect 284260 634788 284266 634840
rect 347774 634788 347780 634840
rect 347832 634828 347838 634840
rect 347958 634828 347964 634840
rect 347832 634800 347964 634828
rect 347832 634788 347838 634800
rect 347958 634788 347964 634800
rect 348016 634788 348022 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 72789 627963 72847 627969
rect 72789 627929 72801 627963
rect 72835 627960 72847 627963
rect 73062 627960 73068 627972
rect 72835 627932 73068 627960
rect 72835 627929 72847 627932
rect 72789 627923 72847 627929
rect 73062 627920 73068 627932
rect 73120 627920 73126 627972
rect 219069 627963 219127 627969
rect 219069 627929 219081 627963
rect 219115 627960 219127 627963
rect 219342 627960 219348 627972
rect 219115 627932 219348 627960
rect 219115 627929 219127 627932
rect 219069 627923 219127 627929
rect 219342 627920 219348 627932
rect 219400 627920 219406 627972
rect 571978 626560 571984 626612
rect 572036 626600 572042 626612
rect 580166 626600 580172 626612
rect 572036 626572 580172 626600
rect 572036 626560 572042 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 8938 623812 8944 623824
rect 3292 623784 8944 623812
rect 3292 623772 3298 623784
rect 8938 623772 8944 623784
rect 8996 623772 9002 623824
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 284018 615476 284024 615528
rect 284076 615516 284082 615528
rect 284202 615516 284208 615528
rect 284076 615488 284208 615516
rect 284076 615476 284082 615488
rect 284202 615476 284208 615488
rect 284260 615476 284266 615528
rect 347774 615476 347780 615528
rect 347832 615516 347838 615528
rect 347958 615516 347964 615528
rect 347832 615488 347964 615516
rect 347832 615476 347838 615488
rect 347958 615476 347964 615488
rect 348016 615476 348022 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 477494 615476 477500 615528
rect 477552 615516 477558 615528
rect 477678 615516 477684 615528
rect 477552 615488 477684 615516
rect 477552 615476 477558 615488
rect 477678 615476 477684 615488
rect 477736 615476 477742 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 300762 604392 300768 604444
rect 300820 604432 300826 604444
rect 307478 604432 307484 604444
rect 300820 604404 307484 604432
rect 300820 604392 300826 604404
rect 307478 604392 307484 604404
rect 307536 604392 307542 604444
rect 89622 603984 89628 604036
rect 89680 604024 89686 604036
rect 151906 604024 151912 604036
rect 89680 603996 151912 604024
rect 89680 603984 89686 603996
rect 151906 603984 151912 603996
rect 151964 603984 151970 604036
rect 73062 603916 73068 603968
rect 73120 603956 73126 603968
rect 136358 603956 136364 603968
rect 73120 603928 136364 603956
rect 73120 603916 73126 603928
rect 136358 603916 136364 603928
rect 136416 603916 136422 603968
rect 41322 603848 41328 603900
rect 41380 603888 41386 603900
rect 120810 603888 120816 603900
rect 41380 603860 120816 603888
rect 41380 603848 41386 603860
rect 120810 603848 120816 603860
rect 120868 603848 120874 603900
rect 154298 603848 154304 603900
rect 154356 603888 154362 603900
rect 198550 603888 198556 603900
rect 154356 603860 198556 603888
rect 154356 603848 154362 603860
rect 198550 603848 198556 603860
rect 198608 603848 198614 603900
rect 385218 603848 385224 603900
rect 385276 603888 385282 603900
rect 412726 603888 412732 603900
rect 385276 603860 412732 603888
rect 385276 603848 385282 603860
rect 412726 603848 412732 603860
rect 412784 603848 412790 603900
rect 447410 603848 447416 603900
rect 447468 603888 447474 603900
rect 494238 603888 494244 603900
rect 447468 603860 494244 603888
rect 447468 603848 447474 603860
rect 494238 603848 494244 603860
rect 494296 603848 494302 603900
rect 494330 603848 494336 603900
rect 494388 603888 494394 603900
rect 559006 603888 559012 603900
rect 494388 603860 559012 603888
rect 494388 603848 494394 603860
rect 559006 603848 559012 603860
rect 559064 603848 559070 603900
rect 24762 603780 24768 603832
rect 24820 603820 24826 603832
rect 105262 603820 105268 603832
rect 24820 603792 105268 603820
rect 24820 603780 24826 603792
rect 105262 603780 105268 603792
rect 105320 603780 105326 603832
rect 137738 603780 137744 603832
rect 137796 603820 137802 603832
rect 183002 603820 183008 603832
rect 137796 603792 183008 603820
rect 137796 603780 137802 603792
rect 183002 603780 183008 603792
rect 183060 603780 183066 603832
rect 202782 603780 202788 603832
rect 202840 603820 202846 603832
rect 229646 603820 229652 603832
rect 202840 603792 229652 603820
rect 202840 603780 202846 603792
rect 229646 603780 229652 603792
rect 229704 603780 229710 603832
rect 235902 603780 235908 603832
rect 235960 603820 235966 603832
rect 260742 603820 260748 603832
rect 235960 603792 260748 603820
rect 235960 603780 235966 603792
rect 260742 603780 260748 603792
rect 260800 603780 260806 603832
rect 400766 603780 400772 603832
rect 400824 603820 400830 603832
rect 429286 603820 429292 603832
rect 400824 603792 429292 603820
rect 400824 603780 400830 603792
rect 429286 603780 429292 603792
rect 429344 603780 429350 603832
rect 431862 603780 431868 603832
rect 431920 603820 431926 603832
rect 477678 603820 477684 603832
rect 431920 603792 477684 603820
rect 431920 603780 431926 603792
rect 477678 603780 477684 603792
rect 477736 603780 477742 603832
rect 478506 603780 478512 603832
rect 478564 603820 478570 603832
rect 542446 603820 542452 603832
rect 478564 603792 542452 603820
rect 478564 603780 478570 603792
rect 542446 603780 542452 603792
rect 542504 603780 542510 603832
rect 8018 603712 8024 603764
rect 8076 603752 8082 603764
rect 89714 603752 89720 603764
rect 8076 603724 89720 603752
rect 8076 603712 8082 603724
rect 89714 603712 89720 603724
rect 89772 603712 89778 603764
rect 106182 603712 106188 603764
rect 106240 603752 106246 603764
rect 167454 603752 167460 603764
rect 106240 603724 167460 603752
rect 106240 603712 106246 603724
rect 167454 603712 167460 603724
rect 167512 603712 167518 603764
rect 171042 603712 171048 603764
rect 171100 603752 171106 603764
rect 214098 603752 214104 603764
rect 171100 603724 214104 603752
rect 171100 603712 171106 603724
rect 214098 603712 214104 603724
rect 214156 603712 214162 603764
rect 219342 603712 219348 603764
rect 219400 603752 219406 603764
rect 245194 603752 245200 603764
rect 219400 603724 245200 603752
rect 219400 603712 219406 603724
rect 245194 603712 245200 603724
rect 245252 603712 245258 603764
rect 267642 603712 267648 603764
rect 267700 603752 267706 603764
rect 276290 603752 276296 603764
rect 267700 603724 276296 603752
rect 267700 603712 267706 603724
rect 276290 603712 276296 603724
rect 276348 603712 276354 603764
rect 284018 603712 284024 603764
rect 284076 603752 284082 603764
rect 291838 603752 291844 603764
rect 284076 603724 291844 603752
rect 284076 603712 284082 603724
rect 291838 603712 291844 603724
rect 291896 603712 291902 603764
rect 323026 603712 323032 603764
rect 323084 603752 323090 603764
rect 331214 603752 331220 603764
rect 323084 603724 331220 603752
rect 323084 603712 323090 603724
rect 331214 603712 331220 603724
rect 331272 603712 331278 603764
rect 338574 603712 338580 603764
rect 338632 603752 338638 603764
rect 347958 603752 347964 603764
rect 338632 603724 347964 603752
rect 338632 603712 338638 603724
rect 347958 603712 347964 603724
rect 348016 603712 348022 603764
rect 354122 603712 354128 603764
rect 354180 603752 354186 603764
rect 364518 603752 364524 603764
rect 354180 603724 364524 603752
rect 354180 603712 354186 603724
rect 364518 603712 364524 603724
rect 364576 603712 364582 603764
rect 369670 603712 369676 603764
rect 369728 603752 369734 603764
rect 397454 603752 397460 603764
rect 369728 603724 397460 603752
rect 369728 603712 369734 603724
rect 397454 603712 397460 603724
rect 397512 603712 397518 603764
rect 416314 603712 416320 603764
rect 416372 603752 416378 603764
rect 462314 603752 462320 603764
rect 416372 603724 462320 603752
rect 416372 603712 416378 603724
rect 462314 603712 462320 603724
rect 462372 603712 462378 603764
rect 462958 603712 462964 603764
rect 463016 603752 463022 603764
rect 527174 603752 527180 603764
rect 463016 603724 527180 603752
rect 463016 603712 463022 603724
rect 527174 603712 527180 603724
rect 527232 603712 527238 603764
rect 565078 603100 565084 603152
rect 565136 603140 565142 603152
rect 580166 603140 580172 603152
rect 565136 603112 580172 603140
rect 565136 603100 565142 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 505002 597456 505008 597508
rect 505060 597496 505066 597508
rect 538858 597496 538864 597508
rect 505060 597468 538864 597496
rect 505060 597456 505066 597468
rect 538858 597456 538864 597468
rect 538916 597456 538922 597508
rect 32398 596096 32404 596148
rect 32456 596136 32462 596148
rect 78674 596136 78680 596148
rect 32456 596108 78680 596136
rect 32456 596096 32462 596108
rect 78674 596096 78680 596108
rect 78732 596096 78738 596148
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 13078 594844 13084 594856
rect 3384 594816 13084 594844
rect 3384 594804 3390 594816
rect 13078 594804 13084 594816
rect 13136 594804 13142 594856
rect 507118 592016 507124 592068
rect 507176 592056 507182 592068
rect 579890 592056 579896 592068
rect 507176 592028 579896 592056
rect 507176 592016 507182 592028
rect 579890 592016 579896 592028
rect 579948 592016 579954 592068
rect 504634 586440 504640 586492
rect 504692 586480 504698 586492
rect 580258 586480 580264 586492
rect 504692 586452 580264 586480
rect 504692 586440 504698 586452
rect 580258 586440 580264 586452
rect 580316 586440 580322 586492
rect 3418 585080 3424 585132
rect 3476 585120 3482 585132
rect 78674 585120 78680 585132
rect 3476 585092 78680 585120
rect 3476 585080 3482 585092
rect 78674 585080 78680 585092
rect 78732 585080 78738 585132
rect 511258 579640 511264 579692
rect 511316 579680 511322 579692
rect 580166 579680 580172 579692
rect 511316 579652 580172 579680
rect 511316 579640 511322 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 505002 573996 505008 574048
rect 505060 574036 505066 574048
rect 536098 574036 536104 574048
rect 505060 574008 536104 574036
rect 505060 573996 505066 574008
rect 536098 573996 536104 574008
rect 536156 573996 536162 574048
rect 10318 572636 10324 572688
rect 10376 572676 10382 572688
rect 78674 572676 78680 572688
rect 10376 572648 78680 572676
rect 10376 572636 10382 572648
rect 78674 572636 78680 572648
rect 78732 572636 78738 572688
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 10318 567236 10324 567248
rect 3476 567208 10324 567236
rect 3476 567196 3482 567208
rect 10318 567196 10324 567208
rect 10376 567196 10382 567248
rect 505002 562980 505008 563032
rect 505060 563020 505066 563032
rect 529198 563020 529204 563032
rect 505060 562992 529204 563020
rect 505060 562980 505066 562992
rect 529198 562980 529204 562992
rect 529256 562980 529262 563032
rect 8938 560192 8944 560244
rect 8996 560232 9002 560244
rect 78674 560232 78680 560244
rect 8996 560204 78680 560232
rect 8996 560192 9002 560204
rect 78674 560192 78680 560204
rect 78732 560192 78738 560244
rect 504358 556180 504364 556232
rect 504416 556220 504422 556232
rect 580166 556220 580172 556232
rect 504416 556192 580172 556220
rect 504416 556180 504422 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 505002 551964 505008 552016
rect 505060 552004 505066 552016
rect 580350 552004 580356 552016
rect 505060 551976 580356 552004
rect 505060 551964 505066 551976
rect 580350 551964 580356 551976
rect 580408 551964 580414 552016
rect 3510 549176 3516 549228
rect 3568 549216 3574 549228
rect 78674 549216 78680 549228
rect 3568 549188 78680 549216
rect 3568 549176 3574 549188
rect 78674 549176 78680 549188
rect 78732 549176 78738 549228
rect 505002 540880 505008 540932
rect 505060 540920 505066 540932
rect 571978 540920 571984 540932
rect 505060 540892 571984 540920
rect 505060 540880 505066 540892
rect 571978 540880 571984 540892
rect 572036 540880 572042 540932
rect 13078 536732 13084 536784
rect 13136 536772 13142 536784
rect 78674 536772 78680 536784
rect 13136 536744 78680 536772
rect 13136 536732 13142 536744
rect 78674 536732 78680 536744
rect 78732 536732 78738 536784
rect 505738 532720 505744 532772
rect 505796 532760 505802 532772
rect 580166 532760 580172 532772
rect 505796 532732 580172 532760
rect 505796 532720 505802 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 505002 529864 505008 529916
rect 505060 529904 505066 529916
rect 565078 529904 565084 529916
rect 505060 529876 565084 529904
rect 505060 529864 505066 529876
rect 565078 529864 565084 529876
rect 565136 529864 565142 529916
rect 10318 525716 10324 525768
rect 10376 525756 10382 525768
rect 78674 525756 78680 525768
rect 10376 525728 78680 525756
rect 10376 525716 10382 525728
rect 78674 525716 78680 525728
rect 78732 525716 78738 525768
rect 504174 518508 504180 518560
rect 504232 518548 504238 518560
rect 507118 518548 507124 518560
rect 504232 518520 507124 518548
rect 504232 518508 504238 518520
rect 507118 518508 507124 518520
rect 507176 518508 507182 518560
rect 3418 513272 3424 513324
rect 3476 513312 3482 513324
rect 78674 513312 78680 513324
rect 3476 513284 78680 513312
rect 3476 513272 3482 513284
rect 78674 513272 78680 513284
rect 78732 513272 78738 513324
rect 507118 509260 507124 509312
rect 507176 509300 507182 509312
rect 580166 509300 580172 509312
rect 507176 509272 580172 509300
rect 507176 509260 507182 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 505002 507696 505008 507748
rect 505060 507736 505066 507748
rect 511258 507736 511264 507748
rect 505060 507708 511264 507736
rect 505060 507696 505066 507708
rect 511258 507696 511264 507708
rect 511316 507696 511322 507748
rect 3510 500896 3516 500948
rect 3568 500936 3574 500948
rect 78674 500936 78680 500948
rect 3568 500908 78680 500936
rect 3568 500896 3574 500908
rect 78674 500896 78680 500908
rect 78732 500896 78738 500948
rect 3418 489812 3424 489864
rect 3476 489852 3482 489864
rect 78674 489852 78680 489864
rect 3476 489824 78680 489852
rect 3476 489812 3482 489824
rect 78674 489812 78680 489824
rect 78732 489812 78738 489864
rect 504358 485800 504364 485852
rect 504416 485840 504422 485852
rect 580166 485840 580172 485852
rect 504416 485812 580172 485840
rect 504416 485800 504422 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 505002 485732 505008 485784
rect 505060 485772 505066 485784
rect 580258 485772 580264 485784
rect 505060 485744 580264 485772
rect 505060 485732 505066 485744
rect 580258 485732 580264 485744
rect 580316 485732 580322 485784
rect 3510 477436 3516 477488
rect 3568 477476 3574 477488
rect 78674 477476 78680 477488
rect 3568 477448 78680 477476
rect 3568 477436 3574 477448
rect 78674 477436 78680 477448
rect 78732 477436 78738 477488
rect 503714 474308 503720 474360
rect 503772 474348 503778 474360
rect 505738 474348 505744 474360
rect 503772 474320 505744 474348
rect 503772 474308 503778 474320
rect 505738 474308 505744 474320
rect 505796 474308 505802 474360
rect 3418 464992 3424 465044
rect 3476 465032 3482 465044
rect 78674 465032 78680 465044
rect 3476 465004 78680 465032
rect 3476 464992 3482 465004
rect 78674 464992 78680 465004
rect 78732 464992 78738 465044
rect 503806 463632 503812 463684
rect 503864 463672 503870 463684
rect 507118 463672 507124 463684
rect 503864 463644 507124 463672
rect 503864 463632 503870 463644
rect 507118 463632 507124 463644
rect 507176 463632 507182 463684
rect 3418 452548 3424 452600
rect 3476 452588 3482 452600
rect 78674 452588 78680 452600
rect 3476 452560 78680 452588
rect 3476 452548 3482 452560
rect 78674 452548 78680 452560
rect 78732 452548 78738 452600
rect 504174 452548 504180 452600
rect 504232 452588 504238 452600
rect 580350 452588 580356 452600
rect 504232 452560 580356 452588
rect 504232 452548 504238 452560
rect 580350 452548 580356 452560
rect 580408 452548 580414 452600
rect 504358 438880 504364 438932
rect 504416 438920 504422 438932
rect 580166 438920 580172 438932
rect 504416 438892 580172 438920
rect 504416 438880 504422 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 78674 438852 78680 438864
rect 3200 438824 78680 438852
rect 3200 438812 3206 438824
rect 78674 438812 78680 438824
rect 78732 438812 78738 438864
rect 505002 430516 505008 430568
rect 505060 430556 505066 430568
rect 580258 430556 580264 430568
rect 505060 430528 580264 430556
rect 505060 430516 505066 430528
rect 580258 430516 580264 430528
rect 580316 430516 580322 430568
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 78674 425048 78680 425060
rect 3292 425020 78680 425048
rect 3292 425008 3298 425020
rect 78674 425008 78680 425020
rect 78732 425008 78738 425060
rect 505002 419432 505008 419484
rect 505060 419472 505066 419484
rect 580442 419472 580448 419484
rect 505060 419444 580448 419472
rect 505060 419432 505066 419444
rect 580442 419432 580448 419444
rect 580500 419432 580506 419484
rect 505002 397400 505008 397452
rect 505060 397440 505066 397452
rect 580350 397440 580356 397452
rect 505060 397412 580356 397440
rect 505060 397400 505066 397412
rect 580350 397400 580356 397412
rect 580408 397400 580414 397452
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 79318 396012 79324 396024
rect 3200 395984 79324 396012
rect 3200 395972 3206 395984
rect 79318 395972 79324 395984
rect 79376 395972 79382 396024
rect 504542 386316 504548 386368
rect 504600 386356 504606 386368
rect 580258 386356 580264 386368
rect 504600 386328 580264 386356
rect 504600 386316 504606 386328
rect 580258 386316 580264 386328
rect 580316 386316 580322 386368
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 79410 380848 79416 380860
rect 3292 380820 79416 380848
rect 3292 380808 3298 380820
rect 79410 380808 79416 380820
rect 79468 380808 79474 380860
rect 505002 375300 505008 375352
rect 505060 375340 505066 375352
rect 580350 375340 580356 375352
rect 505060 375312 580356 375340
rect 505060 375300 505066 375312
rect 580350 375300 580356 375312
rect 580408 375300 580414 375352
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 79318 367044 79324 367056
rect 3200 367016 79324 367044
rect 3200 367004 3206 367016
rect 79318 367004 79324 367016
rect 79376 367004 79382 367056
rect 505002 362856 505008 362908
rect 505060 362896 505066 362908
rect 580258 362896 580264 362908
rect 505060 362868 580264 362896
rect 505060 362856 505066 362868
rect 580258 362856 580264 362868
rect 580316 362856 580322 362908
rect 504634 353200 504640 353252
rect 504692 353240 504698 353252
rect 580258 353240 580264 353252
rect 504692 353212 580264 353240
rect 504692 353200 504698 353212
rect 580258 353200 580264 353212
rect 580316 353200 580322 353252
rect 505002 340824 505008 340876
rect 505060 340864 505066 340876
rect 580902 340864 580908 340876
rect 505060 340836 580908 340864
rect 505060 340824 505066 340836
rect 580902 340824 580908 340836
rect 580960 340824 580966 340876
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 79594 338076 79600 338088
rect 3476 338048 79600 338076
rect 3476 338036 3482 338048
rect 79594 338036 79600 338048
rect 79652 338036 79658 338088
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 79502 324272 79508 324284
rect 3292 324244 79508 324272
rect 3292 324232 3298 324244
rect 79502 324232 79508 324244
rect 79560 324232 79566 324284
rect 504358 322872 504364 322924
rect 504416 322912 504422 322924
rect 580166 322912 580172 322924
rect 504416 322884 580172 322912
rect 504416 322872 504422 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 503806 311788 503812 311840
rect 503864 311828 503870 311840
rect 580166 311828 580172 311840
rect 503864 311800 580172 311828
rect 503864 311788 503870 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 79410 309108 79416 309120
rect 3384 309080 79416 309108
rect 3384 309068 3390 309080
rect 79410 309068 79416 309080
rect 79468 309068 79474 309120
rect 504358 299412 504364 299464
rect 504416 299452 504422 299464
rect 579798 299452 579804 299464
rect 504416 299424 579804 299452
rect 504416 299412 504422 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 79318 295304 79324 295316
rect 3476 295276 79324 295304
rect 3476 295264 3482 295276
rect 79318 295264 79324 295276
rect 79376 295264 79382 295316
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 79686 280140 79692 280152
rect 3476 280112 79692 280140
rect 3476 280100 3482 280112
rect 79686 280100 79692 280112
rect 79744 280100 79750 280152
rect 504358 275952 504364 276004
rect 504416 275992 504422 276004
rect 580166 275992 580172 276004
rect 504416 275964 580172 275992
rect 504416 275952 504422 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 10318 273232 10324 273284
rect 10376 273272 10382 273284
rect 78674 273272 78680 273284
rect 10376 273244 78680 273272
rect 10376 273232 10382 273244
rect 78674 273232 78680 273244
rect 78732 273232 78738 273284
rect 3142 266296 3148 266348
rect 3200 266336 3206 266348
rect 79594 266336 79600 266348
rect 3200 266308 79600 266336
rect 3200 266296 3206 266308
rect 79594 266296 79600 266308
rect 79652 266296 79658 266348
rect 504450 264868 504456 264920
rect 504508 264908 504514 264920
rect 580166 264908 580172 264920
rect 504508 264880 580172 264908
rect 504508 264868 504514 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 79502 252532 79508 252544
rect 3476 252504 79508 252532
rect 3476 252492 3482 252504
rect 79502 252492 79508 252504
rect 79560 252492 79566 252544
rect 504358 252492 504364 252544
rect 504416 252532 504422 252544
rect 579798 252532 579804 252544
rect 504416 252504 579804 252532
rect 504416 252492 504422 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 25498 238756 25504 238808
rect 25556 238796 25562 238808
rect 78674 238796 78680 238808
rect 25556 238768 78680 238796
rect 25556 238756 25562 238768
rect 78674 238756 78680 238768
rect 78732 238756 78738 238808
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 79410 237368 79416 237380
rect 3476 237340 79416 237368
rect 3476 237328 3482 237340
rect 79410 237328 79416 237340
rect 79468 237328 79474 237380
rect 504450 229032 504456 229084
rect 504508 229072 504514 229084
rect 580166 229072 580172 229084
rect 504508 229044 580172 229072
rect 504508 229032 504514 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 79318 223564 79324 223576
rect 3200 223536 79324 223564
rect 3200 223524 3206 223536
rect 79318 223524 79324 223536
rect 79376 223524 79382 223576
rect 504726 217948 504732 218000
rect 504784 217988 504790 218000
rect 580166 217988 580172 218000
rect 504784 217960 580172 217988
rect 504784 217948 504790 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 10318 208332 10324 208344
rect 3476 208304 10324 208332
rect 3476 208292 3482 208304
rect 10318 208292 10324 208304
rect 10376 208292 10382 208344
rect 504358 205572 504364 205624
rect 504416 205612 504422 205624
rect 579798 205612 579804 205624
rect 504416 205584 579804 205612
rect 504416 205572 504422 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 24118 202852 24124 202904
rect 24176 202892 24182 202904
rect 78674 202892 78680 202904
rect 24176 202864 78680 202892
rect 24176 202852 24182 202864
rect 78674 202852 78680 202864
rect 78732 202852 78738 202904
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 79594 194528 79600 194540
rect 3200 194500 79600 194528
rect 3200 194488 3206 194500
rect 79594 194488 79600 194500
rect 79652 194488 79658 194540
rect 504542 182112 504548 182164
rect 504600 182152 504606 182164
rect 580166 182152 580172 182164
rect 504600 182124 580172 182152
rect 504600 182112 504606 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 79502 180792 79508 180804
rect 3292 180764 79508 180792
rect 3292 180752 3298 180764
rect 79502 180752 79508 180764
rect 79560 180752 79566 180804
rect 504634 171028 504640 171080
rect 504692 171068 504698 171080
rect 580166 171068 580172 171080
rect 504692 171040 580172 171068
rect 504692 171028 504698 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 8938 167016 8944 167068
rect 8996 167056 9002 167068
rect 78674 167056 78680 167068
rect 8996 167028 78680 167056
rect 8996 167016 9002 167028
rect 78674 167016 78680 167028
rect 78732 167016 78738 167068
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 25498 165560 25504 165572
rect 3568 165532 25504 165560
rect 3568 165520 3574 165532
rect 25498 165520 25504 165532
rect 25556 165520 25562 165572
rect 504450 158652 504456 158704
rect 504508 158692 504514 158704
rect 579798 158692 579804 158704
rect 504508 158664 579804 158692
rect 504508 158652 504514 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 79410 151756 79416 151768
rect 3200 151728 79416 151756
rect 3200 151716 3206 151728
rect 79410 151716 79416 151728
rect 79468 151716 79474 151768
rect 505002 140768 505008 140820
rect 505060 140808 505066 140820
rect 527818 140808 527824 140820
rect 505060 140780 527824 140808
rect 505060 140768 505066 140780
rect 527818 140768 527824 140780
rect 527876 140768 527882 140820
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 79318 136592 79324 136604
rect 3292 136564 79324 136592
rect 3292 136552 3298 136564
rect 79318 136552 79324 136564
rect 79376 136552 79382 136604
rect 504358 135192 504364 135244
rect 504416 135232 504422 135244
rect 580166 135232 580172 135244
rect 504416 135204 580172 135232
rect 504416 135192 504422 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 14458 131112 14464 131164
rect 14516 131152 14522 131164
rect 78674 131152 78680 131164
rect 14516 131124 78680 131152
rect 14516 131112 14522 131124
rect 78674 131112 78680 131124
rect 78732 131112 78738 131164
rect 504818 124108 504824 124160
rect 504876 124148 504882 124160
rect 580166 124148 580172 124160
rect 504876 124120 580172 124148
rect 504876 124108 504882 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 24118 122788 24124 122800
rect 3476 122760 24124 122788
rect 3476 122748 3482 122760
rect 24118 122748 24124 122760
rect 24176 122748 24182 122800
rect 504726 111732 504732 111784
rect 504784 111772 504790 111784
rect 579798 111772 579804 111784
rect 504784 111744 579804 111772
rect 504784 111732 504790 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 79778 108984 79784 108996
rect 3292 108956 79784 108984
rect 3292 108944 3298 108956
rect 79778 108944 79784 108956
rect 79836 108944 79842 108996
rect 504266 106292 504272 106344
rect 504324 106332 504330 106344
rect 571978 106332 571984 106344
rect 504324 106304 571984 106332
rect 504324 106292 504330 106304
rect 571978 106292 571984 106304
rect 572036 106292 572042 106344
rect 84562 100648 84568 100700
rect 84620 100688 84626 100700
rect 85482 100688 85488 100700
rect 84620 100660 85488 100688
rect 84620 100648 84626 100660
rect 85482 100648 85488 100660
rect 85540 100648 85546 100700
rect 88886 100648 88892 100700
rect 88944 100688 88950 100700
rect 89622 100688 89628 100700
rect 88944 100660 89628 100688
rect 88944 100648 88950 100660
rect 89622 100648 89628 100660
rect 89680 100648 89686 100700
rect 94406 100648 94412 100700
rect 94464 100688 94470 100700
rect 95142 100688 95148 100700
rect 94464 100660 95148 100688
rect 94464 100648 94470 100660
rect 95142 100648 95148 100660
rect 95200 100648 95206 100700
rect 95418 100648 95424 100700
rect 95476 100688 95482 100700
rect 96430 100688 96436 100700
rect 95476 100660 96436 100688
rect 95476 100648 95482 100660
rect 96430 100648 96436 100660
rect 96488 100648 96494 100700
rect 99834 100648 99840 100700
rect 99892 100688 99898 100700
rect 100662 100688 100668 100700
rect 99892 100660 100668 100688
rect 99892 100648 99898 100660
rect 100662 100648 100668 100660
rect 100720 100648 100726 100700
rect 100938 100648 100944 100700
rect 100996 100688 101002 100700
rect 102778 100688 102784 100700
rect 100996 100660 102784 100688
rect 100996 100648 101002 100660
rect 102778 100648 102784 100660
rect 102836 100648 102842 100700
rect 105262 100648 105268 100700
rect 105320 100688 105326 100700
rect 106182 100688 106188 100700
rect 105320 100660 106188 100688
rect 105320 100648 105326 100660
rect 106182 100648 106188 100660
rect 106240 100648 106246 100700
rect 106366 100648 106372 100700
rect 106424 100688 106430 100700
rect 107562 100688 107568 100700
rect 106424 100660 107568 100688
rect 106424 100648 106430 100660
rect 107562 100648 107568 100660
rect 107620 100648 107626 100700
rect 156414 100648 156420 100700
rect 156472 100688 156478 100700
rect 157242 100688 157248 100700
rect 156472 100660 157248 100688
rect 156472 100648 156478 100660
rect 157242 100648 157248 100660
rect 157300 100648 157306 100700
rect 228174 100648 228180 100700
rect 228232 100688 228238 100700
rect 229002 100688 229008 100700
rect 228232 100660 229008 100688
rect 228232 100648 228238 100660
rect 229002 100648 229008 100660
rect 229060 100648 229066 100700
rect 229278 100648 229284 100700
rect 229336 100688 229342 100700
rect 230382 100688 230388 100700
rect 229336 100660 230388 100688
rect 229336 100648 229342 100660
rect 230382 100648 230388 100660
rect 230440 100648 230446 100700
rect 233602 100648 233608 100700
rect 233660 100688 233666 100700
rect 234522 100688 234528 100700
rect 233660 100660 234528 100688
rect 233660 100648 233666 100660
rect 234522 100648 234528 100660
rect 234580 100648 234586 100700
rect 243446 100648 243452 100700
rect 243504 100688 243510 100700
rect 244182 100688 244188 100700
rect 243504 100660 244188 100688
rect 243504 100648 243510 100660
rect 244182 100648 244188 100660
rect 244240 100648 244246 100700
rect 321738 100648 321744 100700
rect 321796 100688 321802 100700
rect 322750 100688 322756 100700
rect 321796 100660 322756 100688
rect 321796 100648 321802 100660
rect 322750 100648 322756 100660
rect 322808 100648 322814 100700
rect 327166 100648 327172 100700
rect 327224 100688 327230 100700
rect 329098 100688 329104 100700
rect 327224 100660 329104 100688
rect 327224 100648 327230 100660
rect 329098 100648 329104 100660
rect 329156 100648 329162 100700
rect 331582 100648 331588 100700
rect 331640 100688 331646 100700
rect 332502 100688 332508 100700
rect 331640 100660 332508 100688
rect 331640 100648 331646 100660
rect 332502 100648 332508 100660
rect 332560 100648 332566 100700
rect 337010 100648 337016 100700
rect 337068 100688 337074 100700
rect 338022 100688 338028 100700
rect 337068 100660 338028 100688
rect 337068 100648 337074 100660
rect 338022 100648 338028 100660
rect 338080 100648 338086 100700
rect 338114 100648 338120 100700
rect 338172 100688 338178 100700
rect 339310 100688 339316 100700
rect 338172 100660 339316 100688
rect 338172 100648 338178 100660
rect 339310 100648 339316 100660
rect 339368 100648 339374 100700
rect 392486 100648 392492 100700
rect 392544 100688 392550 100700
rect 393222 100688 393228 100700
rect 392544 100660 393228 100688
rect 392544 100648 392550 100660
rect 393222 100648 393228 100660
rect 393280 100648 393286 100700
rect 397914 100648 397920 100700
rect 397972 100688 397978 100700
rect 398742 100688 398748 100700
rect 397972 100660 398748 100688
rect 397972 100648 397978 100660
rect 398742 100648 398748 100660
rect 398800 100648 398806 100700
rect 408770 100648 408776 100700
rect 408828 100688 408834 100700
rect 409782 100688 409788 100700
rect 408828 100660 409788 100688
rect 408828 100648 408834 100660
rect 409782 100648 409788 100660
rect 409840 100648 409846 100700
rect 418614 100648 418620 100700
rect 418672 100688 418678 100700
rect 419442 100688 419448 100700
rect 418672 100660 419448 100688
rect 418672 100648 418678 100660
rect 419442 100648 419448 100660
rect 419500 100648 419506 100700
rect 424042 100648 424048 100700
rect 424100 100688 424106 100700
rect 424962 100688 424968 100700
rect 424100 100660 424968 100688
rect 424100 100648 424106 100660
rect 424962 100648 424968 100660
rect 425020 100648 425026 100700
rect 425146 100648 425152 100700
rect 425204 100688 425210 100700
rect 427078 100688 427084 100700
rect 425204 100660 427084 100688
rect 425204 100648 425210 100660
rect 427078 100648 427084 100660
rect 427136 100648 427142 100700
rect 459922 100648 459928 100700
rect 459980 100688 459986 100700
rect 460842 100688 460848 100700
rect 459980 100660 460848 100688
rect 459980 100648 459986 100660
rect 460842 100648 460848 100660
rect 460900 100648 460906 100700
rect 461026 100648 461032 100700
rect 461084 100688 461090 100700
rect 462958 100688 462964 100700
rect 461084 100660 462964 100688
rect 461084 100648 461090 100660
rect 462958 100648 462964 100660
rect 463016 100648 463022 100700
rect 476298 100648 476304 100700
rect 476356 100688 476362 100700
rect 478230 100688 478236 100700
rect 476356 100660 478236 100688
rect 476356 100648 476362 100660
rect 478230 100648 478236 100660
rect 478288 100648 478294 100700
rect 480622 100648 480628 100700
rect 480680 100688 480686 100700
rect 481542 100688 481548 100700
rect 480680 100660 481548 100688
rect 480680 100648 480686 100660
rect 481542 100648 481548 100660
rect 481600 100648 481606 100700
rect 481726 100648 481732 100700
rect 481784 100688 481790 100700
rect 482922 100688 482928 100700
rect 481784 100660 482928 100688
rect 481784 100648 481790 100660
rect 482922 100648 482928 100660
rect 482980 100648 482986 100700
rect 91094 100580 91100 100632
rect 91152 100620 91158 100632
rect 92382 100620 92388 100632
rect 91152 100592 92388 100620
rect 91152 100580 91158 100592
rect 92382 100580 92388 100592
rect 92440 100580 92446 100632
rect 240134 100580 240140 100632
rect 240192 100620 240198 100632
rect 241330 100620 241336 100632
rect 240192 100592 241336 100620
rect 240192 100580 240198 100592
rect 241330 100580 241336 100592
rect 241388 100580 241394 100632
rect 326154 100512 326160 100564
rect 326212 100552 326218 100564
rect 326982 100552 326988 100564
rect 326212 100524 326988 100552
rect 326212 100512 326218 100524
rect 326982 100512 326988 100524
rect 327040 100512 327046 100564
rect 153102 100444 153108 100496
rect 153160 100484 153166 100496
rect 153838 100484 153844 100496
rect 153160 100456 153844 100484
rect 153160 100444 153166 100456
rect 153838 100444 153844 100456
rect 153896 100444 153902 100496
rect 295610 100172 295616 100224
rect 295668 100212 295674 100224
rect 296622 100212 296628 100224
rect 295668 100184 296628 100212
rect 295668 100172 295674 100184
rect 296622 100172 296628 100184
rect 296680 100172 296686 100224
rect 301130 100172 301136 100224
rect 301188 100212 301194 100224
rect 302142 100212 302148 100224
rect 301188 100184 302148 100212
rect 301188 100172 301194 100184
rect 302142 100172 302148 100184
rect 302200 100172 302206 100224
rect 211890 100036 211896 100088
rect 211948 100076 211954 100088
rect 231118 100076 231124 100088
rect 211948 100048 231124 100076
rect 211948 100036 211954 100048
rect 231118 100036 231124 100048
rect 231176 100036 231182 100088
rect 286962 100036 286968 100088
rect 287020 100076 287026 100088
rect 323578 100076 323584 100088
rect 287020 100048 323584 100076
rect 287020 100036 287026 100048
rect 323578 100036 323584 100048
rect 323636 100036 323642 100088
rect 325050 100036 325056 100088
rect 325108 100076 325114 100088
rect 337378 100076 337384 100088
rect 325108 100048 337384 100076
rect 325108 100036 325114 100048
rect 337378 100036 337384 100048
rect 337436 100036 337442 100088
rect 353294 100036 353300 100088
rect 353352 100076 353358 100088
rect 362218 100076 362224 100088
rect 353352 100048 362224 100076
rect 353352 100036 353358 100048
rect 362218 100036 362224 100048
rect 362276 100036 362282 100088
rect 385954 100036 385960 100088
rect 386012 100076 386018 100088
rect 411898 100076 411904 100088
rect 386012 100048 411904 100076
rect 386012 100036 386018 100048
rect 411898 100036 411904 100048
rect 411956 100036 411962 100088
rect 414290 100036 414296 100088
rect 414348 100076 414354 100088
rect 438118 100076 438124 100088
rect 414348 100048 438124 100076
rect 414348 100036 414354 100048
rect 438118 100036 438124 100048
rect 438176 100036 438182 100088
rect 492582 100036 492588 100088
rect 492640 100076 492646 100088
rect 560938 100076 560944 100088
rect 492640 100048 560944 100076
rect 492640 100036 492646 100048
rect 560938 100036 560944 100048
rect 560996 100036 561002 100088
rect 85666 99968 85672 100020
rect 85724 100008 85730 100020
rect 97258 100008 97264 100020
rect 85724 99980 97264 100008
rect 85724 99968 85730 99980
rect 97258 99968 97264 99980
rect 97316 99968 97322 100020
rect 117222 99968 117228 100020
rect 117280 100008 117286 100020
rect 161566 100008 161572 100020
rect 117280 99980 161572 100008
rect 117280 99968 117286 99980
rect 161566 99968 161572 99980
rect 161624 99968 161630 100020
rect 162946 99968 162952 100020
rect 163004 100008 163010 100020
rect 211154 100008 211160 100020
rect 163004 99980 211160 100008
rect 163004 99968 163010 99980
rect 211154 99968 211160 99980
rect 211212 99968 211218 100020
rect 231486 99968 231492 100020
rect 231544 100008 231550 100020
rect 287238 100008 287244 100020
rect 231544 99980 287244 100008
rect 231544 99968 231550 99980
rect 287238 99968 287244 99980
rect 287296 99968 287302 100020
rect 329374 99968 329380 100020
rect 329432 100008 329438 100020
rect 393406 100008 393412 100020
rect 329432 99980 393412 100008
rect 329432 99968 329438 99980
rect 393406 99968 393412 99980
rect 393464 99968 393470 100020
rect 430574 99968 430580 100020
rect 430632 100008 430638 100020
rect 502978 100008 502984 100020
rect 430632 99980 502984 100008
rect 430632 99968 430638 99980
rect 502978 99968 502984 99980
rect 503036 99968 503042 100020
rect 224954 99764 224960 99816
rect 225012 99804 225018 99816
rect 226242 99804 226248 99816
rect 225012 99776 226248 99804
rect 225012 99764 225018 99776
rect 226242 99764 226248 99776
rect 226300 99764 226306 99816
rect 409874 99764 409880 99816
rect 409932 99804 409938 99816
rect 411162 99804 411168 99816
rect 409932 99776 411168 99804
rect 409932 99764 409938 99776
rect 411162 99764 411168 99776
rect 411220 99764 411226 99816
rect 419718 99764 419724 99816
rect 419776 99804 419782 99816
rect 420730 99804 420736 99816
rect 419776 99776 420736 99804
rect 419776 99764 419782 99776
rect 420730 99764 420736 99776
rect 420788 99764 420794 99816
rect 239122 99696 239128 99748
rect 239180 99736 239186 99748
rect 240042 99736 240048 99748
rect 239180 99708 240048 99736
rect 239180 99696 239186 99708
rect 240042 99696 240048 99708
rect 240100 99696 240106 99748
rect 332686 99696 332692 99748
rect 332744 99736 332750 99748
rect 333882 99736 333888 99748
rect 332744 99708 333888 99736
rect 332744 99696 332750 99708
rect 333882 99696 333888 99708
rect 333940 99696 333946 99748
rect 393590 99696 393596 99748
rect 393648 99736 393654 99748
rect 394602 99736 394608 99748
rect 393648 99708 394608 99736
rect 393648 99696 393654 99708
rect 394602 99696 394608 99708
rect 394660 99696 394666 99748
rect 465350 99696 465356 99748
rect 465408 99736 465414 99748
rect 466362 99736 466368 99748
rect 465408 99708 466368 99736
rect 465408 99696 465414 99708
rect 466362 99696 466368 99708
rect 466420 99696 466426 99748
rect 89990 99560 89996 99612
rect 90048 99600 90054 99612
rect 91002 99600 91008 99612
rect 90048 99572 91008 99600
rect 90048 99560 90054 99572
rect 91002 99560 91008 99572
rect 91060 99560 91066 99612
rect 296714 99560 296720 99612
rect 296772 99600 296778 99612
rect 298002 99600 298008 99612
rect 296772 99572 298008 99600
rect 296772 99560 296778 99572
rect 298002 99560 298008 99572
rect 298060 99560 298066 99612
rect 394694 99560 394700 99612
rect 394752 99600 394758 99612
rect 395982 99600 395988 99612
rect 394752 99572 395988 99600
rect 394752 99560 394758 99572
rect 395982 99560 395988 99572
rect 396040 99560 396046 99612
rect 107470 99424 107476 99476
rect 107528 99464 107534 99476
rect 113818 99464 113824 99476
rect 107528 99436 113824 99464
rect 107528 99424 107534 99436
rect 113818 99424 113824 99436
rect 113876 99424 113882 99476
rect 110690 99356 110696 99408
rect 110748 99396 110754 99408
rect 111702 99396 111708 99408
rect 110748 99368 111708 99396
rect 110748 99356 110754 99368
rect 111702 99356 111708 99368
rect 111760 99356 111766 99408
rect 115014 99356 115020 99408
rect 115072 99396 115078 99408
rect 115842 99396 115848 99408
rect 115072 99368 115848 99396
rect 115072 99356 115078 99368
rect 115842 99356 115848 99368
rect 115900 99356 115906 99408
rect 116118 99356 116124 99408
rect 116176 99396 116182 99408
rect 117222 99396 117228 99408
rect 116176 99368 117228 99396
rect 116176 99356 116182 99368
rect 117222 99356 117228 99368
rect 117280 99356 117286 99408
rect 120442 99356 120448 99408
rect 120500 99396 120506 99408
rect 121362 99396 121368 99408
rect 120500 99368 121368 99396
rect 120500 99356 120506 99368
rect 121362 99356 121368 99368
rect 121420 99356 121426 99408
rect 121546 99356 121552 99408
rect 121604 99396 121610 99408
rect 122742 99396 122748 99408
rect 121604 99368 122748 99396
rect 121604 99356 121610 99368
rect 122742 99356 122748 99368
rect 122800 99356 122806 99408
rect 125962 99356 125968 99408
rect 126020 99396 126026 99408
rect 126882 99396 126888 99408
rect 126020 99368 126888 99396
rect 126020 99356 126026 99368
rect 126882 99356 126888 99368
rect 126940 99356 126946 99408
rect 126974 99356 126980 99408
rect 127032 99396 127038 99408
rect 128998 99396 129004 99408
rect 127032 99368 129004 99396
rect 127032 99356 127038 99368
rect 128998 99356 129004 99368
rect 129056 99356 129062 99408
rect 130286 99356 130292 99408
rect 130344 99396 130350 99408
rect 131022 99396 131028 99408
rect 130344 99368 131028 99396
rect 130344 99356 130350 99368
rect 131022 99356 131028 99368
rect 131080 99356 131086 99408
rect 131390 99356 131396 99408
rect 131448 99396 131454 99408
rect 132402 99396 132408 99408
rect 131448 99368 132408 99396
rect 131448 99356 131454 99368
rect 132402 99356 132408 99368
rect 132460 99356 132466 99408
rect 132494 99356 132500 99408
rect 132552 99396 132558 99408
rect 133690 99396 133696 99408
rect 132552 99368 133696 99396
rect 132552 99356 132558 99368
rect 133690 99356 133696 99368
rect 133748 99356 133754 99408
rect 135714 99356 135720 99408
rect 135772 99396 135778 99408
rect 136542 99396 136548 99408
rect 135772 99368 136548 99396
rect 135772 99356 135778 99368
rect 136542 99356 136548 99368
rect 136600 99356 136606 99408
rect 136818 99356 136824 99408
rect 136876 99396 136882 99408
rect 138658 99396 138664 99408
rect 136876 99368 138664 99396
rect 136876 99356 136882 99368
rect 138658 99356 138664 99368
rect 138716 99356 138722 99408
rect 141142 99356 141148 99408
rect 141200 99396 141206 99408
rect 142062 99396 142068 99408
rect 141200 99368 142068 99396
rect 141200 99356 141206 99368
rect 142062 99356 142068 99368
rect 142120 99356 142126 99408
rect 142246 99356 142252 99408
rect 142304 99396 142310 99408
rect 143350 99396 143356 99408
rect 142304 99368 143356 99396
rect 142304 99356 142310 99368
rect 143350 99356 143356 99368
rect 143408 99356 143414 99408
rect 146570 99356 146576 99408
rect 146628 99396 146634 99408
rect 147582 99396 147588 99408
rect 146628 99368 147588 99396
rect 146628 99356 146634 99368
rect 147582 99356 147588 99368
rect 147640 99356 147646 99408
rect 151998 99356 152004 99408
rect 152056 99396 152062 99408
rect 152056 99368 153056 99396
rect 152056 99356 152062 99368
rect 153028 99340 153056 99368
rect 157518 99356 157524 99408
rect 157576 99396 157582 99408
rect 158622 99396 158628 99408
rect 157576 99368 158628 99396
rect 157576 99356 157582 99368
rect 158622 99356 158628 99368
rect 158680 99356 158686 99408
rect 161842 99356 161848 99408
rect 161900 99396 161906 99408
rect 162762 99396 162768 99408
rect 161900 99368 162768 99396
rect 161900 99356 161906 99368
rect 162762 99356 162768 99368
rect 162820 99356 162826 99408
rect 166166 99356 166172 99408
rect 166224 99396 166230 99408
rect 166902 99396 166908 99408
rect 166224 99368 166908 99396
rect 166224 99356 166230 99368
rect 166902 99356 166908 99368
rect 166960 99356 166966 99408
rect 167270 99356 167276 99408
rect 167328 99396 167334 99408
rect 168282 99396 168288 99408
rect 167328 99368 168288 99396
rect 167328 99356 167334 99368
rect 168282 99356 168288 99368
rect 168340 99356 168346 99408
rect 168374 99356 168380 99408
rect 168432 99396 168438 99408
rect 169570 99396 169576 99408
rect 168432 99368 169576 99396
rect 168432 99356 168438 99368
rect 169570 99356 169576 99368
rect 169628 99356 169634 99408
rect 171594 99356 171600 99408
rect 171652 99396 171658 99408
rect 172422 99396 172428 99408
rect 171652 99368 172428 99396
rect 171652 99356 171658 99368
rect 172422 99356 172428 99368
rect 172480 99356 172486 99408
rect 172698 99356 172704 99408
rect 172756 99396 172762 99408
rect 173802 99396 173808 99408
rect 172756 99368 173808 99396
rect 172756 99356 172762 99368
rect 173802 99356 173808 99368
rect 173860 99356 173866 99408
rect 177022 99356 177028 99408
rect 177080 99396 177086 99408
rect 177942 99396 177948 99408
rect 177080 99368 177948 99396
rect 177080 99356 177086 99368
rect 177942 99356 177948 99368
rect 178000 99356 178006 99408
rect 178126 99356 178132 99408
rect 178184 99396 178190 99408
rect 179230 99396 179236 99408
rect 178184 99368 179236 99396
rect 178184 99356 178190 99368
rect 179230 99356 179236 99368
rect 179288 99356 179294 99408
rect 182542 99356 182548 99408
rect 182600 99396 182606 99408
rect 183462 99396 183468 99408
rect 182600 99368 183468 99396
rect 182600 99356 182606 99368
rect 183462 99356 183468 99368
rect 183520 99356 183526 99408
rect 183554 99356 183560 99408
rect 183612 99396 183618 99408
rect 185578 99396 185584 99408
rect 183612 99368 185584 99396
rect 183612 99356 183618 99368
rect 185578 99356 185584 99368
rect 185636 99356 185642 99408
rect 187970 99356 187976 99408
rect 188028 99396 188034 99408
rect 188028 99368 188936 99396
rect 188028 99356 188034 99368
rect 153010 99288 153016 99340
rect 153068 99288 153074 99340
rect 188908 99260 188936 99368
rect 188982 99356 188988 99408
rect 189040 99396 189046 99408
rect 189718 99396 189724 99408
rect 189040 99368 189724 99396
rect 189040 99356 189046 99368
rect 189718 99356 189724 99368
rect 189776 99356 189782 99408
rect 192294 99356 192300 99408
rect 192352 99396 192358 99408
rect 193122 99396 193128 99408
rect 192352 99368 193128 99396
rect 192352 99356 192358 99368
rect 193122 99356 193128 99368
rect 193180 99356 193186 99408
rect 193398 99356 193404 99408
rect 193456 99396 193462 99408
rect 194502 99396 194508 99408
rect 193456 99368 194508 99396
rect 193456 99356 193462 99368
rect 194502 99356 194508 99368
rect 194560 99356 194566 99408
rect 197722 99356 197728 99408
rect 197780 99396 197786 99408
rect 198642 99396 198648 99408
rect 197780 99368 198648 99396
rect 197780 99356 197786 99368
rect 198642 99356 198648 99368
rect 198700 99356 198706 99408
rect 202046 99356 202052 99408
rect 202104 99396 202110 99408
rect 202782 99396 202788 99408
rect 202104 99368 202788 99396
rect 202104 99356 202110 99368
rect 202782 99356 202788 99368
rect 202840 99356 202846 99408
rect 203150 99356 203156 99408
rect 203208 99396 203214 99408
rect 204162 99396 204168 99408
rect 203208 99368 204168 99396
rect 203208 99356 203214 99368
rect 204162 99356 204168 99368
rect 204220 99356 204226 99408
rect 204254 99356 204260 99408
rect 204312 99396 204318 99408
rect 205450 99396 205456 99408
rect 204312 99368 205456 99396
rect 204312 99356 204318 99368
rect 205450 99356 205456 99368
rect 205508 99356 205514 99408
rect 207566 99356 207572 99408
rect 207624 99396 207630 99408
rect 208302 99396 208308 99408
rect 207624 99368 208308 99396
rect 207624 99356 207630 99368
rect 208302 99356 208308 99368
rect 208360 99356 208366 99408
rect 208578 99356 208584 99408
rect 208636 99396 208642 99408
rect 209682 99396 209688 99408
rect 208636 99368 209688 99396
rect 208636 99356 208642 99368
rect 209682 99356 209688 99368
rect 209740 99356 209746 99408
rect 212994 99356 213000 99408
rect 213052 99396 213058 99408
rect 213822 99396 213828 99408
rect 213052 99368 213828 99396
rect 213052 99356 213058 99368
rect 213822 99356 213828 99368
rect 213880 99356 213886 99408
rect 214006 99356 214012 99408
rect 214064 99396 214070 99408
rect 215110 99396 215116 99408
rect 214064 99368 215116 99396
rect 214064 99356 214070 99368
rect 215110 99356 215116 99368
rect 215168 99356 215174 99408
rect 218422 99356 218428 99408
rect 218480 99396 218486 99408
rect 219342 99396 219348 99408
rect 218480 99368 219348 99396
rect 218480 99356 218486 99368
rect 219342 99356 219348 99368
rect 219400 99356 219406 99408
rect 220538 99356 220544 99408
rect 220596 99396 220602 99408
rect 221458 99396 221464 99408
rect 220596 99368 221464 99396
rect 220596 99356 220602 99368
rect 221458 99356 221464 99368
rect 221516 99356 221522 99408
rect 223850 99356 223856 99408
rect 223908 99396 223914 99408
rect 224862 99396 224868 99408
rect 223908 99368 224868 99396
rect 223908 99356 223914 99368
rect 224862 99356 224868 99368
rect 224920 99356 224926 99408
rect 244550 99356 244556 99408
rect 244608 99396 244614 99408
rect 245562 99396 245568 99408
rect 244608 99368 245568 99396
rect 244608 99356 244614 99368
rect 245562 99356 245568 99368
rect 245620 99356 245626 99408
rect 248874 99356 248880 99408
rect 248932 99396 248938 99408
rect 249702 99396 249708 99408
rect 248932 99368 249708 99396
rect 248932 99356 248938 99368
rect 249702 99356 249708 99368
rect 249760 99356 249766 99408
rect 249978 99356 249984 99408
rect 250036 99396 250042 99408
rect 250990 99396 250996 99408
rect 250036 99368 250996 99396
rect 250036 99356 250042 99368
rect 250990 99356 250996 99368
rect 251048 99356 251054 99408
rect 254302 99356 254308 99408
rect 254360 99396 254366 99408
rect 255222 99396 255228 99408
rect 254360 99368 255228 99396
rect 254360 99356 254366 99368
rect 255222 99356 255228 99368
rect 255280 99356 255286 99408
rect 255406 99356 255412 99408
rect 255464 99396 255470 99408
rect 256602 99396 256608 99408
rect 255464 99368 256608 99396
rect 255464 99356 255470 99368
rect 256602 99356 256608 99368
rect 256660 99356 256666 99408
rect 259730 99356 259736 99408
rect 259788 99396 259794 99408
rect 260742 99396 260748 99408
rect 259788 99368 260748 99396
rect 259788 99356 259794 99368
rect 260742 99356 260748 99368
rect 260800 99356 260806 99408
rect 260834 99356 260840 99408
rect 260892 99396 260898 99408
rect 262030 99396 262036 99408
rect 260892 99368 262036 99396
rect 260892 99356 260898 99368
rect 262030 99356 262036 99368
rect 262088 99356 262094 99408
rect 265158 99356 265164 99408
rect 265216 99396 265222 99408
rect 266170 99396 266176 99408
rect 265216 99368 266176 99396
rect 265216 99356 265222 99368
rect 266170 99356 266176 99368
rect 266228 99356 266234 99408
rect 269574 99356 269580 99408
rect 269632 99396 269638 99408
rect 270402 99396 270408 99408
rect 269632 99368 270408 99396
rect 269632 99356 269638 99368
rect 270402 99356 270408 99368
rect 270460 99356 270466 99408
rect 275002 99356 275008 99408
rect 275060 99396 275066 99408
rect 275922 99396 275928 99408
rect 275060 99368 275928 99396
rect 275060 99356 275066 99368
rect 275922 99356 275928 99368
rect 275980 99356 275986 99408
rect 276106 99356 276112 99408
rect 276164 99396 276170 99408
rect 277210 99396 277216 99408
rect 276164 99368 277216 99396
rect 276164 99356 276170 99368
rect 277210 99356 277216 99368
rect 277268 99356 277274 99408
rect 279326 99356 279332 99408
rect 279384 99396 279390 99408
rect 280062 99396 280068 99408
rect 279384 99368 280068 99396
rect 279384 99356 279390 99368
rect 280062 99356 280068 99368
rect 280120 99356 280126 99408
rect 280430 99356 280436 99408
rect 280488 99396 280494 99408
rect 281442 99396 281448 99408
rect 280488 99368 281448 99396
rect 280488 99356 280494 99368
rect 281442 99356 281448 99368
rect 281500 99356 281506 99408
rect 284754 99356 284760 99408
rect 284812 99396 284818 99408
rect 285582 99396 285588 99408
rect 284812 99368 285588 99396
rect 284812 99356 284818 99368
rect 285582 99356 285588 99368
rect 285640 99356 285646 99408
rect 285858 99356 285864 99408
rect 285916 99396 285922 99408
rect 286962 99396 286968 99408
rect 285916 99368 286968 99396
rect 285916 99356 285922 99368
rect 286962 99356 286968 99368
rect 287020 99356 287026 99408
rect 290182 99356 290188 99408
rect 290240 99396 290246 99408
rect 291102 99396 291108 99408
rect 290240 99368 291108 99396
rect 290240 99356 290246 99368
rect 291102 99356 291108 99368
rect 291160 99356 291166 99408
rect 291286 99356 291292 99408
rect 291344 99396 291350 99408
rect 292482 99396 292488 99408
rect 291344 99368 292488 99396
rect 291344 99356 291350 99368
rect 292482 99356 292488 99368
rect 292540 99356 292546 99408
rect 305454 99356 305460 99408
rect 305512 99396 305518 99408
rect 306282 99396 306288 99408
rect 305512 99368 306288 99396
rect 305512 99356 305518 99368
rect 306282 99356 306288 99368
rect 306340 99356 306346 99408
rect 306558 99356 306564 99408
rect 306616 99396 306622 99408
rect 309778 99396 309784 99408
rect 306616 99368 309784 99396
rect 306616 99356 306622 99368
rect 309778 99356 309784 99368
rect 309836 99356 309842 99408
rect 310882 99356 310888 99408
rect 310940 99396 310946 99408
rect 311802 99396 311808 99408
rect 310940 99368 311808 99396
rect 310940 99356 310946 99368
rect 311802 99356 311808 99368
rect 311860 99356 311866 99408
rect 311986 99356 311992 99408
rect 312044 99396 312050 99408
rect 313090 99396 313096 99408
rect 312044 99368 313096 99396
rect 312044 99356 312050 99368
rect 313090 99356 313096 99368
rect 313148 99356 313154 99408
rect 315206 99356 315212 99408
rect 315264 99396 315270 99408
rect 315942 99396 315948 99408
rect 315264 99368 315948 99396
rect 315264 99356 315270 99368
rect 315942 99356 315948 99368
rect 316000 99356 316006 99408
rect 316310 99356 316316 99408
rect 316368 99396 316374 99408
rect 317322 99396 317328 99408
rect 316368 99368 317328 99396
rect 316368 99356 316374 99368
rect 317322 99356 317328 99368
rect 317380 99356 317386 99408
rect 320634 99356 320640 99408
rect 320692 99396 320698 99408
rect 321462 99396 321468 99408
rect 320692 99368 321468 99396
rect 320692 99356 320698 99368
rect 321462 99356 321468 99368
rect 321520 99356 321526 99408
rect 341334 99356 341340 99408
rect 341392 99396 341398 99408
rect 342162 99396 342168 99408
rect 341392 99368 342168 99396
rect 341392 99356 341398 99368
rect 342162 99356 342168 99368
rect 342220 99356 342226 99408
rect 343542 99356 343548 99408
rect 343600 99396 343606 99408
rect 345658 99396 345664 99408
rect 343600 99368 345664 99396
rect 343600 99356 343606 99368
rect 345658 99356 345664 99368
rect 345716 99356 345722 99408
rect 346762 99356 346768 99408
rect 346820 99396 346826 99408
rect 347682 99396 347688 99408
rect 346820 99368 347688 99396
rect 346820 99356 346826 99368
rect 347682 99356 347688 99368
rect 347740 99356 347746 99408
rect 347866 99356 347872 99408
rect 347924 99396 347930 99408
rect 348970 99396 348976 99408
rect 347924 99368 348976 99396
rect 347924 99356 347930 99368
rect 348970 99356 348976 99368
rect 349028 99356 349034 99408
rect 352190 99356 352196 99408
rect 352248 99396 352254 99408
rect 353202 99396 353208 99408
rect 352248 99368 353208 99396
rect 352248 99356 352254 99368
rect 353202 99356 353208 99368
rect 353260 99356 353266 99408
rect 356606 99356 356612 99408
rect 356664 99396 356670 99408
rect 357342 99396 357348 99408
rect 356664 99368 357348 99396
rect 356664 99356 356670 99368
rect 357342 99356 357348 99368
rect 357400 99356 357406 99408
rect 357710 99356 357716 99408
rect 357768 99396 357774 99408
rect 358630 99396 358636 99408
rect 357768 99368 358636 99396
rect 357768 99356 357774 99368
rect 358630 99356 358636 99368
rect 358688 99356 358694 99408
rect 362034 99356 362040 99408
rect 362092 99396 362098 99408
rect 362862 99396 362868 99408
rect 362092 99368 362868 99396
rect 362092 99356 362098 99368
rect 362862 99356 362868 99368
rect 362920 99356 362926 99408
rect 363138 99356 363144 99408
rect 363196 99396 363202 99408
rect 364150 99396 364156 99408
rect 363196 99368 364156 99396
rect 363196 99356 363202 99368
rect 364150 99356 364156 99368
rect 364208 99356 364214 99408
rect 367462 99356 367468 99408
rect 367520 99396 367526 99408
rect 368382 99396 368388 99408
rect 367520 99368 368388 99396
rect 367520 99356 367526 99368
rect 368382 99356 368388 99368
rect 368440 99356 368446 99408
rect 368566 99356 368572 99408
rect 368624 99396 368630 99408
rect 369762 99396 369768 99408
rect 368624 99368 369768 99396
rect 368624 99356 368630 99368
rect 369762 99356 369768 99368
rect 369820 99356 369826 99408
rect 372890 99356 372896 99408
rect 372948 99396 372954 99408
rect 373902 99396 373908 99408
rect 372948 99368 373908 99396
rect 372948 99356 372954 99368
rect 373902 99356 373908 99368
rect 373960 99356 373966 99408
rect 373994 99356 374000 99408
rect 374052 99396 374058 99408
rect 375190 99396 375196 99408
rect 374052 99368 375196 99396
rect 374052 99356 374058 99368
rect 375190 99356 375196 99368
rect 375248 99356 375254 99408
rect 377214 99356 377220 99408
rect 377272 99396 377278 99408
rect 378042 99396 378048 99408
rect 377272 99368 378048 99396
rect 377272 99356 377278 99368
rect 378042 99356 378048 99368
rect 378100 99356 378106 99408
rect 378318 99356 378324 99408
rect 378376 99396 378382 99408
rect 380158 99396 380164 99408
rect 378376 99368 380164 99396
rect 378376 99356 378382 99368
rect 380158 99356 380164 99368
rect 380216 99356 380222 99408
rect 382734 99356 382740 99408
rect 382792 99396 382798 99408
rect 383562 99396 383568 99408
rect 382792 99368 383568 99396
rect 382792 99356 382798 99368
rect 383562 99356 383568 99368
rect 383620 99356 383626 99408
rect 383746 99356 383752 99408
rect 383804 99396 383810 99408
rect 384942 99396 384948 99408
rect 383804 99368 384948 99396
rect 383804 99356 383810 99368
rect 384942 99356 384948 99368
rect 385000 99356 385006 99408
rect 388162 99356 388168 99408
rect 388220 99396 388226 99408
rect 389082 99396 389088 99408
rect 388220 99368 389088 99396
rect 388220 99356 388226 99368
rect 389082 99356 389088 99368
rect 389140 99356 389146 99408
rect 399018 99356 399024 99408
rect 399076 99396 399082 99408
rect 400030 99396 400036 99408
rect 399076 99368 400036 99396
rect 399076 99356 399082 99368
rect 400030 99356 400036 99368
rect 400088 99356 400094 99408
rect 403342 99356 403348 99408
rect 403400 99396 403406 99408
rect 404262 99396 404268 99408
rect 403400 99368 404268 99396
rect 403400 99356 403406 99368
rect 404262 99356 404268 99368
rect 404320 99356 404326 99408
rect 404446 99356 404452 99408
rect 404504 99396 404510 99408
rect 405642 99396 405648 99408
rect 404504 99368 405648 99396
rect 404504 99356 404510 99368
rect 405642 99356 405648 99368
rect 405700 99356 405706 99408
rect 428366 99356 428372 99408
rect 428424 99396 428430 99408
rect 429102 99396 429108 99408
rect 428424 99368 429108 99396
rect 428424 99356 428430 99368
rect 429102 99356 429108 99368
rect 429160 99356 429166 99408
rect 429470 99356 429476 99408
rect 429528 99396 429534 99408
rect 430482 99396 430488 99408
rect 429528 99368 430488 99396
rect 429528 99356 429534 99368
rect 430482 99356 430488 99368
rect 430540 99356 430546 99408
rect 433794 99356 433800 99408
rect 433852 99396 433858 99408
rect 434622 99396 434628 99408
rect 433852 99368 434628 99396
rect 433852 99356 433858 99368
rect 434622 99356 434628 99368
rect 434680 99356 434686 99408
rect 434898 99356 434904 99408
rect 434956 99396 434962 99408
rect 435910 99396 435916 99408
rect 434956 99368 435916 99396
rect 434956 99356 434962 99368
rect 435910 99356 435916 99368
rect 435968 99356 435974 99408
rect 439314 99356 439320 99408
rect 439372 99396 439378 99408
rect 440142 99396 440148 99408
rect 439372 99368 440148 99396
rect 439372 99356 439378 99368
rect 440142 99356 440148 99368
rect 440200 99356 440206 99408
rect 444742 99356 444748 99408
rect 444800 99396 444806 99408
rect 445662 99396 445668 99408
rect 444800 99368 445668 99396
rect 444800 99356 444806 99368
rect 445662 99356 445668 99368
rect 445720 99356 445726 99408
rect 445846 99356 445852 99408
rect 445904 99396 445910 99408
rect 447042 99396 447048 99408
rect 445904 99368 447048 99396
rect 445904 99356 445910 99368
rect 447042 99356 447048 99368
rect 447100 99356 447106 99408
rect 450170 99356 450176 99408
rect 450228 99396 450234 99408
rect 451182 99396 451188 99408
rect 450228 99368 451188 99396
rect 450228 99356 450234 99368
rect 451182 99356 451188 99368
rect 451240 99356 451246 99408
rect 451274 99356 451280 99408
rect 451332 99396 451338 99408
rect 452562 99396 452568 99408
rect 451332 99368 452568 99396
rect 451332 99356 451338 99368
rect 452562 99356 452568 99368
rect 452620 99356 452626 99408
rect 454494 99356 454500 99408
rect 454552 99396 454558 99408
rect 455322 99396 455328 99408
rect 454552 99368 455328 99396
rect 454552 99356 454558 99368
rect 455322 99356 455328 99368
rect 455380 99356 455386 99408
rect 455598 99356 455604 99408
rect 455656 99396 455662 99408
rect 456610 99396 456616 99408
rect 455656 99368 456616 99396
rect 455656 99356 455662 99368
rect 456610 99356 456616 99368
rect 456668 99356 456674 99408
rect 466454 99356 466460 99408
rect 466512 99396 466518 99408
rect 467742 99396 467748 99408
rect 466512 99368 467748 99396
rect 466512 99356 466518 99368
rect 467742 99356 467748 99368
rect 467800 99356 467806 99408
rect 469766 99356 469772 99408
rect 469824 99396 469830 99408
rect 470502 99396 470508 99408
rect 469824 99368 470508 99396
rect 469824 99356 469830 99368
rect 470502 99356 470508 99368
rect 470560 99356 470566 99408
rect 470870 99356 470876 99408
rect 470928 99396 470934 99408
rect 471790 99396 471796 99408
rect 470928 99368 471796 99396
rect 470928 99356 470934 99368
rect 471790 99356 471796 99368
rect 471848 99356 471854 99408
rect 475194 99356 475200 99408
rect 475252 99396 475258 99408
rect 476022 99396 476028 99408
rect 475252 99368 476028 99396
rect 475252 99356 475258 99368
rect 476022 99356 476028 99368
rect 476080 99356 476086 99408
rect 486050 99356 486056 99408
rect 486108 99396 486114 99408
rect 487062 99396 487068 99408
rect 486108 99368 487068 99396
rect 486108 99356 486114 99368
rect 487062 99356 487068 99368
rect 487120 99356 487126 99408
rect 487154 99356 487160 99408
rect 487212 99396 487218 99408
rect 488350 99396 488356 99408
rect 487212 99368 488356 99396
rect 487212 99356 487218 99368
rect 488350 99356 488356 99368
rect 488408 99356 488414 99408
rect 490374 99356 490380 99408
rect 490432 99396 490438 99408
rect 491202 99396 491208 99408
rect 490432 99368 491208 99396
rect 490432 99356 490438 99368
rect 491202 99356 491208 99368
rect 491260 99356 491266 99408
rect 491478 99356 491484 99408
rect 491536 99396 491542 99408
rect 492582 99396 492588 99408
rect 491536 99368 492588 99396
rect 491536 99356 491542 99368
rect 492582 99356 492588 99368
rect 492640 99356 492646 99408
rect 495894 99356 495900 99408
rect 495952 99396 495958 99408
rect 496722 99396 496728 99408
rect 495952 99368 496728 99396
rect 495952 99356 495958 99368
rect 496722 99356 496728 99368
rect 496780 99356 496786 99408
rect 496906 99356 496912 99408
rect 496964 99396 496970 99408
rect 498010 99396 498016 99408
rect 496964 99368 498016 99396
rect 496964 99356 496970 99368
rect 498010 99356 498016 99368
rect 498068 99356 498074 99408
rect 501322 99356 501328 99408
rect 501380 99396 501386 99408
rect 502242 99396 502248 99408
rect 501380 99368 502248 99396
rect 501380 99356 501386 99368
rect 502242 99356 502248 99368
rect 502300 99356 502306 99408
rect 188982 99260 188988 99272
rect 188908 99232 188988 99260
rect 188982 99220 188988 99232
rect 189040 99220 189046 99272
rect 147674 98608 147680 98660
rect 147732 98648 147738 98660
rect 194594 98648 194600 98660
rect 147732 98620 194600 98648
rect 147732 98608 147738 98620
rect 194594 98608 194600 98620
rect 194652 98608 194658 98660
rect 198826 98608 198832 98660
rect 198884 98648 198890 98660
rect 251174 98648 251180 98660
rect 198884 98620 251180 98648
rect 198884 98608 198890 98620
rect 251174 98608 251180 98620
rect 251232 98608 251238 98660
rect 270586 98608 270592 98660
rect 270644 98648 270650 98660
rect 329834 98648 329840 98660
rect 270644 98620 329840 98648
rect 270644 98608 270650 98620
rect 329834 98608 329840 98620
rect 329892 98608 329898 98660
rect 342438 98608 342444 98660
rect 342496 98648 342502 98660
rect 408494 98648 408500 98660
rect 342496 98620 408500 98648
rect 342496 98608 342502 98620
rect 408494 98608 408500 98620
rect 408552 98608 408558 98660
rect 440326 98608 440332 98660
rect 440384 98648 440390 98660
rect 514754 98648 514760 98660
rect 440384 98620 514760 98648
rect 440384 98608 440390 98620
rect 514754 98608 514760 98620
rect 514812 98608 514818 98660
rect 111794 97248 111800 97300
rect 111852 97288 111858 97300
rect 155954 97288 155960 97300
rect 111852 97260 155960 97288
rect 111852 97248 111858 97260
rect 155954 97248 155960 97260
rect 156012 97248 156018 97300
rect 234706 97248 234712 97300
rect 234764 97288 234770 97300
rect 289814 97288 289820 97300
rect 234764 97260 289820 97288
rect 234764 97248 234770 97260
rect 289814 97248 289820 97260
rect 289872 97248 289878 97300
rect 317414 97248 317420 97300
rect 317472 97288 317478 97300
rect 380894 97288 380900 97300
rect 317472 97260 380900 97288
rect 317472 97248 317478 97260
rect 380894 97248 380900 97260
rect 380952 97248 380958 97300
rect 443638 97248 443644 97300
rect 443696 97288 443702 97300
rect 518894 97288 518900 97300
rect 443696 97260 518900 97288
rect 443696 97248 443702 97260
rect 518894 97248 518900 97260
rect 518952 97248 518958 97300
rect 395801 96611 395859 96617
rect 395801 96577 395813 96611
rect 395847 96608 395859 96611
rect 395890 96608 395896 96620
rect 395847 96580 395896 96608
rect 395847 96577 395859 96580
rect 395801 96571 395859 96577
rect 395890 96568 395896 96580
rect 395948 96568 395954 96620
rect 219526 95888 219532 95940
rect 219584 95928 219590 95940
rect 273254 95928 273260 95940
rect 219584 95900 273260 95928
rect 219584 95888 219590 95900
rect 273254 95888 273260 95900
rect 273312 95888 273318 95940
rect 281534 95888 281540 95940
rect 281592 95928 281598 95940
rect 340874 95928 340880 95940
rect 281592 95900 340880 95928
rect 281592 95888 281598 95900
rect 340874 95888 340880 95900
rect 340932 95888 340938 95940
rect 370774 95888 370780 95940
rect 370832 95928 370838 95940
rect 438854 95928 438860 95940
rect 370832 95900 438860 95928
rect 370832 95888 370838 95900
rect 438854 95888 438860 95900
rect 438912 95888 438918 95940
rect 446858 95888 446864 95940
rect 446916 95928 446922 95940
rect 521654 95928 521660 95940
rect 446916 95900 521660 95928
rect 446916 95888 446922 95900
rect 521654 95888 521660 95900
rect 521712 95888 521718 95940
rect 389266 94460 389272 94512
rect 389324 94500 389330 94512
rect 459646 94500 459652 94512
rect 389324 94472 459652 94500
rect 389324 94460 389330 94472
rect 459646 94460 459652 94472
rect 459704 94460 459710 94512
rect 478230 94460 478236 94512
rect 478288 94500 478294 94512
rect 554774 94500 554780 94512
rect 478288 94472 554780 94500
rect 478288 94460 478294 94472
rect 554774 94460 554780 94472
rect 554832 94460 554838 94512
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 79686 93820 79692 93832
rect 3476 93792 79692 93820
rect 3476 93780 3482 93792
rect 79686 93780 79692 93792
rect 79744 93780 79750 93832
rect 368382 93100 368388 93152
rect 368440 93140 368446 93152
rect 434714 93140 434720 93152
rect 368440 93112 434720 93140
rect 368440 93100 368446 93112
rect 434714 93100 434720 93112
rect 434772 93100 434778 93152
rect 480162 93100 480168 93152
rect 480220 93140 480226 93152
rect 557534 93140 557540 93152
rect 480220 93112 557540 93140
rect 480220 93100 480226 93112
rect 557534 93100 557540 93112
rect 557592 93100 557598 93152
rect 354582 91740 354588 91792
rect 354640 91780 354646 91792
rect 420914 91780 420920 91792
rect 354640 91752 420920 91780
rect 354640 91740 354646 91752
rect 420914 91740 420920 91752
rect 420972 91740 420978 91792
rect 435910 91740 435916 91792
rect 435968 91780 435974 91792
rect 509234 91780 509240 91792
rect 435968 91752 509240 91780
rect 435968 91740 435974 91752
rect 509234 91740 509240 91752
rect 509292 91740 509298 91792
rect 364150 90312 364156 90364
rect 364208 90352 364214 90364
rect 430574 90352 430580 90364
rect 364208 90324 430580 90352
rect 364208 90312 364214 90324
rect 430574 90312 430580 90324
rect 430632 90312 430638 90364
rect 441430 90312 441436 90364
rect 441488 90352 441494 90364
rect 516134 90352 516140 90364
rect 441488 90324 516140 90352
rect 441488 90312 441494 90324
rect 516134 90312 516140 90324
rect 516192 90312 516198 90364
rect 148686 89700 148692 89752
rect 148744 89740 148750 89752
rect 148870 89740 148876 89752
rect 148744 89712 148876 89740
rect 148744 89700 148750 89712
rect 148870 89700 148876 89712
rect 148928 89700 148934 89752
rect 225966 89700 225972 89752
rect 226024 89740 226030 89752
rect 226150 89740 226156 89752
rect 226024 89712 226156 89740
rect 226024 89700 226030 89712
rect 226150 89700 226156 89712
rect 226208 89700 226214 89752
rect 235718 89700 235724 89752
rect 235776 89740 235782 89752
rect 235902 89740 235908 89752
rect 235776 89712 235908 89740
rect 235776 89700 235782 89712
rect 235902 89700 235908 89712
rect 235960 89700 235966 89752
rect 297726 89700 297732 89752
rect 297784 89740 297790 89752
rect 297910 89740 297916 89752
rect 297784 89712 297916 89740
rect 297784 89700 297790 89712
rect 297910 89700 297916 89712
rect 297968 89700 297974 89752
rect 462038 89700 462044 89752
rect 462096 89740 462102 89752
rect 462222 89740 462228 89752
rect 462096 89712 462228 89740
rect 462096 89700 462102 89712
rect 462222 89700 462228 89712
rect 462280 89700 462286 89752
rect 419442 88952 419448 89004
rect 419500 88992 419506 89004
rect 491294 88992 491300 89004
rect 419500 88964 491300 88992
rect 419500 88952 419506 88964
rect 491294 88952 491300 88964
rect 491352 88952 491358 89004
rect 498010 88952 498016 89004
rect 498068 88992 498074 89004
rect 574738 88992 574744 89004
rect 498068 88964 574744 88992
rect 498068 88952 498074 88964
rect 574738 88952 574744 88964
rect 574796 88952 574802 89004
rect 504542 88272 504548 88324
rect 504600 88312 504606 88324
rect 580166 88312 580172 88324
rect 504600 88284 580172 88312
rect 504600 88272 504606 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 351822 87592 351828 87644
rect 351880 87632 351886 87644
rect 416774 87632 416780 87644
rect 351880 87604 416780 87632
rect 351880 87592 351886 87604
rect 416774 87592 416780 87604
rect 416832 87592 416838 87644
rect 395798 87020 395804 87032
rect 395759 86992 395804 87020
rect 395798 86980 395804 86992
rect 395856 86980 395862 87032
rect 410978 86980 410984 87032
rect 411036 87020 411042 87032
rect 411070 87020 411076 87032
rect 411036 86992 411076 87020
rect 411036 86980 411042 86992
rect 411070 86980 411076 86992
rect 411128 86980 411134 87032
rect 152829 86955 152887 86961
rect 152829 86921 152841 86955
rect 152875 86952 152887 86955
rect 152918 86952 152924 86964
rect 152875 86924 152924 86952
rect 152875 86921 152887 86924
rect 152829 86915 152887 86921
rect 152918 86912 152924 86924
rect 152976 86912 152982 86964
rect 342162 86232 342168 86284
rect 342220 86272 342226 86284
rect 407114 86272 407120 86284
rect 342220 86244 407120 86272
rect 342220 86232 342226 86244
rect 407114 86232 407120 86244
rect 407172 86232 407178 86284
rect 462958 86232 462964 86284
rect 463016 86272 463022 86284
rect 536834 86272 536840 86284
rect 463016 86244 536840 86272
rect 463016 86232 463022 86244
rect 536834 86232 536840 86244
rect 536892 86232 536898 86284
rect 339310 84804 339316 84856
rect 339368 84844 339374 84856
rect 402974 84844 402980 84856
rect 339368 84816 402980 84844
rect 339368 84804 339374 84816
rect 402974 84804 402980 84816
rect 403032 84804 403038 84856
rect 467558 84804 467564 84856
rect 467616 84844 467622 84856
rect 545114 84844 545120 84856
rect 467616 84816 545120 84844
rect 467616 84804 467622 84816
rect 545114 84804 545120 84816
rect 545172 84804 545178 84856
rect 322750 83444 322756 83496
rect 322808 83484 322814 83496
rect 385034 83484 385040 83496
rect 322808 83456 385040 83484
rect 322808 83444 322814 83456
rect 385034 83444 385040 83456
rect 385092 83444 385098 83496
rect 491202 83444 491208 83496
rect 491260 83484 491266 83496
rect 569954 83484 569960 83496
rect 491260 83456 569960 83484
rect 491260 83444 491266 83456
rect 569954 83444 569960 83456
rect 570012 83444 570018 83496
rect 188706 82084 188712 82136
rect 188764 82124 188770 82136
rect 188890 82124 188896 82136
rect 188764 82096 188896 82124
rect 188764 82084 188770 82096
rect 188890 82084 188896 82096
rect 188948 82084 188954 82136
rect 328362 82084 328368 82136
rect 328420 82124 328426 82136
rect 391934 82124 391940 82136
rect 328420 82096 391940 82124
rect 328420 82084 328426 82096
rect 391934 82084 391940 82096
rect 391992 82084 391998 82136
rect 410978 82124 410984 82136
rect 410939 82096 410984 82124
rect 410978 82084 410984 82096
rect 411036 82084 411042 82136
rect 433242 82084 433248 82136
rect 433300 82124 433306 82136
rect 506474 82124 506480 82136
rect 433300 82096 506480 82124
rect 433300 82084 433306 82096
rect 506474 82084 506480 82096
rect 506532 82084 506538 82136
rect 315942 80724 315948 80776
rect 316000 80764 316006 80776
rect 378226 80764 378232 80776
rect 316000 80736 378232 80764
rect 316000 80724 316006 80736
rect 378226 80724 378232 80736
rect 378284 80724 378290 80776
rect 375190 80656 375196 80708
rect 375248 80696 375254 80708
rect 442994 80696 443000 80708
rect 375248 80668 443000 80696
rect 375248 80656 375254 80668
rect 442994 80656 443000 80668
rect 443052 80656 443058 80708
rect 452470 80656 452476 80708
rect 452528 80696 452534 80708
rect 528554 80696 528560 80708
rect 452528 80668 528560 80696
rect 452528 80656 452534 80668
rect 528554 80656 528560 80668
rect 528612 80656 528618 80708
rect 395798 80112 395804 80164
rect 395856 80112 395862 80164
rect 462130 80112 462136 80164
rect 462188 80112 462194 80164
rect 395816 80028 395844 80112
rect 462148 80028 462176 80112
rect 395798 79976 395804 80028
rect 395856 79976 395862 80028
rect 462130 79976 462136 80028
rect 462188 79976 462194 80028
rect 3510 79432 3516 79484
rect 3568 79472 3574 79484
rect 8938 79472 8944 79484
rect 3568 79444 8944 79472
rect 3568 79432 3574 79444
rect 8938 79432 8944 79444
rect 8996 79432 9002 79484
rect 302050 79364 302056 79416
rect 302108 79404 302114 79416
rect 364334 79404 364340 79416
rect 302108 79376 364340 79404
rect 302108 79364 302114 79376
rect 364334 79364 364340 79376
rect 364392 79364 364398 79416
rect 364242 79296 364248 79348
rect 364300 79336 364306 79348
rect 431954 79336 431960 79348
rect 364300 79308 431960 79336
rect 364300 79296 364306 79308
rect 431954 79296 431960 79308
rect 432012 79296 432018 79348
rect 456610 79296 456616 79348
rect 456668 79336 456674 79348
rect 531314 79336 531320 79348
rect 456668 79308 531320 79336
rect 456668 79296 456674 79308
rect 531314 79296 531320 79308
rect 531372 79296 531378 79348
rect 299382 77936 299388 77988
rect 299440 77976 299446 77988
rect 360194 77976 360200 77988
rect 299440 77948 360200 77976
rect 299440 77936 299446 77948
rect 360194 77936 360200 77948
rect 360252 77936 360258 77988
rect 361482 77936 361488 77988
rect 361540 77976 361546 77988
rect 427814 77976 427820 77988
rect 361540 77948 427820 77976
rect 361540 77936 361546 77948
rect 427814 77936 427820 77948
rect 427872 77936 427878 77988
rect 459462 77936 459468 77988
rect 459520 77976 459526 77988
rect 535454 77976 535460 77988
rect 459520 77948 535460 77976
rect 459520 77936 459526 77948
rect 535454 77936 535460 77948
rect 535512 77936 535518 77988
rect 410978 77364 410984 77376
rect 410939 77336 410984 77364
rect 410978 77324 410984 77336
rect 411036 77324 411042 77376
rect 152826 77296 152832 77308
rect 152787 77268 152832 77296
rect 152826 77256 152832 77268
rect 152884 77256 152890 77308
rect 148873 77231 148931 77237
rect 148873 77197 148885 77231
rect 148919 77228 148931 77231
rect 148962 77228 148968 77240
rect 148919 77200 148968 77228
rect 148919 77197 148931 77200
rect 148873 77191 148931 77197
rect 148962 77188 148968 77200
rect 149020 77188 149026 77240
rect 188525 77231 188583 77237
rect 188525 77197 188537 77231
rect 188571 77228 188583 77231
rect 188614 77228 188620 77240
rect 188571 77200 188620 77228
rect 188571 77197 188583 77200
rect 188525 77191 188583 77197
rect 188614 77188 188620 77200
rect 188672 77188 188678 77240
rect 225877 77231 225935 77237
rect 225877 77197 225889 77231
rect 225923 77228 225935 77231
rect 225966 77228 225972 77240
rect 225923 77200 225972 77228
rect 225923 77197 225935 77200
rect 225877 77191 225935 77197
rect 225966 77188 225972 77200
rect 226024 77188 226030 77240
rect 235629 77231 235687 77237
rect 235629 77197 235641 77231
rect 235675 77228 235687 77231
rect 235718 77228 235724 77240
rect 235675 77200 235724 77228
rect 235675 77197 235687 77200
rect 235629 77191 235687 77197
rect 235718 77188 235724 77200
rect 235776 77188 235782 77240
rect 297726 77228 297732 77240
rect 297687 77200 297732 77228
rect 297726 77188 297732 77200
rect 297784 77188 297790 77240
rect 378134 77228 378140 77240
rect 378095 77200 378140 77228
rect 378134 77188 378140 77200
rect 378192 77188 378198 77240
rect 504634 77188 504640 77240
rect 504692 77228 504698 77240
rect 580166 77228 580172 77240
rect 504692 77200 580172 77228
rect 504692 77188 504698 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 296622 76508 296628 76560
rect 296680 76548 296686 76560
rect 356054 76548 356060 76560
rect 296680 76520 356060 76548
rect 296680 76508 296686 76520
rect 356054 76508 356060 76520
rect 356112 76508 356118 76560
rect 358630 76508 358636 76560
rect 358688 76548 358694 76560
rect 425054 76548 425060 76560
rect 358688 76520 425060 76548
rect 358688 76508 358694 76520
rect 425054 76508 425060 76520
rect 425112 76508 425118 76560
rect 430482 76508 430488 76560
rect 430540 76548 430546 76560
rect 502334 76548 502340 76560
rect 430540 76520 502340 76548
rect 430540 76508 430546 76520
rect 502334 76508 502340 76520
rect 502392 76508 502398 76560
rect 260742 75148 260748 75200
rect 260800 75188 260806 75200
rect 317414 75188 317420 75200
rect 260800 75160 317420 75188
rect 260800 75148 260806 75160
rect 317414 75148 317420 75160
rect 317472 75148 317478 75200
rect 318702 75148 318708 75200
rect 318760 75188 318766 75200
rect 382274 75188 382280 75200
rect 318760 75160 382280 75188
rect 318760 75148 318766 75160
rect 382274 75148 382280 75160
rect 382332 75148 382338 75200
rect 426342 75148 426348 75200
rect 426400 75188 426406 75200
rect 499574 75188 499580 75200
rect 426400 75160 499580 75188
rect 426400 75148 426406 75160
rect 499574 75148 499580 75160
rect 499632 75148 499638 75200
rect 256510 73856 256516 73908
rect 256568 73896 256574 73908
rect 313274 73896 313280 73908
rect 256568 73868 313280 73896
rect 256568 73856 256574 73868
rect 313274 73856 313280 73868
rect 313332 73856 313338 73908
rect 313090 73788 313096 73840
rect 313148 73828 313154 73840
rect 373994 73828 374000 73840
rect 313148 73800 374000 73828
rect 313148 73788 313154 73800
rect 373994 73788 374000 73800
rect 374052 73788 374058 73840
rect 423582 73788 423588 73840
rect 423640 73828 423646 73840
rect 495434 73828 495440 73840
rect 423640 73800 495440 73828
rect 423640 73788 423646 73800
rect 495434 73788 495440 73800
rect 495492 73788 495498 73840
rect 246942 72428 246948 72480
rect 247000 72468 247006 72480
rect 303614 72468 303620 72480
rect 247000 72440 303620 72468
rect 247000 72428 247006 72440
rect 303614 72428 303620 72440
rect 303672 72428 303678 72480
rect 309042 72428 309048 72480
rect 309100 72468 309106 72480
rect 371234 72468 371240 72480
rect 309100 72440 371240 72468
rect 309100 72428 309106 72440
rect 371234 72428 371240 72440
rect 371292 72428 371298 72480
rect 420730 72428 420736 72480
rect 420788 72468 420794 72480
rect 492674 72468 492680 72480
rect 420788 72440 492680 72468
rect 420788 72428 420794 72440
rect 492674 72428 492680 72440
rect 492732 72428 492738 72480
rect 280062 71068 280068 71120
rect 280120 71108 280126 71120
rect 339494 71108 339500 71120
rect 280120 71080 339500 71108
rect 280120 71068 280126 71080
rect 339494 71068 339500 71080
rect 339552 71068 339558 71120
rect 224862 71000 224868 71052
rect 224920 71040 224926 71052
rect 278774 71040 278780 71052
rect 224920 71012 278780 71040
rect 224920 71000 224926 71012
rect 278774 71000 278780 71012
rect 278832 71000 278838 71052
rect 335262 71000 335268 71052
rect 335320 71040 335326 71052
rect 400214 71040 400220 71052
rect 335320 71012 400220 71040
rect 335320 71000 335326 71012
rect 400214 71000 400220 71012
rect 400272 71000 400278 71052
rect 409782 71000 409788 71052
rect 409840 71040 409846 71052
rect 480254 71040 480260 71052
rect 409840 71012 480260 71040
rect 409840 71000 409846 71012
rect 480254 71000 480260 71012
rect 480312 71000 480318 71052
rect 153010 70428 153016 70440
rect 152936 70400 153016 70428
rect 152936 70304 152964 70400
rect 153010 70388 153016 70400
rect 153068 70388 153074 70440
rect 410886 70388 410892 70440
rect 410944 70388 410950 70440
rect 152918 70252 152924 70304
rect 152976 70252 152982 70304
rect 410904 70292 410932 70388
rect 410978 70292 410984 70304
rect 410904 70264 410984 70292
rect 410978 70252 410984 70264
rect 411036 70252 411042 70304
rect 230290 69640 230296 69692
rect 230348 69680 230354 69692
rect 285674 69680 285680 69692
rect 230348 69652 285680 69680
rect 230348 69640 230354 69652
rect 285674 69640 285680 69652
rect 285732 69640 285738 69692
rect 286962 69640 286968 69692
rect 287020 69680 287026 69692
rect 346394 69680 346400 69692
rect 287020 69652 346400 69680
rect 287020 69640 287026 69652
rect 346394 69640 346400 69652
rect 346452 69640 346458 69692
rect 405550 69640 405556 69692
rect 405608 69680 405614 69692
rect 477586 69680 477592 69692
rect 405608 69652 477592 69680
rect 405608 69640 405614 69652
rect 477586 69640 477592 69652
rect 477644 69640 477650 69692
rect 215110 68280 215116 68332
rect 215168 68320 215174 68332
rect 267734 68320 267740 68332
rect 215168 68292 267740 68320
rect 215168 68280 215174 68292
rect 267734 68280 267740 68292
rect 267792 68280 267798 68332
rect 273162 68280 273168 68332
rect 273220 68320 273226 68332
rect 331214 68320 331220 68332
rect 273220 68292 331220 68320
rect 273220 68280 273226 68292
rect 331214 68280 331220 68292
rect 331272 68280 331278 68332
rect 332502 68280 332508 68332
rect 332560 68320 332566 68332
rect 396074 68320 396080 68332
rect 332560 68292 396080 68320
rect 332560 68280 332566 68292
rect 396074 68280 396080 68292
rect 396132 68280 396138 68332
rect 402882 68280 402888 68332
rect 402940 68320 402946 68332
rect 473354 68320 473360 68332
rect 402940 68292 473360 68320
rect 402940 68280 402946 68292
rect 473354 68280 473360 68292
rect 473412 68280 473418 68332
rect 378134 67708 378140 67720
rect 378095 67680 378140 67708
rect 378134 67668 378140 67680
rect 378192 67668 378198 67720
rect 148870 67640 148876 67652
rect 148831 67612 148876 67640
rect 148870 67600 148876 67612
rect 148928 67600 148934 67652
rect 188522 67640 188528 67652
rect 188483 67612 188528 67640
rect 188522 67600 188528 67612
rect 188580 67600 188586 67652
rect 225874 67640 225880 67652
rect 225835 67612 225880 67640
rect 225874 67600 225880 67612
rect 225932 67600 225938 67652
rect 235626 67640 235632 67652
rect 235587 67612 235632 67640
rect 235626 67600 235632 67612
rect 235684 67600 235690 67652
rect 297729 67643 297787 67649
rect 297729 67609 297741 67643
rect 297775 67640 297787 67643
rect 297818 67640 297824 67652
rect 297775 67612 297824 67640
rect 297775 67609 297787 67612
rect 297729 67603 297787 67609
rect 297818 67600 297824 67612
rect 297876 67600 297882 67652
rect 378134 67572 378140 67584
rect 378095 67544 378140 67572
rect 378134 67532 378140 67544
rect 378192 67532 378198 67584
rect 499574 67572 499580 67584
rect 499535 67544 499580 67572
rect 499574 67532 499580 67544
rect 499632 67532 499638 67584
rect 237282 66920 237288 66972
rect 237340 66960 237346 66972
rect 292574 66960 292580 66972
rect 237340 66932 292580 66960
rect 237340 66920 237346 66932
rect 292574 66920 292580 66932
rect 292632 66920 292638 66972
rect 395798 66920 395804 66972
rect 395856 66960 395862 66972
rect 466454 66960 466460 66972
rect 395856 66932 466460 66960
rect 395856 66920 395862 66932
rect 466454 66920 466460 66932
rect 466512 66920 466518 66972
rect 184842 66852 184848 66904
rect 184900 66892 184906 66904
rect 235994 66892 236000 66904
rect 184900 66864 236000 66892
rect 184900 66852 184906 66864
rect 235994 66852 236000 66864
rect 236052 66852 236058 66904
rect 292390 66852 292396 66904
rect 292448 66892 292454 66904
rect 353386 66892 353392 66904
rect 292448 66864 353392 66892
rect 292448 66852 292454 66864
rect 353386 66852 353392 66864
rect 353444 66852 353450 66904
rect 466362 66852 466368 66904
rect 466420 66892 466426 66904
rect 542354 66892 542360 66904
rect 466420 66864 542360 66892
rect 466420 66852 466426 66864
rect 542354 66852 542360 66864
rect 542412 66852 542418 66904
rect 371234 66212 371240 66224
rect 371195 66184 371240 66212
rect 371234 66172 371240 66184
rect 371292 66172 371298 66224
rect 393222 65560 393228 65612
rect 393280 65600 393286 65612
rect 462314 65600 462320 65612
rect 393280 65572 462320 65600
rect 393280 65560 393286 65572
rect 462314 65560 462320 65572
rect 462372 65560 462378 65612
rect 182082 65492 182088 65544
rect 182140 65532 182146 65544
rect 231854 65532 231860 65544
rect 182140 65504 231860 65532
rect 182140 65492 182146 65504
rect 231854 65492 231860 65504
rect 231912 65492 231918 65544
rect 234522 65492 234528 65544
rect 234580 65532 234586 65544
rect 288434 65532 288440 65544
rect 234580 65504 288440 65532
rect 234580 65492 234586 65504
rect 288434 65492 288440 65504
rect 288492 65492 288498 65544
rect 289722 65492 289728 65544
rect 289780 65532 289786 65544
rect 349154 65532 349160 65544
rect 289780 65504 349160 65532
rect 289780 65492 289786 65504
rect 349154 65492 349160 65504
rect 349212 65492 349218 65544
rect 462038 65492 462044 65544
rect 462096 65532 462102 65544
rect 538214 65532 538220 65544
rect 462096 65504 538220 65532
rect 462096 65492 462102 65504
rect 538214 65492 538220 65504
rect 538272 65492 538278 65544
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 79594 64852 79600 64864
rect 3384 64824 79600 64852
rect 3384 64812 3390 64824
rect 79594 64812 79600 64824
rect 79652 64812 79658 64864
rect 527818 64812 527824 64864
rect 527876 64852 527882 64864
rect 579798 64852 579804 64864
rect 527876 64824 579804 64852
rect 527876 64812 527882 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 179230 64200 179236 64252
rect 179288 64240 179294 64252
rect 227714 64240 227720 64252
rect 179288 64212 227720 64240
rect 179288 64200 179294 64212
rect 227714 64200 227720 64212
rect 227772 64200 227778 64252
rect 227622 64132 227628 64184
rect 227680 64172 227686 64184
rect 281534 64172 281540 64184
rect 227680 64144 281540 64172
rect 227680 64132 227686 64144
rect 281534 64132 281540 64144
rect 281592 64132 281598 64184
rect 282822 64132 282828 64184
rect 282880 64172 282886 64184
rect 342254 64172 342260 64184
rect 282880 64144 342260 64172
rect 282880 64132 282886 64144
rect 342254 64132 342260 64144
rect 342312 64132 342318 64184
rect 383562 64132 383568 64184
rect 383620 64172 383626 64184
rect 451274 64172 451280 64184
rect 383620 64144 451280 64172
rect 383620 64132 383626 64144
rect 451274 64132 451280 64144
rect 451332 64132 451338 64184
rect 452562 64132 452568 64184
rect 452620 64172 452626 64184
rect 527174 64172 527180 64184
rect 452620 64144 527180 64172
rect 452620 64132 452626 64144
rect 527174 64132 527180 64144
rect 527232 64132 527238 64184
rect 172422 62772 172428 62824
rect 172480 62812 172486 62824
rect 220814 62812 220820 62824
rect 172480 62784 220820 62812
rect 172480 62772 172486 62784
rect 220814 62772 220820 62784
rect 220872 62772 220878 62824
rect 221458 62772 221464 62824
rect 221516 62812 221522 62824
rect 274634 62812 274640 62824
rect 221516 62784 274640 62812
rect 221516 62772 221522 62784
rect 274634 62772 274640 62784
rect 274692 62772 274698 62824
rect 277210 62772 277216 62824
rect 277268 62812 277274 62824
rect 335354 62812 335360 62824
rect 277268 62784 335360 62812
rect 277268 62772 277274 62784
rect 335354 62772 335360 62784
rect 335412 62772 335418 62824
rect 376662 62772 376668 62824
rect 376720 62812 376726 62824
rect 444374 62812 444380 62824
rect 376720 62784 444380 62812
rect 376720 62772 376726 62784
rect 444374 62772 444380 62784
rect 444432 62772 444438 62824
rect 447042 62772 447048 62824
rect 447100 62812 447106 62824
rect 520274 62812 520280 62824
rect 447100 62784 520280 62812
rect 447100 62772 447106 62784
rect 520274 62772 520280 62784
rect 520332 62772 520338 62824
rect 211062 61412 211068 61464
rect 211120 61452 211126 61464
rect 263594 61452 263600 61464
rect 211120 61424 263600 61452
rect 211120 61412 211126 61424
rect 263594 61412 263600 61424
rect 263652 61412 263658 61464
rect 410702 61412 410708 61464
rect 410760 61452 410766 61464
rect 410978 61452 410984 61464
rect 410760 61424 410984 61452
rect 410760 61412 410766 61424
rect 410978 61412 410984 61424
rect 411036 61412 411042 61464
rect 158530 61344 158536 61396
rect 158588 61384 158594 61396
rect 207014 61384 207020 61396
rect 158588 61356 207020 61384
rect 158588 61344 158594 61356
rect 207014 61344 207020 61356
rect 207072 61344 207078 61396
rect 263502 61344 263508 61396
rect 263560 61384 263566 61396
rect 321554 61384 321560 61396
rect 263560 61356 321560 61384
rect 263560 61344 263566 61356
rect 321554 61344 321560 61356
rect 321612 61344 321618 61396
rect 347682 61344 347688 61396
rect 347740 61384 347746 61396
rect 412634 61384 412640 61396
rect 347740 61356 412640 61384
rect 347740 61344 347746 61356
rect 412634 61344 412640 61356
rect 412692 61344 412698 61396
rect 413922 61344 413928 61396
rect 413980 61384 413986 61396
rect 485774 61384 485780 61396
rect 413980 61356 485780 61384
rect 413980 61344 413986 61356
rect 485774 61344 485780 61356
rect 485832 61344 485838 61396
rect 148870 60840 148876 60852
rect 148796 60812 148876 60840
rect 148796 60716 148824 60812
rect 148870 60800 148876 60812
rect 148928 60800 148934 60852
rect 297818 60840 297824 60852
rect 297744 60812 297824 60840
rect 297744 60716 297772 60812
rect 297818 60800 297824 60812
rect 297876 60800 297882 60852
rect 148778 60664 148784 60716
rect 148836 60664 148842 60716
rect 297726 60664 297732 60716
rect 297784 60664 297790 60716
rect 217962 60052 217968 60104
rect 218020 60092 218026 60104
rect 270494 60092 270500 60104
rect 218020 60064 270500 60092
rect 218020 60052 218026 60064
rect 270494 60052 270500 60064
rect 270552 60052 270558 60104
rect 169570 59984 169576 60036
rect 169628 60024 169634 60036
rect 218054 60024 218060 60036
rect 169628 59996 218060 60024
rect 169628 59984 169634 59996
rect 218054 59984 218060 59996
rect 218112 59984 218118 60036
rect 270402 59984 270408 60036
rect 270460 60024 270466 60036
rect 328454 60024 328460 60036
rect 270460 59996 328460 60024
rect 270460 59984 270466 59996
rect 328454 59984 328460 59996
rect 328512 59984 328518 60036
rect 369670 59984 369676 60036
rect 369728 60024 369734 60036
rect 437474 60024 437480 60036
rect 369728 59996 437480 60024
rect 369728 59984 369734 59996
rect 437474 59984 437480 59996
rect 437532 59984 437538 60036
rect 440142 59984 440148 60036
rect 440200 60024 440206 60036
rect 513374 60024 513380 60036
rect 440200 59996 513380 60024
rect 440200 59984 440206 59996
rect 513374 59984 513380 59996
rect 513432 59984 513438 60036
rect 155862 58624 155868 58676
rect 155920 58664 155926 58676
rect 202874 58664 202880 58676
rect 155920 58636 202880 58664
rect 155920 58624 155926 58636
rect 202874 58624 202880 58636
rect 202932 58624 202938 58676
rect 208302 58624 208308 58676
rect 208360 58664 208366 58676
rect 260834 58664 260840 58676
rect 208360 58636 260840 58664
rect 208360 58624 208366 58636
rect 260834 58624 260840 58636
rect 260892 58624 260898 58676
rect 314562 58624 314568 58676
rect 314620 58664 314626 58676
rect 376754 58664 376760 58676
rect 314620 58636 376760 58664
rect 314620 58624 314626 58636
rect 376754 58624 376760 58636
rect 376812 58624 376818 58676
rect 379422 58624 379428 58676
rect 379480 58664 379486 58676
rect 448514 58664 448520 58676
rect 379480 58636 448520 58664
rect 379480 58624 379486 58636
rect 448514 58624 448520 58636
rect 448572 58624 448578 58676
rect 449802 58624 449808 58676
rect 449860 58664 449866 58676
rect 524414 58664 524420 58676
rect 449860 58636 524420 58664
rect 449860 58624 449866 58636
rect 524414 58624 524420 58636
rect 524472 58624 524478 58676
rect 333698 57944 333704 57996
rect 333756 57984 333762 57996
rect 333790 57984 333796 57996
rect 333756 57956 333796 57984
rect 333756 57944 333762 57956
rect 333790 57944 333796 57956
rect 333848 57944 333854 57996
rect 378134 57984 378140 57996
rect 378095 57956 378140 57984
rect 378134 57944 378140 57956
rect 378192 57944 378198 57996
rect 499574 57984 499580 57996
rect 499535 57956 499580 57984
rect 499574 57944 499580 57956
rect 499632 57944 499638 57996
rect 353294 57916 353300 57928
rect 353255 57888 353300 57916
rect 353294 57876 353300 57888
rect 353352 57876 353358 57928
rect 495434 57916 495440 57928
rect 495395 57888 495440 57916
rect 495434 57876 495440 57888
rect 495492 57876 495498 57928
rect 378134 57848 378140 57860
rect 378095 57820 378140 57848
rect 378134 57808 378140 57820
rect 378192 57808 378198 57860
rect 205450 57264 205456 57316
rect 205508 57304 205514 57316
rect 256694 57304 256700 57316
rect 205508 57276 256700 57304
rect 205508 57264 205514 57276
rect 256694 57264 256700 57276
rect 256752 57264 256758 57316
rect 306282 57264 306288 57316
rect 306340 57304 306346 57316
rect 367094 57304 367100 57316
rect 306340 57276 367100 57304
rect 306340 57264 306346 57276
rect 367094 57264 367100 57276
rect 367152 57264 367158 57316
rect 152918 57196 152924 57248
rect 152976 57236 152982 57248
rect 200114 57236 200120 57248
rect 152976 57208 200120 57236
rect 152976 57196 152982 57208
rect 200114 57196 200120 57208
rect 200172 57196 200178 57248
rect 253842 57196 253848 57248
rect 253900 57236 253906 57248
rect 310514 57236 310520 57248
rect 253900 57208 310520 57236
rect 253900 57196 253906 57208
rect 310514 57196 310520 57208
rect 310572 57196 310578 57248
rect 367002 57196 367008 57248
rect 367060 57236 367066 57248
rect 433334 57236 433340 57248
rect 367060 57208 433340 57236
rect 367060 57196 367066 57208
rect 433334 57196 433340 57208
rect 433392 57196 433398 57248
rect 436002 57196 436008 57248
rect 436060 57236 436066 57248
rect 510614 57236 510620 57248
rect 436060 57208 510620 57236
rect 436060 57196 436066 57208
rect 510614 57196 510620 57208
rect 510672 57196 510678 57248
rect 371234 56624 371240 56636
rect 371195 56596 371240 56624
rect 371234 56584 371240 56596
rect 371292 56584 371298 56636
rect 410702 56556 410708 56568
rect 410663 56528 410708 56556
rect 410702 56516 410708 56528
rect 410760 56516 410766 56568
rect 201402 55904 201408 55956
rect 201460 55944 201466 55956
rect 252554 55944 252560 55956
rect 201460 55916 252560 55944
rect 201460 55904 201466 55916
rect 252554 55904 252560 55916
rect 252612 55904 252618 55956
rect 148778 55836 148784 55888
rect 148836 55876 148842 55888
rect 195974 55876 195980 55888
rect 148836 55848 195980 55876
rect 148836 55836 148842 55848
rect 195974 55836 195980 55848
rect 196032 55836 196038 55888
rect 250990 55836 250996 55888
rect 251048 55876 251054 55888
rect 306374 55876 306380 55888
rect 251048 55848 306380 55876
rect 251048 55836 251054 55848
rect 306374 55836 306380 55848
rect 306432 55836 306438 55888
rect 307662 55836 307668 55888
rect 307720 55876 307726 55888
rect 369854 55876 369860 55888
rect 307720 55848 369860 55876
rect 307720 55836 307726 55848
rect 369854 55836 369860 55848
rect 369912 55836 369918 55888
rect 373902 55836 373908 55888
rect 373960 55876 373966 55888
rect 441614 55876 441620 55888
rect 373960 55848 441620 55876
rect 373960 55836 373966 55848
rect 441614 55836 441620 55848
rect 441672 55836 441678 55888
rect 442902 55836 442908 55888
rect 442960 55876 442966 55888
rect 517514 55876 517520 55888
rect 442960 55848 517520 55876
rect 442960 55836 442966 55848
rect 517514 55836 517520 55848
rect 517572 55836 517578 55888
rect 194410 54544 194416 54596
rect 194468 54584 194474 54596
rect 245654 54584 245660 54596
rect 194468 54556 245660 54584
rect 194468 54544 194474 54556
rect 245654 54544 245660 54556
rect 245712 54544 245718 54596
rect 350442 54544 350448 54596
rect 350500 54584 350506 54596
rect 416866 54584 416872 54596
rect 350500 54556 416872 54584
rect 350500 54544 350506 54556
rect 416866 54544 416872 54556
rect 416924 54544 416930 54596
rect 146202 54476 146208 54528
rect 146260 54516 146266 54528
rect 193214 54516 193220 54528
rect 146260 54488 193220 54516
rect 146260 54476 146266 54488
rect 193214 54476 193220 54488
rect 193272 54476 193278 54528
rect 244182 54476 244188 54528
rect 244240 54516 244246 54528
rect 299474 54516 299480 54528
rect 244240 54488 299480 54516
rect 244240 54476 244246 54488
rect 299474 54476 299480 54488
rect 299532 54476 299538 54528
rect 416682 54476 416688 54528
rect 416740 54516 416746 54528
rect 488534 54516 488540 54528
rect 416740 54488 488540 54516
rect 416740 54476 416746 54488
rect 488534 54476 488540 54488
rect 488592 54476 488598 54528
rect 191742 53116 191748 53168
rect 191800 53156 191806 53168
rect 242894 53156 242900 53168
rect 191800 53128 242900 53156
rect 191800 53116 191806 53128
rect 242894 53116 242900 53128
rect 242952 53116 242958 53168
rect 143350 53048 143356 53100
rect 143408 53088 143414 53100
rect 189074 53088 189080 53100
rect 143408 53060 189080 53088
rect 143408 53048 143414 53060
rect 189074 53048 189080 53060
rect 189132 53048 189138 53100
rect 241330 53048 241336 53100
rect 241388 53088 241394 53100
rect 296714 53088 296720 53100
rect 241388 53060 296720 53088
rect 241388 53048 241394 53060
rect 296714 53048 296720 53060
rect 296772 53048 296778 53100
rect 297726 53048 297732 53100
rect 297784 53088 297790 53100
rect 358814 53088 358820 53100
rect 297784 53060 358820 53088
rect 297784 53048 297790 53060
rect 358814 53048 358820 53060
rect 358872 53048 358878 53100
rect 360102 53048 360108 53100
rect 360160 53088 360166 53100
rect 426434 53088 426440 53100
rect 360160 53060 426440 53088
rect 360160 53048 360166 53060
rect 426434 53048 426440 53060
rect 426492 53048 426498 53100
rect 458082 53048 458088 53100
rect 458140 53088 458146 53100
rect 534074 53088 534080 53100
rect 458140 53060 534080 53088
rect 458140 53048 458146 53060
rect 534074 53048 534080 53060
rect 534132 53048 534138 53100
rect 139302 51688 139308 51740
rect 139360 51728 139366 51740
rect 184934 51728 184940 51740
rect 139360 51700 184940 51728
rect 139360 51688 139366 51700
rect 184934 51688 184940 51700
rect 184992 51688 184998 51740
rect 188706 51688 188712 51740
rect 188764 51728 188770 51740
rect 238754 51728 238760 51740
rect 188764 51700 238760 51728
rect 188764 51688 188770 51700
rect 238754 51688 238760 51700
rect 238812 51688 238818 51740
rect 242802 51688 242808 51740
rect 242860 51728 242866 51740
rect 298094 51728 298100 51740
rect 242860 51700 298100 51728
rect 242860 51688 242866 51700
rect 298094 51688 298100 51700
rect 298152 51688 298158 51740
rect 340782 51688 340788 51740
rect 340840 51728 340846 51740
rect 405734 51728 405740 51740
rect 340840 51700 405740 51728
rect 340840 51688 340846 51700
rect 405734 51688 405740 51700
rect 405792 51688 405798 51740
rect 455322 51688 455328 51740
rect 455380 51728 455386 51740
rect 529934 51728 529940 51740
rect 455380 51700 529940 51728
rect 455380 51688 455386 51700
rect 529934 51688 529940 51700
rect 529992 51688 529998 51740
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 79502 51048 79508 51060
rect 3476 51020 79508 51048
rect 3476 51008 3482 51020
rect 79502 51008 79508 51020
rect 79560 51008 79566 51060
rect 410705 50983 410763 50989
rect 410705 50949 410717 50983
rect 410751 50980 410763 50983
rect 410978 50980 410984 50992
rect 410751 50952 410984 50980
rect 410751 50949 410763 50952
rect 410705 50943 410763 50949
rect 410978 50940 410984 50952
rect 411036 50940 411042 50992
rect 235810 50436 235816 50448
rect 235771 50408 235816 50436
rect 235810 50396 235816 50408
rect 235868 50396 235874 50448
rect 136542 50328 136548 50380
rect 136600 50368 136606 50380
rect 182174 50368 182180 50380
rect 136600 50340 182180 50368
rect 136600 50328 136606 50340
rect 182174 50328 182180 50340
rect 182232 50328 182238 50380
rect 209590 50328 209596 50380
rect 209648 50368 209654 50380
rect 262214 50368 262220 50380
rect 209648 50340 262220 50368
rect 209648 50328 209654 50340
rect 262214 50328 262220 50340
rect 262272 50328 262278 50380
rect 275922 50328 275928 50380
rect 275980 50368 275986 50380
rect 333974 50368 333980 50380
rect 275980 50340 333980 50368
rect 275980 50328 275986 50340
rect 333974 50328 333980 50340
rect 334032 50328 334038 50380
rect 338022 50328 338028 50380
rect 338080 50368 338086 50380
rect 401594 50368 401600 50380
rect 338080 50340 401600 50368
rect 338080 50328 338086 50340
rect 401594 50328 401600 50340
rect 401652 50328 401658 50380
rect 431862 50328 431868 50380
rect 431920 50368 431926 50380
rect 505094 50368 505100 50380
rect 431920 50340 505100 50368
rect 431920 50328 431926 50340
rect 505094 50328 505100 50340
rect 505152 50328 505158 50380
rect 133690 49036 133696 49088
rect 133748 49076 133754 49088
rect 178034 49076 178040 49088
rect 133748 49048 178040 49076
rect 133748 49036 133754 49048
rect 178034 49036 178040 49048
rect 178092 49036 178098 49088
rect 175182 48968 175188 49020
rect 175240 49008 175246 49020
rect 224954 49008 224960 49020
rect 175240 48980 224960 49008
rect 175240 48968 175246 48980
rect 224954 48968 224960 48980
rect 225012 48968 225018 49020
rect 225966 48968 225972 49020
rect 226024 49008 226030 49020
rect 280154 49008 280160 49020
rect 226024 48980 280160 49008
rect 226024 48968 226030 48980
rect 280154 48968 280160 48980
rect 280212 48968 280218 49020
rect 292482 48968 292488 49020
rect 292540 49008 292546 49020
rect 351914 49008 351920 49020
rect 292540 48980 351920 49008
rect 292540 48968 292546 48980
rect 351914 48968 351920 48980
rect 351972 48968 351978 49020
rect 357342 48968 357348 49020
rect 357400 49008 357406 49020
rect 423674 49008 423680 49020
rect 357400 48980 423680 49008
rect 357400 48968 357406 48980
rect 423674 48968 423680 48980
rect 423732 48968 423738 49020
rect 427078 48968 427084 49020
rect 427136 49008 427142 49020
rect 498194 49008 498200 49020
rect 427136 48980 498200 49008
rect 427136 48968 427142 48980
rect 498194 48968 498200 48980
rect 498252 48968 498258 49020
rect 353294 48328 353300 48340
rect 353255 48300 353300 48328
rect 353294 48288 353300 48300
rect 353352 48288 353358 48340
rect 378134 48328 378140 48340
rect 378095 48300 378140 48328
rect 378134 48288 378140 48300
rect 378192 48288 378198 48340
rect 495434 48328 495440 48340
rect 495395 48300 495440 48328
rect 495434 48288 495440 48300
rect 495492 48288 495498 48340
rect 333790 48192 333796 48204
rect 333751 48164 333796 48192
rect 333790 48152 333796 48164
rect 333848 48152 333854 48204
rect 164142 47540 164148 47592
rect 164200 47580 164206 47592
rect 212534 47580 212540 47592
rect 164200 47552 212540 47580
rect 164200 47540 164206 47552
rect 212534 47540 212540 47552
rect 212592 47540 212598 47592
rect 213822 47540 213828 47592
rect 213880 47580 213886 47592
rect 266354 47580 266360 47592
rect 213880 47552 266360 47580
rect 213880 47540 213886 47552
rect 266354 47540 266360 47552
rect 266412 47540 266418 47592
rect 271690 47540 271696 47592
rect 271748 47580 271754 47592
rect 331306 47580 331312 47592
rect 271748 47552 331312 47580
rect 271748 47540 271754 47552
rect 331306 47540 331312 47552
rect 331364 47540 331370 47592
rect 333793 47583 333851 47589
rect 333793 47549 333805 47583
rect 333839 47580 333851 47583
rect 398834 47580 398840 47592
rect 333839 47552 398840 47580
rect 333839 47549 333851 47552
rect 333793 47543 333851 47549
rect 398834 47540 398840 47552
rect 398892 47540 398898 47592
rect 400030 47540 400036 47592
rect 400088 47580 400094 47592
rect 469214 47580 469220 47592
rect 400088 47552 469220 47580
rect 400088 47540 400094 47552
rect 469214 47540 469220 47552
rect 469272 47540 469278 47592
rect 473262 47540 473268 47592
rect 473320 47580 473326 47592
rect 550634 47580 550640 47592
rect 473320 47552 550640 47580
rect 473320 47540 473326 47552
rect 550634 47540 550640 47552
rect 550692 47540 550698 47592
rect 371234 46900 371240 46912
rect 371195 46872 371240 46900
rect 371234 46860 371240 46872
rect 371292 46860 371298 46912
rect 129642 46180 129648 46232
rect 129700 46220 129706 46232
rect 175274 46220 175280 46232
rect 129700 46192 175280 46220
rect 129700 46180 129706 46192
rect 175274 46180 175280 46192
rect 175332 46180 175338 46232
rect 197262 46180 197268 46232
rect 197320 46220 197326 46232
rect 248414 46220 248420 46232
rect 197320 46192 248420 46220
rect 197320 46180 197326 46192
rect 248414 46180 248420 46192
rect 248472 46180 248478 46232
rect 269022 46180 269028 46232
rect 269080 46220 269086 46232
rect 327074 46220 327080 46232
rect 269080 46192 327080 46220
rect 269080 46180 269086 46192
rect 327074 46180 327080 46192
rect 327132 46180 327138 46232
rect 329098 46180 329104 46232
rect 329156 46220 329162 46232
rect 390554 46220 390560 46232
rect 329156 46192 390560 46220
rect 329156 46180 329162 46192
rect 390554 46180 390560 46192
rect 390612 46180 390618 46232
rect 429102 46180 429108 46232
rect 429160 46220 429166 46232
rect 502426 46220 502432 46232
rect 429160 46192 502432 46220
rect 429160 46180 429166 46192
rect 502426 46180 502432 46192
rect 502484 46180 502490 46232
rect 235813 45611 235871 45617
rect 235813 45577 235825 45611
rect 235859 45608 235871 45611
rect 235902 45608 235908 45620
rect 235859 45580 235908 45608
rect 235859 45577 235871 45580
rect 235813 45571 235871 45577
rect 235902 45568 235908 45580
rect 235960 45568 235966 45620
rect 169662 44820 169668 44872
rect 169720 44860 169726 44872
rect 218146 44860 218152 44872
rect 169720 44832 218152 44860
rect 169720 44820 169726 44832
rect 218146 44820 218152 44832
rect 218204 44820 218210 44872
rect 262030 44820 262036 44872
rect 262088 44860 262094 44872
rect 318794 44860 318800 44872
rect 262088 44832 318800 44860
rect 262088 44820 262094 44832
rect 318794 44820 318800 44832
rect 318852 44820 318858 44872
rect 324222 44820 324228 44872
rect 324280 44860 324286 44872
rect 387794 44860 387800 44872
rect 324280 44832 387800 44860
rect 324280 44820 324286 44832
rect 387794 44820 387800 44832
rect 387852 44820 387858 44872
rect 422202 44820 422208 44872
rect 422260 44860 422266 44872
rect 494054 44860 494060 44872
rect 422260 44832 494060 44860
rect 422260 44820 422266 44832
rect 494054 44820 494060 44832
rect 494112 44820 494118 44872
rect 126882 43392 126888 43444
rect 126940 43432 126946 43444
rect 171134 43432 171140 43444
rect 126940 43404 171140 43432
rect 126940 43392 126946 43404
rect 171134 43392 171140 43404
rect 171192 43392 171198 43444
rect 194502 43392 194508 43444
rect 194560 43432 194566 43444
rect 244274 43432 244280 43444
rect 194560 43404 244280 43432
rect 194560 43392 194566 43404
rect 244274 43392 244280 43404
rect 244332 43392 244338 43444
rect 245470 43392 245476 43444
rect 245528 43432 245534 43444
rect 302234 43432 302240 43444
rect 245528 43404 302240 43432
rect 245528 43392 245534 43404
rect 302234 43392 302240 43404
rect 302292 43392 302298 43444
rect 304902 43392 304908 43444
rect 304960 43432 304966 43444
rect 365714 43432 365720 43444
rect 304960 43404 365720 43432
rect 304960 43392 304966 43404
rect 365714 43392 365720 43404
rect 365772 43392 365778 43444
rect 415302 43392 415308 43444
rect 415360 43432 415366 43444
rect 487154 43432 487160 43444
rect 415360 43404 487160 43432
rect 415360 43392 415366 43404
rect 487154 43392 487160 43404
rect 487212 43392 487218 43444
rect 488350 43392 488356 43444
rect 488408 43432 488414 43444
rect 565814 43432 565820 43444
rect 488408 43404 565820 43432
rect 488408 43392 488414 43404
rect 565814 43392 565820 43404
rect 565872 43392 565878 43444
rect 122650 42100 122656 42152
rect 122708 42140 122714 42152
rect 166994 42140 167000 42152
rect 122708 42112 167000 42140
rect 122708 42100 122714 42112
rect 166994 42100 167000 42112
rect 167052 42100 167058 42152
rect 348970 42100 348976 42152
rect 349028 42140 349034 42152
rect 414014 42140 414020 42152
rect 349028 42112 414020 42140
rect 349028 42100 349034 42112
rect 414014 42100 414020 42112
rect 414072 42100 414078 42152
rect 165522 42032 165528 42084
rect 165580 42072 165586 42084
rect 213914 42072 213920 42084
rect 165580 42044 213920 42072
rect 165580 42032 165586 42044
rect 213914 42032 213920 42044
rect 213972 42032 213978 42084
rect 229002 42032 229008 42084
rect 229060 42072 229066 42084
rect 282914 42072 282920 42084
rect 229060 42044 282920 42072
rect 229060 42032 229066 42044
rect 282914 42032 282920 42044
rect 282972 42032 282978 42084
rect 295242 42032 295248 42084
rect 295300 42072 295306 42084
rect 356146 42072 356152 42084
rect 295300 42044 356152 42072
rect 295300 42032 295306 42044
rect 356146 42032 356152 42044
rect 356204 42032 356210 42084
rect 412542 42032 412548 42084
rect 412600 42072 412606 42084
rect 484394 42072 484400 42084
rect 412600 42044 484400 42072
rect 412600 42032 412606 42044
rect 484394 42032 484400 42044
rect 484452 42032 484458 42084
rect 493962 42032 493968 42084
rect 494020 42072 494026 42084
rect 572714 42072 572720 42084
rect 494020 42044 572720 42072
rect 494020 42032 494026 42044
rect 572714 42032 572720 42044
rect 572772 42032 572778 42084
rect 235721 41463 235779 41469
rect 235721 41429 235733 41463
rect 235767 41460 235779 41463
rect 235810 41460 235816 41472
rect 235767 41432 235816 41460
rect 235767 41429 235779 41432
rect 235721 41423 235779 41429
rect 235810 41420 235816 41432
rect 235868 41420 235874 41472
rect 504450 41352 504456 41404
rect 504508 41392 504514 41404
rect 580166 41392 580172 41404
rect 504508 41364 580172 41392
rect 504508 41352 504514 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 345658 40740 345664 40792
rect 345716 40780 345722 40792
rect 408586 40780 408592 40792
rect 345716 40752 408592 40780
rect 345716 40740 345722 40752
rect 408586 40740 408592 40752
rect 408644 40740 408650 40792
rect 119982 40672 119988 40724
rect 120040 40712 120046 40724
rect 164234 40712 164240 40724
rect 120040 40684 164240 40712
rect 120040 40672 120046 40684
rect 164234 40672 164240 40684
rect 164292 40672 164298 40724
rect 173710 40672 173716 40724
rect 173768 40712 173774 40724
rect 223574 40712 223580 40724
rect 173768 40684 223580 40712
rect 173768 40672 173774 40684
rect 223574 40672 223580 40684
rect 223632 40672 223638 40724
rect 230382 40672 230388 40724
rect 230440 40712 230446 40724
rect 284294 40712 284300 40724
rect 230440 40684 284300 40712
rect 230440 40672 230446 40684
rect 284294 40672 284300 40684
rect 284352 40672 284358 40724
rect 285582 40672 285588 40724
rect 285640 40712 285646 40724
rect 345014 40712 345020 40724
rect 285640 40684 345020 40712
rect 285640 40672 285646 40684
rect 345014 40672 345020 40684
rect 345072 40672 345078 40724
rect 408402 40672 408408 40724
rect 408460 40712 408466 40724
rect 478874 40712 478880 40724
rect 408460 40684 478880 40712
rect 408460 40672 408466 40684
rect 478874 40672 478880 40684
rect 478932 40672 478938 40724
rect 115842 39312 115848 39364
rect 115900 39352 115906 39364
rect 158714 39352 158720 39364
rect 115900 39324 158720 39352
rect 115900 39312 115906 39324
rect 158714 39312 158720 39324
rect 158772 39312 158778 39364
rect 162762 39312 162768 39364
rect 162820 39352 162826 39364
rect 209774 39352 209780 39364
rect 162820 39324 209780 39352
rect 162820 39312 162826 39324
rect 209774 39312 209780 39324
rect 209832 39312 209838 39364
rect 215202 39312 215208 39364
rect 215260 39352 215266 39364
rect 269114 39352 269120 39364
rect 215260 39324 269120 39352
rect 215260 39312 215266 39324
rect 269114 39312 269120 39324
rect 269172 39312 269178 39364
rect 291102 39312 291108 39364
rect 291160 39352 291166 39364
rect 350534 39352 350540 39364
rect 291160 39324 350540 39352
rect 291160 39312 291166 39324
rect 350534 39312 350540 39324
rect 350592 39312 350598 39364
rect 365622 39312 365628 39364
rect 365680 39352 365686 39364
rect 433426 39352 433432 39364
rect 365680 39324 433432 39352
rect 365680 39312 365686 39324
rect 433426 39312 433432 39324
rect 433484 39312 433490 39364
rect 438762 39312 438768 39364
rect 438820 39352 438826 39364
rect 511994 39352 512000 39364
rect 438820 39324 512000 39352
rect 438820 39312 438826 39324
rect 511994 39312 512000 39324
rect 512052 39312 512058 39364
rect 353294 38564 353300 38616
rect 353352 38604 353358 38616
rect 353386 38604 353392 38616
rect 353352 38576 353392 38604
rect 353352 38564 353358 38576
rect 353386 38564 353392 38576
rect 353444 38564 353450 38616
rect 378134 38604 378140 38616
rect 378095 38576 378140 38604
rect 378134 38564 378140 38576
rect 378192 38564 378198 38616
rect 495434 38604 495440 38616
rect 495395 38576 495440 38604
rect 495434 38564 495440 38576
rect 495492 38564 495498 38616
rect 108942 37884 108948 37936
rect 109000 37924 109006 37936
rect 151814 37924 151820 37936
rect 109000 37896 151820 37924
rect 109000 37884 109006 37896
rect 151814 37884 151820 37896
rect 151872 37884 151878 37936
rect 158622 37884 158628 37936
rect 158680 37924 158686 37936
rect 205634 37924 205640 37936
rect 158680 37896 205640 37924
rect 158680 37884 158686 37896
rect 205634 37884 205640 37896
rect 205692 37884 205698 37936
rect 206922 37884 206928 37936
rect 206980 37924 206986 37936
rect 259454 37924 259460 37936
rect 206980 37896 259460 37924
rect 206980 37884 206986 37896
rect 259454 37884 259460 37896
rect 259512 37884 259518 37936
rect 262122 37884 262128 37936
rect 262180 37924 262186 37936
rect 320174 37924 320180 37936
rect 262180 37896 320180 37924
rect 262180 37884 262186 37896
rect 320174 37884 320180 37896
rect 320232 37884 320238 37936
rect 331122 37884 331128 37936
rect 331180 37924 331186 37936
rect 394694 37924 394700 37936
rect 331180 37896 394700 37924
rect 331180 37884 331186 37896
rect 394694 37884 394700 37896
rect 394752 37884 394758 37936
rect 405642 37884 405648 37936
rect 405700 37924 405706 37936
rect 476114 37924 476120 37936
rect 405700 37896 476120 37924
rect 405700 37884 405706 37896
rect 476114 37884 476120 37896
rect 476172 37884 476178 37936
rect 477402 37884 477408 37936
rect 477460 37924 477466 37936
rect 554866 37924 554872 37936
rect 477460 37896 554872 37924
rect 477460 37884 477466 37896
rect 554866 37884 554872 37896
rect 554924 37884 554930 37936
rect 371234 37312 371240 37324
rect 371195 37284 371240 37312
rect 371234 37272 371240 37284
rect 371292 37272 371298 37324
rect 154482 36592 154488 36644
rect 154540 36632 154546 36644
rect 201494 36632 201500 36644
rect 154540 36604 201500 36632
rect 154540 36592 154546 36604
rect 201494 36592 201500 36604
rect 201552 36592 201558 36644
rect 106182 36524 106188 36576
rect 106240 36564 106246 36576
rect 149054 36564 149060 36576
rect 106240 36536 149060 36564
rect 106240 36524 106246 36536
rect 149054 36524 149060 36536
rect 149112 36524 149118 36576
rect 198642 36524 198648 36576
rect 198700 36564 198706 36576
rect 249794 36564 249800 36576
rect 198700 36536 249800 36564
rect 198700 36524 198706 36536
rect 249794 36524 249800 36536
rect 249852 36524 249858 36576
rect 251082 36524 251088 36576
rect 251140 36564 251146 36576
rect 307754 36564 307760 36576
rect 251140 36536 307760 36564
rect 251140 36524 251146 36536
rect 307754 36524 307760 36536
rect 307812 36524 307818 36576
rect 311802 36524 311808 36576
rect 311860 36564 311866 36576
rect 374086 36564 374092 36576
rect 311860 36536 374092 36564
rect 311860 36524 311866 36536
rect 374086 36524 374092 36536
rect 374144 36524 374150 36576
rect 401502 36524 401508 36576
rect 401560 36564 401566 36576
rect 471974 36564 471980 36576
rect 401560 36536 471980 36564
rect 401560 36524 401566 36536
rect 471974 36524 471980 36536
rect 472032 36524 472038 36576
rect 484302 36524 484308 36576
rect 484360 36564 484366 36576
rect 563146 36564 563152 36576
rect 484360 36536 563152 36564
rect 484360 36524 484366 36536
rect 563146 36524 563152 36536
rect 563204 36524 563210 36576
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 14458 35884 14464 35896
rect 3476 35856 14464 35884
rect 3476 35844 3482 35856
rect 14458 35844 14464 35856
rect 14516 35844 14522 35896
rect 410886 35884 410892 35896
rect 410847 35856 410892 35884
rect 410886 35844 410892 35856
rect 410944 35844 410950 35896
rect 102042 35164 102048 35216
rect 102100 35204 102106 35216
rect 144914 35204 144920 35216
rect 102100 35176 144920 35204
rect 102100 35164 102106 35176
rect 144914 35164 144920 35176
rect 144972 35164 144978 35216
rect 151722 35164 151728 35216
rect 151780 35204 151786 35216
rect 198734 35204 198740 35216
rect 151780 35176 198740 35204
rect 151780 35164 151786 35176
rect 198734 35164 198740 35176
rect 198792 35164 198798 35216
rect 199930 35164 199936 35216
rect 199988 35204 199994 35216
rect 252646 35204 252652 35216
rect 199988 35176 252652 35204
rect 199988 35164 199994 35176
rect 252646 35164 252652 35176
rect 252704 35164 252710 35216
rect 259362 35164 259368 35216
rect 259420 35204 259426 35216
rect 316034 35204 316040 35216
rect 259420 35176 316040 35204
rect 259420 35164 259426 35176
rect 316034 35164 316040 35176
rect 316092 35164 316098 35216
rect 321462 35164 321468 35216
rect 321520 35204 321526 35216
rect 383654 35204 383660 35216
rect 321520 35176 383660 35204
rect 321520 35164 321526 35176
rect 383654 35164 383660 35176
rect 383712 35164 383718 35216
rect 398742 35164 398748 35216
rect 398800 35204 398806 35216
rect 467926 35204 467932 35216
rect 398800 35176 467932 35204
rect 398800 35164 398806 35176
rect 467926 35164 467932 35176
rect 467984 35164 467990 35216
rect 481542 35164 481548 35216
rect 481600 35204 481606 35216
rect 558914 35204 558920 35216
rect 481600 35176 558920 35204
rect 481600 35164 481606 35176
rect 558914 35164 558920 35176
rect 558972 35164 558978 35216
rect 144822 33804 144828 33856
rect 144880 33844 144886 33856
rect 191834 33844 191840 33856
rect 144880 33816 191840 33844
rect 144880 33804 144886 33816
rect 191834 33804 191840 33816
rect 191892 33804 191898 33856
rect 99282 33736 99288 33788
rect 99340 33776 99346 33788
rect 140774 33776 140780 33788
rect 99340 33748 140780 33776
rect 99340 33736 99346 33748
rect 140774 33736 140780 33748
rect 140832 33736 140838 33788
rect 190362 33736 190368 33788
rect 190420 33776 190426 33788
rect 241514 33776 241520 33788
rect 190420 33748 241520 33776
rect 190420 33736 190426 33748
rect 241514 33736 241520 33748
rect 241572 33736 241578 33788
rect 277302 33736 277308 33788
rect 277360 33776 277366 33788
rect 336734 33776 336740 33788
rect 277360 33748 336740 33776
rect 277360 33736 277366 33748
rect 336734 33736 336740 33748
rect 336792 33736 336798 33788
rect 337378 33736 337384 33788
rect 337436 33776 337442 33788
rect 389174 33776 389180 33788
rect 337436 33748 389180 33776
rect 337436 33736 337442 33748
rect 389174 33736 389180 33748
rect 389232 33736 389238 33788
rect 395982 33736 395988 33788
rect 396040 33776 396046 33788
rect 465074 33776 465080 33788
rect 396040 33748 465080 33776
rect 396040 33736 396046 33748
rect 465074 33736 465080 33748
rect 465132 33736 465138 33788
rect 474642 33736 474648 33788
rect 474700 33776 474706 33788
rect 552014 33776 552020 33788
rect 474700 33748 552020 33776
rect 474700 33736 474706 33748
rect 552014 33736 552020 33748
rect 552072 33736 552078 33788
rect 142062 32444 142068 32496
rect 142120 32484 142126 32496
rect 187694 32484 187700 32496
rect 142120 32456 187700 32484
rect 142120 32444 142126 32456
rect 187694 32444 187700 32456
rect 187752 32444 187758 32496
rect 249702 32444 249708 32496
rect 249760 32484 249766 32496
rect 304994 32484 305000 32496
rect 249760 32456 305000 32484
rect 249760 32444 249766 32456
rect 304994 32444 305000 32456
rect 305052 32444 305058 32496
rect 96430 32376 96436 32428
rect 96488 32416 96494 32428
rect 138014 32416 138020 32428
rect 96488 32388 138020 32416
rect 96488 32376 96494 32388
rect 138014 32376 138020 32388
rect 138072 32376 138078 32428
rect 187602 32376 187608 32428
rect 187660 32416 187666 32428
rect 237374 32416 237380 32428
rect 187660 32388 237380 32416
rect 187660 32376 187666 32388
rect 237374 32376 237380 32388
rect 237432 32376 237438 32428
rect 302142 32376 302148 32428
rect 302200 32416 302206 32428
rect 362954 32416 362960 32428
rect 302200 32388 362960 32416
rect 302200 32376 302206 32388
rect 362954 32376 362960 32388
rect 363012 32376 363018 32428
rect 391842 32376 391848 32428
rect 391900 32416 391906 32428
rect 460934 32416 460940 32428
rect 391900 32388 460940 32416
rect 391900 32376 391906 32388
rect 460934 32376 460940 32388
rect 460992 32376 460998 32428
rect 471790 32376 471796 32428
rect 471848 32416 471854 32428
rect 547874 32416 547880 32428
rect 471848 32388 547880 32416
rect 471848 32376 471854 32388
rect 547874 32376 547880 32388
rect 547932 32376 547938 32428
rect 137922 31016 137928 31068
rect 137980 31056 137986 31068
rect 183554 31056 183560 31068
rect 137980 31028 183560 31056
rect 137980 31016 137986 31028
rect 183554 31016 183560 31028
rect 183612 31016 183618 31068
rect 185578 31016 185584 31068
rect 185636 31056 185642 31068
rect 234614 31056 234620 31068
rect 185636 31028 234620 31056
rect 185636 31016 185642 31028
rect 234614 31016 234620 31028
rect 234672 31016 234678 31068
rect 240042 31016 240048 31068
rect 240100 31056 240106 31068
rect 295334 31056 295340 31068
rect 240100 31028 295340 31056
rect 240100 31016 240106 31028
rect 295334 31016 295340 31028
rect 295392 31016 295398 31068
rect 313182 31016 313188 31068
rect 313240 31056 313246 31068
rect 375374 31056 375380 31068
rect 313240 31028 375380 31056
rect 313240 31016 313246 31028
rect 375374 31016 375380 31028
rect 375432 31016 375438 31068
rect 389082 31016 389088 31068
rect 389140 31056 389146 31068
rect 458174 31056 458180 31068
rect 389140 31028 458180 31056
rect 389140 31016 389146 31028
rect 458174 31016 458180 31028
rect 458232 31016 458238 31068
rect 464982 31016 464988 31068
rect 465040 31056 465046 31068
rect 540974 31056 540980 31068
rect 465040 31028 540980 31056
rect 465040 31016 465046 31028
rect 540974 31016 540980 31028
rect 541032 31016 541038 31068
rect 504358 30268 504364 30320
rect 504416 30308 504422 30320
rect 580166 30308 580172 30320
rect 504416 30280 580172 30308
rect 504416 30268 504422 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 135162 29656 135168 29708
rect 135220 29696 135226 29708
rect 180794 29696 180800 29708
rect 135220 29668 180800 29696
rect 135220 29656 135226 29668
rect 180794 29656 180800 29668
rect 180852 29656 180858 29708
rect 92290 29588 92296 29640
rect 92348 29628 92354 29640
rect 133874 29628 133880 29640
rect 92348 29600 133880 29628
rect 92348 29588 92354 29600
rect 133874 29588 133880 29600
rect 133932 29588 133938 29640
rect 180702 29588 180708 29640
rect 180760 29628 180766 29640
rect 230474 29628 230480 29640
rect 180760 29600 230480 29628
rect 180760 29588 180766 29600
rect 230474 29588 230480 29600
rect 230532 29588 230538 29640
rect 235721 29631 235779 29637
rect 235721 29597 235733 29631
rect 235767 29628 235779 29631
rect 291194 29628 291200 29640
rect 235767 29600 291200 29628
rect 235767 29597 235779 29600
rect 235721 29591 235779 29597
rect 291194 29588 291200 29600
rect 291252 29588 291258 29640
rect 310422 29588 310428 29640
rect 310480 29628 310486 29640
rect 372614 29628 372620 29640
rect 310480 29600 372620 29628
rect 310480 29588 310486 29600
rect 372614 29588 372620 29600
rect 372672 29588 372678 29640
rect 380158 29588 380164 29640
rect 380216 29628 380222 29640
rect 447134 29628 447140 29640
rect 380216 29600 447140 29628
rect 380216 29588 380222 29600
rect 447134 29588 447140 29600
rect 447192 29588 447198 29640
rect 378134 29084 378140 29096
rect 378095 29056 378140 29084
rect 378134 29044 378140 29056
rect 378192 29044 378198 29096
rect 495434 29016 495440 29028
rect 495395 28988 495440 29016
rect 495434 28976 495440 28988
rect 495492 28976 495498 29028
rect 378134 28908 378140 28960
rect 378192 28948 378198 28960
rect 378226 28948 378232 28960
rect 378192 28920 378232 28948
rect 378192 28908 378198 28920
rect 378226 28908 378232 28920
rect 378284 28908 378290 28960
rect 89622 28228 89628 28280
rect 89680 28268 89686 28280
rect 131114 28268 131120 28280
rect 89680 28240 131120 28268
rect 89680 28228 89686 28240
rect 131114 28228 131120 28240
rect 131172 28228 131178 28280
rect 132402 28228 132408 28280
rect 132460 28268 132466 28280
rect 176654 28268 176660 28280
rect 132460 28240 176660 28268
rect 132460 28228 132466 28240
rect 176654 28228 176660 28240
rect 176712 28228 176718 28280
rect 177942 28228 177948 28280
rect 178000 28268 178006 28280
rect 227806 28268 227812 28280
rect 178000 28240 227812 28268
rect 178000 28228 178006 28240
rect 227806 28228 227812 28240
rect 227864 28228 227870 28280
rect 233142 28228 233148 28280
rect 233200 28268 233206 28280
rect 287146 28268 287152 28280
rect 233200 28240 287152 28268
rect 233200 28228 233206 28240
rect 287146 28228 287152 28240
rect 287204 28228 287210 28280
rect 288342 28228 288348 28280
rect 288400 28268 288406 28280
rect 347774 28268 347780 28280
rect 288400 28240 347780 28268
rect 288400 28228 288406 28240
rect 347774 28228 347780 28240
rect 347832 28228 347838 28280
rect 375282 28228 375288 28280
rect 375340 28268 375346 28280
rect 443086 28268 443092 28280
rect 375340 28240 443092 28268
rect 375340 28228 375346 28240
rect 443086 28228 443092 28240
rect 443144 28228 443150 28280
rect 448422 28228 448428 28280
rect 448480 28268 448486 28280
rect 523034 28268 523040 28280
rect 448480 28240 523040 28268
rect 448480 28228 448486 28240
rect 523034 28228 523040 28240
rect 523092 28228 523098 28280
rect 353294 27548 353300 27600
rect 353352 27588 353358 27600
rect 353846 27588 353852 27600
rect 353352 27560 353852 27588
rect 353352 27548 353358 27560
rect 353846 27548 353852 27560
rect 353904 27548 353910 27600
rect 371234 27588 371240 27600
rect 371195 27560 371240 27588
rect 371234 27548 371240 27560
rect 371292 27548 371298 27600
rect 128262 26936 128268 26988
rect 128320 26976 128326 26988
rect 173894 26976 173900 26988
rect 128320 26948 173900 26976
rect 128320 26936 128326 26948
rect 173894 26936 173900 26948
rect 173952 26936 173958 26988
rect 171042 26868 171048 26920
rect 171100 26908 171106 26920
rect 219434 26908 219440 26920
rect 171100 26880 219440 26908
rect 171100 26868 171106 26880
rect 219434 26868 219440 26880
rect 219492 26868 219498 26920
rect 223482 26868 223488 26920
rect 223540 26908 223546 26920
rect 277394 26908 277400 26920
rect 223540 26880 277400 26908
rect 223540 26868 223546 26880
rect 277394 26868 277400 26880
rect 277452 26868 277458 26920
rect 278682 26868 278688 26920
rect 278740 26908 278746 26920
rect 338114 26908 338120 26920
rect 278740 26880 338120 26908
rect 278740 26868 278746 26880
rect 338114 26868 338120 26880
rect 338172 26868 338178 26920
rect 372522 26868 372528 26920
rect 372580 26908 372586 26920
rect 440234 26908 440240 26920
rect 372580 26880 440240 26908
rect 372580 26868 372586 26880
rect 440234 26868 440240 26880
rect 440292 26868 440298 26920
rect 445662 26868 445668 26920
rect 445720 26908 445726 26920
rect 520366 26908 520372 26920
rect 445720 26880 520372 26908
rect 445720 26868 445726 26880
rect 520366 26868 520372 26880
rect 520424 26868 520430 26920
rect 410889 26299 410947 26305
rect 410889 26265 410901 26299
rect 410935 26296 410947 26299
rect 410978 26296 410984 26308
rect 410935 26268 410984 26296
rect 410935 26265 410947 26268
rect 410889 26259 410947 26265
rect 410978 26256 410984 26268
rect 411036 26256 411042 26308
rect 125502 25576 125508 25628
rect 125560 25616 125566 25628
rect 169754 25616 169760 25628
rect 125560 25588 169760 25616
rect 125560 25576 125566 25588
rect 169754 25576 169760 25588
rect 169812 25576 169818 25628
rect 216582 25576 216588 25628
rect 216640 25616 216646 25628
rect 270586 25616 270592 25628
rect 216640 25588 270592 25616
rect 216640 25576 216646 25588
rect 270586 25576 270592 25588
rect 270644 25576 270650 25628
rect 168282 25508 168288 25560
rect 168340 25548 168346 25560
rect 216674 25548 216680 25560
rect 168340 25520 216680 25548
rect 168340 25508 168346 25520
rect 216674 25508 216680 25520
rect 216732 25508 216738 25560
rect 266170 25508 266176 25560
rect 266228 25548 266234 25560
rect 322934 25548 322940 25560
rect 266228 25520 322940 25548
rect 266228 25508 266234 25520
rect 322934 25508 322940 25520
rect 322992 25508 322998 25560
rect 362862 25508 362868 25560
rect 362920 25548 362926 25560
rect 429194 25548 429200 25560
rect 362920 25520 429200 25548
rect 362920 25508 362926 25520
rect 429194 25508 429200 25520
rect 429252 25508 429258 25560
rect 482830 25508 482836 25560
rect 482888 25548 482894 25560
rect 561674 25548 561680 25560
rect 482888 25520 561680 25548
rect 482888 25508 482894 25520
rect 561674 25508 561680 25520
rect 561732 25508 561738 25560
rect 202782 24148 202788 24200
rect 202840 24188 202846 24200
rect 253934 24188 253940 24200
rect 202840 24160 253940 24188
rect 202840 24148 202846 24160
rect 253934 24148 253940 24160
rect 253992 24148 253998 24200
rect 122742 24080 122748 24132
rect 122800 24120 122806 24132
rect 167086 24120 167092 24132
rect 122800 24092 167092 24120
rect 122800 24080 122806 24092
rect 167086 24080 167092 24092
rect 167144 24080 167150 24132
rect 252462 24080 252468 24132
rect 252520 24120 252526 24132
rect 309134 24120 309140 24132
rect 252520 24092 309140 24120
rect 252520 24080 252526 24092
rect 309134 24080 309140 24092
rect 309192 24080 309198 24132
rect 349062 24080 349068 24132
rect 349120 24120 349126 24132
rect 415394 24120 415400 24132
rect 349120 24092 415400 24120
rect 349120 24080 349126 24092
rect 415394 24080 415400 24092
rect 415452 24080 415458 24132
rect 470502 24080 470508 24132
rect 470560 24120 470566 24132
rect 546586 24120 546592 24132
rect 470560 24092 546592 24120
rect 470560 24080 470566 24092
rect 546586 24080 546592 24092
rect 546644 24080 546650 24132
rect 161382 22788 161388 22840
rect 161440 22828 161446 22840
rect 209866 22828 209872 22840
rect 161440 22800 209872 22828
rect 161440 22788 161446 22800
rect 209866 22788 209872 22800
rect 209924 22788 209930 22840
rect 118602 22720 118608 22772
rect 118660 22760 118666 22772
rect 162854 22760 162860 22772
rect 118660 22732 162860 22760
rect 118660 22720 118666 22732
rect 162854 22720 162860 22732
rect 162912 22720 162918 22772
rect 204162 22720 204168 22772
rect 204220 22760 204226 22772
rect 255314 22760 255320 22772
rect 204220 22732 255320 22760
rect 204220 22720 204226 22732
rect 255314 22720 255320 22732
rect 255372 22720 255378 22772
rect 256602 22720 256608 22772
rect 256660 22760 256666 22772
rect 313366 22760 313372 22772
rect 256660 22732 313372 22760
rect 256660 22720 256666 22732
rect 313366 22720 313372 22732
rect 313424 22720 313430 22772
rect 333882 22720 333888 22772
rect 333940 22760 333946 22772
rect 397546 22760 397552 22772
rect 333940 22732 397552 22760
rect 333940 22720 333946 22732
rect 397546 22720 397552 22732
rect 397604 22720 397610 22772
rect 453942 22720 453948 22772
rect 454000 22760 454006 22772
rect 528646 22760 528652 22772
rect 454000 22732 528652 22760
rect 454000 22720 454006 22732
rect 528646 22720 528652 22732
rect 528704 22720 528710 22772
rect 410889 22151 410947 22157
rect 410889 22117 410901 22151
rect 410935 22148 410947 22151
rect 410978 22148 410984 22160
rect 410935 22120 410984 22148
rect 410935 22117 410947 22120
rect 410889 22111 410947 22117
rect 410978 22108 410984 22120
rect 411036 22108 411042 22160
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 79410 22080 79416 22092
rect 3200 22052 79416 22080
rect 3200 22040 3206 22052
rect 79410 22040 79416 22052
rect 79468 22040 79474 22092
rect 226242 21428 226248 21480
rect 226300 21468 226306 21480
rect 278866 21468 278872 21480
rect 226300 21440 278872 21468
rect 226300 21428 226306 21440
rect 278866 21428 278872 21440
rect 278924 21428 278930 21480
rect 322842 21428 322848 21480
rect 322900 21468 322906 21480
rect 386414 21468 386420 21480
rect 322900 21440 386420 21468
rect 322900 21428 322906 21440
rect 386414 21428 386420 21440
rect 386472 21428 386478 21480
rect 114462 21360 114468 21412
rect 114520 21400 114526 21412
rect 158806 21400 158812 21412
rect 114520 21372 158812 21400
rect 114520 21360 114526 21372
rect 158806 21360 158812 21372
rect 158864 21360 158870 21412
rect 166902 21360 166908 21412
rect 166960 21400 166966 21412
rect 215294 21400 215300 21412
rect 166960 21372 215300 21400
rect 166960 21360 166966 21372
rect 215294 21360 215300 21372
rect 215352 21360 215358 21412
rect 266262 21360 266268 21412
rect 266320 21400 266326 21412
rect 324314 21400 324320 21412
rect 266320 21372 324320 21400
rect 266320 21360 266326 21372
rect 324314 21360 324320 21372
rect 324372 21360 324378 21412
rect 384850 21360 384856 21412
rect 384908 21400 384914 21412
rect 454034 21400 454040 21412
rect 384908 21372 454040 21400
rect 384908 21360 384914 21372
rect 454034 21360 454040 21372
rect 454092 21360 454098 21412
rect 467742 21360 467748 21412
rect 467800 21400 467806 21412
rect 543734 21400 543740 21412
rect 467800 21372 543740 21400
rect 467800 21360 467806 21372
rect 543734 21360 543740 21372
rect 543792 21360 543798 21412
rect 111702 19932 111708 19984
rect 111760 19972 111766 19984
rect 154574 19972 154580 19984
rect 111760 19944 154580 19972
rect 111760 19932 111766 19944
rect 154574 19932 154580 19944
rect 154632 19932 154638 19984
rect 157242 19932 157248 19984
rect 157300 19972 157306 19984
rect 204254 19972 204260 19984
rect 157300 19944 204260 19972
rect 157300 19932 157306 19944
rect 204254 19932 204260 19944
rect 204312 19932 204318 19984
rect 205542 19932 205548 19984
rect 205600 19972 205606 19984
rect 258074 19972 258080 19984
rect 205600 19944 258080 19972
rect 205600 19932 205606 19944
rect 258074 19932 258080 19944
rect 258132 19932 258138 19984
rect 293862 19932 293868 19984
rect 293920 19972 293926 19984
rect 354674 19972 354680 19984
rect 293920 19944 354680 19972
rect 293920 19932 293926 19944
rect 354674 19932 354680 19944
rect 354732 19932 354738 19984
rect 355962 19932 355968 19984
rect 356020 19972 356026 19984
rect 422294 19972 422300 19984
rect 356020 19944 422300 19972
rect 356020 19932 356026 19944
rect 422294 19932 422300 19944
rect 422352 19932 422358 19984
rect 463602 19932 463608 19984
rect 463660 19972 463666 19984
rect 539594 19972 539600 19984
rect 463660 19944 539600 19972
rect 463660 19932 463666 19944
rect 539594 19932 539600 19944
rect 539652 19932 539658 19984
rect 369854 19292 369860 19304
rect 369815 19264 369860 19292
rect 369854 19252 369860 19264
rect 369912 19252 369918 19304
rect 378134 19292 378140 19304
rect 378095 19264 378140 19292
rect 378134 19252 378140 19264
rect 378192 19252 378198 19304
rect 389174 19252 389180 19304
rect 389232 19292 389238 19304
rect 389358 19292 389364 19304
rect 389232 19264 389364 19292
rect 389232 19252 389238 19264
rect 389358 19252 389364 19264
rect 389416 19252 389422 19304
rect 397454 19292 397460 19304
rect 397415 19264 397460 19292
rect 397454 19252 397460 19264
rect 397512 19252 397518 19304
rect 408586 19252 408592 19304
rect 408644 19292 408650 19304
rect 409690 19292 409696 19304
rect 408644 19264 409696 19292
rect 408644 19252 408650 19264
rect 409690 19252 409696 19264
rect 409748 19252 409754 19304
rect 414014 19252 414020 19304
rect 414072 19292 414078 19304
rect 414474 19292 414480 19304
rect 414072 19264 414480 19292
rect 414072 19252 414078 19264
rect 414474 19252 414480 19264
rect 414532 19252 414538 19304
rect 415394 19252 415400 19304
rect 415452 19292 415458 19304
rect 415452 19264 415497 19292
rect 415452 19252 415458 19264
rect 495434 19252 495440 19304
rect 495492 19292 495498 19304
rect 495618 19292 495624 19304
rect 495492 19264 495624 19292
rect 495492 19252 495498 19264
rect 495618 19252 495624 19264
rect 495676 19252 495682 19304
rect 561674 19292 561680 19304
rect 561635 19264 561680 19292
rect 561674 19252 561680 19264
rect 561732 19252 561738 19304
rect 113818 18572 113824 18624
rect 113876 18612 113882 18624
rect 150526 18612 150532 18624
rect 113876 18584 150532 18612
rect 113876 18572 113882 18584
rect 150526 18572 150532 18584
rect 150584 18572 150590 18624
rect 153838 18572 153844 18624
rect 153896 18612 153902 18624
rect 201586 18612 201592 18624
rect 153896 18584 201592 18612
rect 153896 18572 153902 18584
rect 201586 18572 201592 18584
rect 201644 18572 201650 18624
rect 222102 18572 222108 18624
rect 222160 18612 222166 18624
rect 276014 18612 276020 18624
rect 222160 18584 276020 18612
rect 222160 18572 222166 18584
rect 276014 18572 276020 18584
rect 276072 18572 276078 18624
rect 284202 18572 284208 18624
rect 284260 18612 284266 18624
rect 343634 18612 343640 18624
rect 284260 18584 343640 18612
rect 284260 18572 284266 18584
rect 343634 18572 343640 18584
rect 343692 18572 343698 18624
rect 346302 18572 346308 18624
rect 346360 18612 346366 18624
rect 346360 18584 407804 18612
rect 346360 18572 346366 18584
rect 407776 18544 407804 18584
rect 411898 18572 411904 18624
rect 411956 18612 411962 18624
rect 455414 18612 455420 18624
rect 411956 18584 455420 18612
rect 411956 18572 411962 18584
rect 455414 18572 455420 18584
rect 455472 18572 455478 18624
rect 456702 18572 456708 18624
rect 456760 18612 456766 18624
rect 532694 18612 532700 18624
rect 456760 18584 532700 18612
rect 456760 18572 456766 18584
rect 532694 18572 532700 18584
rect 532752 18572 532758 18624
rect 412082 18544 412088 18556
rect 407776 18516 412088 18544
rect 412082 18504 412088 18516
rect 412140 18504 412146 18556
rect 371234 18000 371240 18012
rect 371195 17972 371240 18000
rect 371234 17960 371240 17972
rect 371292 17960 371298 18012
rect 571978 17892 571984 17944
rect 572036 17932 572042 17944
rect 579798 17932 579804 17944
rect 572036 17904 579804 17932
rect 572036 17892 572042 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 281442 17280 281448 17332
rect 281500 17320 281506 17332
rect 339586 17320 339592 17332
rect 281500 17292 339592 17320
rect 281500 17280 281506 17292
rect 339586 17280 339592 17292
rect 339644 17280 339650 17332
rect 104802 17212 104808 17264
rect 104860 17252 104866 17264
rect 147674 17252 147680 17264
rect 104860 17224 147680 17252
rect 104860 17212 104866 17224
rect 147674 17212 147680 17224
rect 147732 17212 147738 17264
rect 150342 17212 150348 17264
rect 150400 17252 150406 17264
rect 197354 17252 197360 17264
rect 150400 17224 197360 17252
rect 150400 17212 150406 17224
rect 197354 17212 197360 17224
rect 197412 17212 197418 17264
rect 209682 17212 209688 17264
rect 209740 17252 209746 17264
rect 262306 17252 262312 17264
rect 209740 17224 262312 17252
rect 209740 17212 209746 17224
rect 262306 17212 262312 17224
rect 262364 17212 262370 17264
rect 339402 17212 339408 17264
rect 339460 17252 339466 17264
rect 404354 17252 404360 17264
rect 339460 17224 404360 17252
rect 339460 17212 339466 17224
rect 404354 17212 404360 17224
rect 404412 17212 404418 17264
rect 451182 17212 451188 17264
rect 451240 17252 451246 17264
rect 525794 17252 525800 17264
rect 451240 17224 525800 17252
rect 451240 17212 451246 17224
rect 525794 17212 525800 17224
rect 525852 17212 525858 17264
rect 102778 15852 102784 15904
rect 102836 15892 102842 15904
rect 143534 15892 143540 15904
rect 102836 15864 143540 15892
rect 102836 15852 102842 15864
rect 143534 15852 143540 15864
rect 143592 15852 143598 15904
rect 147582 15852 147588 15904
rect 147640 15892 147646 15904
rect 193306 15892 193312 15904
rect 147640 15864 193312 15892
rect 147640 15852 147646 15864
rect 193306 15852 193312 15864
rect 193364 15852 193370 15904
rect 195882 15852 195888 15904
rect 195940 15892 195946 15904
rect 247034 15892 247040 15904
rect 195940 15864 247040 15892
rect 195940 15852 195946 15864
rect 247034 15852 247040 15864
rect 247092 15852 247098 15904
rect 267642 15852 267648 15904
rect 267700 15892 267706 15904
rect 325694 15892 325700 15904
rect 267700 15864 325700 15892
rect 267700 15852 267706 15864
rect 325694 15852 325700 15864
rect 325752 15852 325758 15904
rect 326982 15852 326988 15904
rect 327040 15892 327046 15904
rect 390646 15892 390652 15904
rect 327040 15864 390652 15892
rect 327040 15852 327046 15864
rect 390646 15852 390652 15864
rect 390704 15852 390710 15904
rect 437382 15852 437388 15904
rect 437440 15892 437446 15904
rect 512086 15892 512092 15904
rect 437440 15864 512092 15892
rect 437440 15852 437446 15864
rect 512086 15852 512092 15864
rect 512144 15852 512150 15904
rect 320082 14492 320088 14544
rect 320140 14532 320146 14544
rect 382366 14532 382372 14544
rect 320140 14504 382372 14532
rect 320140 14492 320146 14504
rect 382366 14492 382372 14504
rect 382424 14492 382430 14544
rect 97902 14424 97908 14476
rect 97960 14464 97966 14476
rect 140866 14464 140872 14476
rect 97960 14436 140872 14464
rect 97960 14424 97966 14436
rect 140866 14424 140872 14436
rect 140924 14424 140930 14476
rect 143442 14424 143448 14476
rect 143500 14464 143506 14476
rect 190454 14464 190460 14476
rect 143500 14436 190460 14464
rect 143500 14424 143506 14436
rect 190454 14424 190460 14436
rect 190512 14424 190518 14476
rect 193122 14424 193128 14476
rect 193180 14464 193186 14476
rect 244366 14464 244372 14476
rect 193180 14436 244372 14464
rect 193180 14424 193186 14436
rect 244366 14424 244372 14436
rect 244424 14424 244430 14476
rect 257982 14424 257988 14476
rect 258040 14464 258046 14476
rect 314654 14464 314660 14476
rect 258040 14436 314660 14464
rect 258040 14424 258046 14436
rect 314654 14424 314660 14436
rect 314712 14424 314718 14476
rect 382182 14424 382188 14476
rect 382240 14464 382246 14476
rect 451366 14464 451372 14476
rect 382240 14436 451372 14464
rect 382240 14424 382246 14436
rect 451366 14424 451372 14436
rect 451424 14424 451430 14476
rect 460842 14424 460848 14476
rect 460900 14464 460906 14476
rect 536926 14464 536932 14476
rect 460900 14436 536932 14464
rect 460900 14424 460906 14436
rect 536926 14424 536932 14436
rect 536984 14424 536990 14476
rect 97258 13064 97264 13116
rect 97316 13104 97322 13116
rect 126974 13104 126980 13116
rect 97316 13076 126980 13104
rect 97316 13064 97322 13076
rect 126974 13064 126980 13076
rect 127032 13064 127038 13116
rect 140682 13064 140688 13116
rect 140740 13104 140746 13116
rect 186314 13104 186320 13116
rect 140740 13076 186320 13104
rect 140740 13064 140746 13076
rect 186314 13064 186320 13076
rect 186372 13064 186378 13116
rect 189718 13064 189724 13116
rect 189776 13104 189782 13116
rect 240134 13104 240140 13116
rect 189776 13076 240140 13104
rect 189776 13064 189782 13076
rect 240134 13064 240140 13076
rect 240192 13064 240198 13116
rect 255222 13064 255228 13116
rect 255280 13104 255286 13116
rect 311894 13104 311900 13116
rect 255280 13076 311900 13104
rect 255280 13064 255286 13076
rect 311894 13064 311900 13076
rect 311952 13064 311958 13116
rect 317322 13064 317328 13116
rect 317380 13104 317386 13116
rect 379514 13104 379520 13116
rect 317380 13076 379520 13104
rect 317380 13064 317386 13076
rect 379514 13064 379520 13076
rect 379572 13064 379578 13116
rect 434622 13064 434628 13116
rect 434680 13104 434686 13116
rect 507854 13104 507860 13116
rect 434680 13076 507860 13104
rect 434680 13064 434686 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 354674 12452 354680 12504
rect 354732 12452 354738 12504
rect 371234 12452 371240 12504
rect 371292 12452 371298 12504
rect 372614 12452 372620 12504
rect 372672 12452 372678 12504
rect 394694 12452 394700 12504
rect 394752 12452 394758 12504
rect 350534 12384 350540 12436
rect 350592 12424 350598 12436
rect 351362 12424 351368 12436
rect 350592 12396 351368 12424
rect 350592 12384 350598 12396
rect 351362 12384 351368 12396
rect 351420 12384 351426 12436
rect 351914 12384 351920 12436
rect 351972 12424 351978 12436
rect 352558 12424 352564 12436
rect 351972 12396 352564 12424
rect 351972 12384 351978 12396
rect 352558 12384 352564 12396
rect 352616 12384 352622 12436
rect 354692 12356 354720 12452
rect 358814 12384 358820 12436
rect 358872 12424 358878 12436
rect 359734 12424 359740 12436
rect 358872 12396 359740 12424
rect 358872 12384 358878 12396
rect 359734 12384 359740 12396
rect 359792 12384 359798 12436
rect 354950 12356 354956 12368
rect 354692 12328 354956 12356
rect 354950 12316 354956 12328
rect 355008 12316 355014 12368
rect 371252 12356 371280 12452
rect 371602 12356 371608 12368
rect 371252 12328 371608 12356
rect 371602 12316 371608 12328
rect 371660 12316 371666 12368
rect 372632 12356 372660 12452
rect 375374 12384 375380 12436
rect 375432 12424 375438 12436
rect 376386 12424 376392 12436
rect 375432 12396 376392 12424
rect 375432 12384 375438 12396
rect 376386 12384 376392 12396
rect 376444 12384 376450 12436
rect 376754 12384 376760 12436
rect 376812 12424 376818 12436
rect 377582 12424 377588 12436
rect 376812 12396 377588 12424
rect 376812 12384 376818 12396
rect 377582 12384 377588 12396
rect 377640 12384 377646 12436
rect 391934 12384 391940 12436
rect 391992 12424 391998 12436
rect 393038 12424 393044 12436
rect 391992 12396 393044 12424
rect 391992 12384 391998 12396
rect 393038 12384 393044 12396
rect 393096 12384 393102 12436
rect 393406 12384 393412 12436
rect 393464 12424 393470 12436
rect 394234 12424 394240 12436
rect 393464 12396 394240 12424
rect 393464 12384 393470 12396
rect 394234 12384 394240 12396
rect 394292 12384 394298 12436
rect 372798 12356 372804 12368
rect 372632 12328 372804 12356
rect 372798 12316 372804 12328
rect 372856 12316 372862 12368
rect 394712 12356 394740 12452
rect 396074 12384 396080 12436
rect 396132 12424 396138 12436
rect 396626 12424 396632 12436
rect 396132 12396 396632 12424
rect 396132 12384 396138 12396
rect 396626 12384 396632 12396
rect 396684 12384 396690 12436
rect 412634 12384 412640 12436
rect 412692 12424 412698 12436
rect 413278 12424 413284 12436
rect 412692 12396 413284 12424
rect 412692 12384 412698 12396
rect 413278 12384 413284 12396
rect 413336 12384 413342 12436
rect 554866 12384 554872 12436
rect 554924 12424 554930 12436
rect 555970 12424 555976 12436
rect 554924 12396 555976 12424
rect 554924 12384 554930 12396
rect 555970 12384 555976 12396
rect 556028 12384 556034 12436
rect 557534 12384 557540 12436
rect 557592 12424 557598 12436
rect 558362 12424 558368 12436
rect 557592 12396 558368 12424
rect 557592 12384 557598 12396
rect 558362 12384 558368 12396
rect 558420 12384 558426 12436
rect 558914 12384 558920 12436
rect 558972 12424 558978 12436
rect 559558 12424 559564 12436
rect 558972 12396 559564 12424
rect 558972 12384 558978 12396
rect 559558 12384 559564 12396
rect 559616 12384 559622 12436
rect 395430 12356 395436 12368
rect 394712 12328 395436 12356
rect 395430 12316 395436 12328
rect 395488 12316 395494 12368
rect 427722 11772 427728 11824
rect 427780 11812 427786 11824
rect 501230 11812 501236 11824
rect 427780 11784 501236 11812
rect 427780 11772 427786 11784
rect 501230 11772 501236 11784
rect 501288 11772 501294 11824
rect 92382 11704 92388 11756
rect 92440 11744 92446 11756
rect 132586 11744 132592 11756
rect 92440 11716 132592 11744
rect 92440 11704 92446 11716
rect 132586 11704 132592 11716
rect 132644 11704 132650 11756
rect 133782 11704 133788 11756
rect 133840 11744 133846 11756
rect 179414 11744 179420 11756
rect 133840 11716 179420 11744
rect 133840 11704 133846 11716
rect 179414 11704 179420 11716
rect 179472 11704 179478 11756
rect 183462 11704 183468 11756
rect 183520 11744 183526 11756
rect 233234 11744 233240 11756
rect 183520 11716 233240 11744
rect 183520 11704 183526 11716
rect 233234 11704 233240 11716
rect 233292 11704 233298 11756
rect 241422 11704 241428 11756
rect 241480 11744 241486 11756
rect 296806 11744 296812 11756
rect 241480 11716 296812 11744
rect 241480 11704 241486 11716
rect 296806 11704 296812 11716
rect 296864 11704 296870 11756
rect 300762 11704 300768 11756
rect 300820 11744 300826 11756
rect 361574 11744 361580 11756
rect 300820 11716 361580 11744
rect 300820 11704 300826 11716
rect 361574 11704 361580 11716
rect 361632 11704 361638 11756
rect 362218 11704 362224 11756
rect 362276 11744 362282 11756
rect 419534 11744 419540 11756
rect 362276 11716 419540 11744
rect 362276 11704 362282 11716
rect 419534 11704 419540 11716
rect 419592 11704 419598 11756
rect 500862 11704 500868 11756
rect 500920 11744 500926 11756
rect 581086 11744 581092 11756
rect 500920 11716 581092 11744
rect 500920 11704 500926 11716
rect 581086 11704 581092 11716
rect 581144 11704 581150 11756
rect 309778 10344 309784 10396
rect 309836 10384 309842 10396
rect 368474 10384 368480 10396
rect 309836 10356 368480 10384
rect 309836 10344 309842 10356
rect 368474 10344 368480 10356
rect 368532 10344 368538 10396
rect 95142 10276 95148 10328
rect 95200 10316 95206 10328
rect 136634 10316 136640 10328
rect 95200 10288 136640 10316
rect 95200 10276 95206 10288
rect 136634 10276 136640 10288
rect 136692 10276 136698 10328
rect 138658 10276 138664 10328
rect 138716 10316 138722 10328
rect 183646 10316 183652 10328
rect 138716 10288 183652 10316
rect 138716 10276 138722 10288
rect 183646 10276 183652 10288
rect 183704 10276 183710 10328
rect 186222 10276 186228 10328
rect 186280 10316 186286 10328
rect 236086 10316 236092 10328
rect 186280 10288 236092 10316
rect 186280 10276 186286 10288
rect 236086 10276 236092 10288
rect 236144 10276 236150 10328
rect 248322 10276 248328 10328
rect 248380 10316 248386 10328
rect 305086 10316 305092 10328
rect 248380 10288 305092 10316
rect 248380 10276 248386 10288
rect 305086 10276 305092 10288
rect 305144 10276 305150 10328
rect 344922 10276 344928 10328
rect 344980 10316 344986 10328
rect 410794 10316 410800 10328
rect 344980 10288 410800 10316
rect 344980 10276 344986 10288
rect 410794 10276 410800 10288
rect 410852 10276 410858 10328
rect 424962 10276 424968 10328
rect 425020 10316 425026 10328
rect 497734 10316 497740 10328
rect 425020 10288 497740 10316
rect 425020 10276 425026 10288
rect 497734 10276 497740 10288
rect 497792 10276 497798 10328
rect 499482 10276 499488 10328
rect 499540 10316 499546 10328
rect 579614 10316 579620 10328
rect 499540 10288 579620 10316
rect 499540 10276 499546 10288
rect 579614 10276 579620 10288
rect 579672 10276 579678 10328
rect 369857 9707 369915 9713
rect 369857 9673 369869 9707
rect 369903 9704 369915 9707
rect 370406 9704 370412 9716
rect 369903 9676 370412 9704
rect 369903 9673 369915 9676
rect 369857 9667 369915 9673
rect 370406 9664 370412 9676
rect 370464 9664 370470 9716
rect 378137 9707 378195 9713
rect 378137 9673 378149 9707
rect 378183 9704 378195 9707
rect 378778 9704 378784 9716
rect 378183 9676 378784 9704
rect 378183 9673 378195 9676
rect 378137 9667 378195 9673
rect 378778 9664 378784 9676
rect 378836 9664 378842 9716
rect 397457 9707 397515 9713
rect 397457 9673 397469 9707
rect 397503 9704 397515 9707
rect 397822 9704 397828 9716
rect 397503 9676 397828 9704
rect 397503 9673 397515 9676
rect 397457 9667 397515 9673
rect 397822 9664 397828 9676
rect 397880 9664 397886 9716
rect 415397 9707 415455 9713
rect 415397 9673 415409 9707
rect 415443 9704 415455 9707
rect 415670 9704 415676 9716
rect 415443 9676 415676 9704
rect 415443 9673 415455 9676
rect 415397 9667 415455 9673
rect 415670 9664 415676 9676
rect 415728 9664 415734 9716
rect 561677 9707 561735 9713
rect 561677 9673 561689 9707
rect 561723 9704 561735 9707
rect 561950 9704 561956 9716
rect 561723 9676 561956 9704
rect 561723 9673 561735 9676
rect 561677 9667 561735 9673
rect 561950 9664 561956 9676
rect 562008 9664 562014 9716
rect 353754 9596 353760 9648
rect 353812 9596 353818 9648
rect 354950 9596 354956 9648
rect 355008 9596 355014 9648
rect 389450 9596 389456 9648
rect 389508 9596 389514 9648
rect 395430 9596 395436 9648
rect 395488 9596 395494 9648
rect 495434 9596 495440 9648
rect 495492 9636 495498 9648
rect 496541 9639 496599 9645
rect 496541 9636 496553 9639
rect 495492 9608 496553 9636
rect 495492 9596 495498 9608
rect 496541 9605 496553 9608
rect 496587 9605 496599 9639
rect 496541 9599 496599 9605
rect 353772 9512 353800 9596
rect 354968 9512 354996 9596
rect 389468 9512 389496 9596
rect 395448 9512 395476 9596
rect 353754 9460 353760 9512
rect 353812 9460 353818 9512
rect 354950 9460 354956 9512
rect 355008 9460 355014 9512
rect 389450 9460 389456 9512
rect 389508 9460 389514 9512
rect 395430 9460 395436 9512
rect 395488 9460 395494 9512
rect 88242 8916 88248 8968
rect 88300 8956 88306 8968
rect 130194 8956 130200 8968
rect 88300 8928 130200 8956
rect 88300 8916 88306 8928
rect 130194 8916 130200 8928
rect 130252 8916 130258 8968
rect 131022 8916 131028 8968
rect 131080 8956 131086 8968
rect 176562 8956 176568 8968
rect 131080 8928 176568 8956
rect 131080 8916 131086 8928
rect 176562 8916 176568 8928
rect 176620 8916 176626 8968
rect 179322 8916 179328 8968
rect 179380 8956 179386 8968
rect 230106 8956 230112 8968
rect 179380 8928 230112 8956
rect 179380 8916 179386 8928
rect 230106 8916 230112 8928
rect 230164 8916 230170 8968
rect 245562 8916 245568 8968
rect 245620 8956 245626 8968
rect 301406 8956 301412 8968
rect 245620 8928 301412 8956
rect 245620 8916 245626 8928
rect 301406 8916 301412 8928
rect 301464 8916 301470 8968
rect 303522 8916 303528 8968
rect 303580 8956 303586 8968
rect 365806 8956 365812 8968
rect 303580 8928 365812 8956
rect 303580 8916 303586 8928
rect 365806 8916 365812 8928
rect 365864 8916 365870 8968
rect 369762 8916 369768 8968
rect 369820 8956 369826 8968
rect 437014 8956 437020 8968
rect 369820 8928 437020 8956
rect 369820 8916 369826 8928
rect 437014 8916 437020 8928
rect 437072 8916 437078 8968
rect 438118 8916 438124 8968
rect 438176 8956 438182 8968
rect 486970 8956 486976 8968
rect 438176 8928 486976 8956
rect 438176 8916 438182 8928
rect 486970 8916 486976 8928
rect 487028 8916 487034 8968
rect 487062 8916 487068 8968
rect 487120 8956 487126 8968
rect 565538 8956 565544 8968
rect 487120 8928 565544 8956
rect 487120 8916 487126 8928
rect 565538 8916 565544 8928
rect 565596 8916 565602 8968
rect 410886 8412 410892 8424
rect 410847 8384 410892 8412
rect 410886 8372 410892 8384
rect 410944 8372 410950 8424
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 79318 8276 79324 8288
rect 3476 8248 79324 8276
rect 3476 8236 3482 8248
rect 79318 8236 79324 8248
rect 79376 8236 79382 8288
rect 410886 8276 410892 8288
rect 410847 8248 410892 8276
rect 410886 8236 410892 8248
rect 410944 8236 410950 8288
rect 86862 7624 86868 7676
rect 86920 7664 86926 7676
rect 128906 7664 128912 7676
rect 86920 7636 128912 7664
rect 86920 7624 86926 7636
rect 128906 7624 128912 7636
rect 128964 7624 128970 7676
rect 358722 7624 358728 7676
rect 358780 7664 358786 7676
rect 426342 7664 426348 7676
rect 358780 7636 426348 7664
rect 358780 7624 358786 7636
rect 426342 7624 426348 7636
rect 426400 7624 426406 7676
rect 124122 7556 124128 7608
rect 124180 7596 124186 7608
rect 169386 7596 169392 7608
rect 124180 7568 169392 7596
rect 124180 7556 124186 7568
rect 169386 7556 169392 7568
rect 169444 7556 169450 7608
rect 176378 7556 176384 7608
rect 176436 7596 176442 7608
rect 226518 7596 226524 7608
rect 176436 7568 226524 7596
rect 176436 7556 176442 7568
rect 226518 7556 226524 7568
rect 226576 7556 226582 7608
rect 238662 7556 238668 7608
rect 238720 7596 238726 7608
rect 294322 7596 294328 7608
rect 238720 7568 294328 7596
rect 238720 7556 238726 7568
rect 294322 7556 294328 7568
rect 294380 7556 294386 7608
rect 298002 7556 298008 7608
rect 298060 7596 298066 7608
rect 298060 7568 354536 7596
rect 298060 7556 298066 7568
rect 354508 7528 354536 7568
rect 356054 7556 356060 7608
rect 356112 7596 356118 7608
rect 357342 7596 357348 7608
rect 356112 7568 357348 7596
rect 356112 7556 356118 7568
rect 357342 7556 357348 7568
rect 357400 7556 357406 7608
rect 373994 7556 374000 7608
rect 374052 7596 374058 7608
rect 375190 7596 375196 7608
rect 374052 7568 375196 7596
rect 374052 7556 374058 7568
rect 375190 7556 375196 7568
rect 375248 7556 375254 7608
rect 390554 7556 390560 7608
rect 390612 7596 390618 7608
rect 391842 7596 391848 7608
rect 390612 7568 391848 7596
rect 390612 7556 390618 7568
rect 391842 7556 391848 7568
rect 391900 7556 391906 7608
rect 416774 7556 416780 7608
rect 416832 7596 416838 7608
rect 417970 7596 417976 7608
rect 416832 7568 417976 7596
rect 416832 7556 416838 7568
rect 417970 7556 417976 7568
rect 418028 7556 418034 7608
rect 420822 7556 420828 7608
rect 420880 7596 420886 7608
rect 494146 7596 494152 7608
rect 420880 7568 494152 7596
rect 420880 7556 420886 7568
rect 494146 7556 494152 7568
rect 494204 7556 494210 7608
rect 496722 7556 496728 7608
rect 496780 7596 496786 7608
rect 576210 7596 576216 7608
rect 496780 7568 576216 7596
rect 496780 7556 496786 7568
rect 576210 7556 576216 7568
rect 576268 7556 576274 7608
rect 358538 7528 358544 7540
rect 354508 7500 358544 7528
rect 358538 7488 358544 7500
rect 358596 7488 358602 7540
rect 121362 6196 121368 6248
rect 121420 6236 121426 6248
rect 165890 6236 165896 6248
rect 121420 6208 165896 6236
rect 121420 6196 121426 6208
rect 165890 6196 165896 6208
rect 165948 6196 165954 6248
rect 160002 6128 160008 6180
rect 160060 6168 160066 6180
rect 208670 6168 208676 6180
rect 160060 6140 208676 6168
rect 160060 6128 160066 6140
rect 208670 6128 208676 6140
rect 208728 6128 208734 6180
rect 219342 6128 219348 6180
rect 219400 6168 219406 6180
rect 272886 6168 272892 6180
rect 219400 6140 272892 6168
rect 219400 6128 219406 6140
rect 272886 6128 272892 6140
rect 272944 6128 272950 6180
rect 274542 6128 274548 6180
rect 274600 6168 274606 6180
rect 333606 6168 333612 6180
rect 274600 6140 333612 6168
rect 274600 6128 274606 6140
rect 333606 6128 333612 6140
rect 333664 6128 333670 6180
rect 336642 6128 336648 6180
rect 336700 6168 336706 6180
rect 401318 6168 401324 6180
rect 336700 6140 401324 6168
rect 336700 6128 336706 6140
rect 401318 6128 401324 6140
rect 401376 6128 401382 6180
rect 410889 6171 410947 6177
rect 410889 6137 410901 6171
rect 410935 6168 410947 6171
rect 483474 6168 483480 6180
rect 410935 6140 483480 6168
rect 410935 6137 410947 6140
rect 410889 6131 410947 6137
rect 483474 6128 483480 6140
rect 483532 6128 483538 6180
rect 489822 6128 489828 6180
rect 489880 6168 489886 6180
rect 569034 6168 569040 6180
rect 489880 6140 569040 6168
rect 489880 6128 489886 6140
rect 569034 6128 569040 6140
rect 569092 6128 569098 6180
rect 502978 5448 502984 5500
rect 503036 5488 503042 5500
rect 504818 5488 504824 5500
rect 503036 5460 504824 5488
rect 503036 5448 503042 5460
rect 504818 5448 504824 5460
rect 504876 5448 504882 5500
rect 356057 5015 356115 5021
rect 356057 4981 356069 5015
rect 356103 5012 356115 5015
rect 365625 5015 365683 5021
rect 365625 5012 365637 5015
rect 356103 4984 365637 5012
rect 356103 4981 356115 4984
rect 356057 4975 356115 4981
rect 365625 4981 365637 4984
rect 365671 4981 365683 5015
rect 365625 4975 365683 4981
rect 365717 5015 365775 5021
rect 365717 4981 365729 5015
rect 365763 5012 365775 5015
rect 370501 5015 370559 5021
rect 370501 5012 370513 5015
rect 365763 4984 370513 5012
rect 365763 4981 365775 4984
rect 365717 4975 365775 4981
rect 370501 4981 370513 4984
rect 370547 4981 370559 5015
rect 370501 4975 370559 4981
rect 231118 4836 231124 4888
rect 231176 4876 231182 4888
rect 265802 4876 265808 4888
rect 231176 4848 265808 4876
rect 231176 4836 231182 4848
rect 265802 4836 265808 4848
rect 265860 4836 265866 4888
rect 353202 4836 353208 4888
rect 353260 4876 353266 4888
rect 356057 4879 356115 4885
rect 356057 4876 356069 4879
rect 353260 4848 356069 4876
rect 353260 4836 353266 4848
rect 356057 4845 356069 4848
rect 356103 4845 356115 4879
rect 356057 4839 356115 4845
rect 365717 4879 365775 4885
rect 365717 4845 365729 4879
rect 365763 4845 365775 4879
rect 365717 4839 365775 4845
rect 370501 4879 370559 4885
rect 370501 4845 370513 4879
rect 370547 4876 370559 4879
rect 419166 4876 419172 4888
rect 370547 4848 376800 4876
rect 370547 4845 370559 4848
rect 370501 4839 370559 4845
rect 85482 4768 85488 4820
rect 85540 4808 85546 4820
rect 126606 4808 126612 4820
rect 85540 4780 126612 4808
rect 85540 4768 85546 4780
rect 126606 4768 126612 4780
rect 126664 4768 126670 4820
rect 128998 4768 129004 4820
rect 129056 4808 129062 4820
rect 172974 4808 172980 4820
rect 129056 4780 172980 4808
rect 129056 4768 129062 4780
rect 172974 4768 172980 4780
rect 173032 4768 173038 4820
rect 173802 4768 173808 4820
rect 173860 4808 173866 4820
rect 222930 4808 222936 4820
rect 173860 4780 222936 4808
rect 173860 4768 173866 4780
rect 222930 4768 222936 4780
rect 222988 4768 222994 4820
rect 264882 4768 264888 4820
rect 264940 4808 264946 4820
rect 322842 4808 322848 4820
rect 264940 4780 322848 4808
rect 264940 4768 264946 4780
rect 322842 4768 322848 4780
rect 322900 4768 322906 4820
rect 323578 4768 323584 4820
rect 323636 4808 323642 4820
rect 347866 4808 347872 4820
rect 323636 4780 347872 4808
rect 323636 4768 323642 4780
rect 347866 4768 347872 4780
rect 347924 4768 347930 4820
rect 365625 4811 365683 4817
rect 365625 4777 365637 4811
rect 365671 4808 365683 4811
rect 365732 4808 365760 4839
rect 376772 4817 376800 4848
rect 391216 4848 419172 4876
rect 365671 4780 365760 4808
rect 376757 4811 376815 4817
rect 365671 4777 365683 4780
rect 365625 4771 365683 4777
rect 376757 4777 376769 4811
rect 376803 4777 376815 4811
rect 376757 4771 376815 4777
rect 376849 4811 376907 4817
rect 376849 4777 376861 4811
rect 376895 4808 376907 4811
rect 391216 4808 391244 4848
rect 419166 4836 419172 4848
rect 419224 4836 419230 4888
rect 376895 4780 391244 4808
rect 376895 4777 376907 4780
rect 376849 4771 376907 4777
rect 418062 4768 418068 4820
rect 418120 4808 418126 4820
rect 490558 4808 490564 4820
rect 418120 4780 490564 4808
rect 418120 4768 418126 4780
rect 490558 4768 490564 4780
rect 490616 4768 490622 4820
rect 560938 4768 560944 4820
rect 560996 4808 561002 4820
rect 572622 4808 572628 4820
rect 560996 4780 572628 4808
rect 560996 4768 561002 4780
rect 572622 4768 572628 4780
rect 572680 4768 572686 4820
rect 520274 4156 520280 4208
rect 520332 4196 520338 4208
rect 521470 4196 521476 4208
rect 520332 4168 521476 4196
rect 520332 4156 520338 4168
rect 521470 4156 521476 4168
rect 521528 4156 521534 4208
rect 528646 4156 528652 4208
rect 528704 4196 528710 4208
rect 529842 4196 529848 4208
rect 528704 4168 529848 4196
rect 528704 4156 528710 4168
rect 529842 4156 529848 4168
rect 529900 4156 529906 4208
rect 384942 4088 384948 4140
rect 385000 4128 385006 4140
rect 453666 4128 453672 4140
rect 385000 4100 453672 4128
rect 385000 4088 385006 4100
rect 453666 4088 453672 4100
rect 453724 4088 453730 4140
rect 471882 4088 471888 4140
rect 471940 4128 471946 4140
rect 550082 4128 550088 4140
rect 471940 4100 550088 4128
rect 471940 4088 471946 4100
rect 550082 4088 550088 4100
rect 550140 4088 550146 4140
rect 378042 4020 378048 4072
rect 378100 4060 378106 4072
rect 446582 4060 446588 4072
rect 378100 4032 446588 4060
rect 378100 4020 378106 4032
rect 446582 4020 446588 4032
rect 446640 4020 446646 4072
rect 476022 4020 476028 4072
rect 476080 4060 476086 4072
rect 553578 4060 553584 4072
rect 476080 4032 553584 4060
rect 476080 4020 476086 4032
rect 553578 4020 553584 4032
rect 553636 4020 553642 4072
rect 91002 3952 91008 4004
rect 91060 3992 91066 4004
rect 132494 3992 132500 4004
rect 91060 3964 132500 3992
rect 91060 3952 91066 3964
rect 132494 3952 132500 3964
rect 132552 3952 132558 4004
rect 394602 3952 394608 4004
rect 394660 3992 394666 4004
rect 464430 3992 464436 4004
rect 394660 3964 464436 3992
rect 394660 3952 394666 3964
rect 464430 3952 464436 3964
rect 464488 3952 464494 4004
rect 478782 3952 478788 4004
rect 478840 3992 478846 4004
rect 557166 3992 557172 4004
rect 478840 3964 557172 3992
rect 478840 3952 478846 3964
rect 557166 3952 557172 3964
rect 557224 3952 557230 4004
rect 574738 3952 574744 4004
rect 574796 3992 574802 4004
rect 577406 3992 577412 4004
rect 574796 3964 577412 3992
rect 574796 3952 574802 3964
rect 577406 3952 577412 3964
rect 577464 3952 577470 4004
rect 93762 3884 93768 3936
rect 93820 3924 93826 3936
rect 136082 3924 136088 3936
rect 93820 3896 136088 3924
rect 93820 3884 93826 3896
rect 136082 3884 136088 3896
rect 136140 3884 136146 3936
rect 390462 3884 390468 3936
rect 390520 3924 390526 3936
rect 460842 3924 460848 3936
rect 390520 3896 460848 3924
rect 390520 3884 390526 3896
rect 460842 3884 460848 3896
rect 460900 3884 460906 3936
rect 482922 3884 482928 3936
rect 482980 3924 482986 3936
rect 560754 3924 560760 3936
rect 482980 3896 560760 3924
rect 482980 3884 482986 3896
rect 560754 3884 560760 3896
rect 560812 3884 560818 3936
rect 100662 3816 100668 3868
rect 100720 3856 100726 3868
rect 143258 3856 143264 3868
rect 100720 3828 143264 3856
rect 100720 3816 100726 3828
rect 143258 3816 143264 3828
rect 143316 3816 143322 3868
rect 387702 3816 387708 3868
rect 387760 3856 387766 3868
rect 457254 3856 457260 3868
rect 387760 3828 457260 3856
rect 387760 3816 387766 3828
rect 457254 3816 457260 3828
rect 457312 3816 457318 3868
rect 485682 3816 485688 3868
rect 485740 3856 485746 3868
rect 564342 3856 564348 3868
rect 485740 3828 564348 3856
rect 485740 3816 485746 3828
rect 564342 3816 564348 3828
rect 564400 3816 564406 3868
rect 96522 3748 96528 3800
rect 96580 3788 96586 3800
rect 139670 3788 139676 3800
rect 96580 3760 139676 3788
rect 96580 3748 96586 3760
rect 139670 3748 139676 3760
rect 139728 3748 139734 3800
rect 380802 3748 380808 3800
rect 380860 3788 380866 3800
rect 450170 3788 450176 3800
rect 380860 3760 450176 3788
rect 380860 3748 380866 3760
rect 450170 3748 450176 3760
rect 450228 3748 450234 3800
rect 469122 3748 469128 3800
rect 469180 3788 469186 3800
rect 546494 3788 546500 3800
rect 469180 3760 546500 3788
rect 469180 3748 469186 3760
rect 546494 3748 546500 3760
rect 546552 3748 546558 3800
rect 547877 3791 547935 3797
rect 547877 3757 547889 3791
rect 547923 3788 547935 3791
rect 558181 3791 558239 3797
rect 558181 3788 558193 3791
rect 547923 3760 558193 3788
rect 547923 3757 547935 3760
rect 547877 3751 547935 3757
rect 558181 3757 558193 3760
rect 558227 3757 558239 3791
rect 558181 3751 558239 3757
rect 103422 3680 103428 3732
rect 103480 3720 103486 3732
rect 146846 3720 146852 3732
rect 103480 3692 146852 3720
rect 103480 3680 103486 3692
rect 146846 3680 146852 3692
rect 146904 3680 146910 3732
rect 397362 3680 397368 3732
rect 397420 3720 397426 3732
rect 467834 3720 467840 3732
rect 397420 3692 467840 3720
rect 397420 3680 397426 3692
rect 467834 3680 467840 3692
rect 467892 3680 467898 3732
rect 492582 3680 492588 3732
rect 492640 3720 492646 3732
rect 492640 3692 500264 3720
rect 492640 3680 492646 3692
rect 107562 3612 107568 3664
rect 107620 3652 107626 3664
rect 150434 3652 150440 3664
rect 107620 3624 150440 3652
rect 107620 3612 107626 3624
rect 150434 3612 150440 3624
rect 150492 3612 150498 3664
rect 404262 3612 404268 3664
rect 404320 3652 404326 3664
rect 475102 3652 475108 3664
rect 404320 3624 475108 3652
rect 404320 3612 404326 3624
rect 475102 3612 475108 3624
rect 475160 3612 475166 3664
rect 488442 3612 488448 3664
rect 488500 3652 488506 3664
rect 500037 3655 500095 3661
rect 500037 3652 500049 3655
rect 488500 3624 500049 3652
rect 488500 3612 488506 3624
rect 500037 3621 500049 3624
rect 500083 3621 500095 3655
rect 500037 3615 500095 3621
rect 110322 3544 110328 3596
rect 110380 3584 110386 3596
rect 153930 3584 153936 3596
rect 110380 3556 153936 3584
rect 110380 3544 110386 3556
rect 153930 3544 153936 3556
rect 153988 3544 153994 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 218146 3544 218152 3596
rect 218204 3584 218210 3596
rect 219342 3584 219348 3596
rect 218204 3556 219348 3584
rect 218204 3544 218210 3556
rect 219342 3544 219348 3556
rect 219400 3544 219406 3596
rect 227714 3544 227720 3596
rect 227772 3584 227778 3596
rect 228910 3584 228916 3596
rect 227772 3556 228916 3584
rect 227772 3544 227778 3556
rect 228910 3544 228916 3556
rect 228968 3544 228974 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 263410 3584 263416 3596
rect 262272 3556 263416 3584
rect 262272 3544 262278 3556
rect 263410 3544 263416 3556
rect 263468 3544 263474 3596
rect 270494 3544 270500 3596
rect 270552 3584 270558 3596
rect 271690 3584 271696 3596
rect 270552 3556 271696 3584
rect 270552 3544 270558 3556
rect 271690 3544 271696 3556
rect 271748 3544 271754 3596
rect 278866 3544 278872 3596
rect 278924 3584 278930 3596
rect 280062 3584 280068 3596
rect 278924 3556 280068 3584
rect 278924 3544 278930 3556
rect 280062 3544 280068 3556
rect 280120 3544 280126 3596
rect 331214 3544 331220 3596
rect 331272 3584 331278 3596
rect 332410 3584 332416 3596
rect 331272 3556 332416 3584
rect 331272 3544 331278 3556
rect 332410 3544 332416 3556
rect 332468 3544 332474 3596
rect 365714 3544 365720 3596
rect 365772 3584 365778 3596
rect 366910 3584 366916 3596
rect 365772 3556 366916 3584
rect 365772 3544 365778 3556
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 382366 3544 382372 3596
rect 382424 3584 382430 3596
rect 383562 3584 383568 3596
rect 382424 3556 383568 3584
rect 382424 3544 382430 3556
rect 383562 3544 383568 3556
rect 383620 3544 383626 3596
rect 400122 3544 400128 3596
rect 400180 3584 400186 3596
rect 471514 3584 471520 3596
rect 400180 3556 471520 3584
rect 400180 3544 400186 3556
rect 471514 3544 471520 3556
rect 471572 3544 471578 3596
rect 495250 3544 495256 3596
rect 495308 3584 495314 3596
rect 500236 3584 500264 3692
rect 502242 3680 502248 3732
rect 502300 3720 502306 3732
rect 582190 3720 582196 3732
rect 502300 3692 582196 3720
rect 502300 3680 502306 3692
rect 582190 3680 582196 3692
rect 582248 3680 582254 3732
rect 500313 3655 500371 3661
rect 500313 3621 500325 3655
rect 500359 3652 500371 3655
rect 547877 3655 547935 3661
rect 547877 3652 547889 3655
rect 500359 3624 547889 3652
rect 500359 3621 500371 3624
rect 500313 3615 500371 3621
rect 547877 3621 547889 3624
rect 547923 3621 547935 3655
rect 547877 3615 547935 3621
rect 558181 3655 558239 3661
rect 558181 3621 558193 3655
rect 558227 3652 558239 3655
rect 567194 3652 567200 3664
rect 558227 3624 567200 3652
rect 558227 3621 558239 3624
rect 558181 3615 558239 3621
rect 567194 3612 567200 3624
rect 567252 3612 567258 3664
rect 571426 3584 571432 3596
rect 495308 3556 495664 3584
rect 500236 3556 571432 3584
rect 495308 3544 495314 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 81434 3516 81440 3528
rect 624 3488 81440 3516
rect 624 3476 630 3488
rect 81434 3476 81440 3488
rect 81492 3476 81498 3528
rect 117222 3476 117228 3528
rect 117280 3516 117286 3528
rect 117280 3488 157656 3516
rect 117280 3476 117286 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 82814 3448 82820 3460
rect 1728 3420 82820 3448
rect 1728 3408 1734 3420
rect 82814 3408 82820 3420
rect 82872 3408 82878 3460
rect 113082 3408 113088 3460
rect 113140 3448 113146 3460
rect 157518 3448 157524 3460
rect 113140 3420 157524 3448
rect 113140 3408 113146 3420
rect 157518 3408 157524 3420
rect 157576 3408 157582 3460
rect 157628 3448 157656 3488
rect 158714 3476 158720 3528
rect 158772 3516 158778 3528
rect 159910 3516 159916 3528
rect 158772 3488 159916 3516
rect 158772 3476 158778 3488
rect 159910 3476 159916 3488
rect 159968 3476 159974 3528
rect 166994 3476 167000 3528
rect 167052 3516 167058 3528
rect 168190 3516 168196 3528
rect 167052 3488 168196 3516
rect 167052 3476 167058 3488
rect 168190 3476 168196 3488
rect 168248 3476 168254 3528
rect 183554 3476 183560 3528
rect 183612 3516 183618 3528
rect 184842 3516 184848 3528
rect 183612 3488 184848 3516
rect 183612 3476 183618 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 211062 3516 211068 3528
rect 209832 3488 211068 3516
rect 209832 3476 209838 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 252554 3476 252560 3528
rect 252612 3516 252618 3528
rect 253842 3516 253848 3528
rect 252612 3488 253848 3516
rect 252612 3476 252618 3488
rect 253842 3476 253848 3488
rect 253900 3476 253906 3528
rect 287146 3476 287152 3528
rect 287204 3516 287210 3528
rect 288342 3516 288348 3528
rect 287204 3488 288348 3516
rect 287204 3476 287210 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 304994 3476 305000 3528
rect 305052 3516 305058 3528
rect 306190 3516 306196 3528
rect 305052 3488 306196 3516
rect 305052 3476 305058 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 313274 3476 313280 3528
rect 313332 3516 313338 3528
rect 314562 3516 314568 3528
rect 313332 3488 314568 3516
rect 313332 3476 313338 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 347774 3476 347780 3528
rect 347832 3516 347838 3528
rect 349062 3516 349068 3528
rect 347832 3488 349068 3516
rect 347832 3476 347838 3488
rect 349062 3476 349068 3488
rect 349120 3476 349126 3528
rect 411162 3476 411168 3528
rect 411220 3516 411226 3528
rect 482278 3516 482284 3528
rect 411220 3488 482284 3516
rect 411220 3476 411226 3488
rect 482278 3476 482284 3488
rect 482336 3476 482342 3528
rect 494054 3476 494060 3528
rect 494112 3516 494118 3528
rect 495342 3516 495348 3528
rect 494112 3488 495348 3516
rect 494112 3476 494118 3488
rect 495342 3476 495348 3488
rect 495400 3476 495406 3528
rect 495636 3516 495664 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 575014 3516 575020 3528
rect 495636 3488 575020 3516
rect 575014 3476 575020 3488
rect 575072 3476 575078 3528
rect 161106 3448 161112 3460
rect 157628 3420 161112 3448
rect 161106 3408 161112 3420
rect 161164 3408 161170 3460
rect 407022 3408 407028 3460
rect 407080 3448 407086 3460
rect 478690 3448 478696 3460
rect 407080 3420 478696 3448
rect 407080 3408 407086 3420
rect 478690 3408 478696 3420
rect 478748 3408 478754 3460
rect 498102 3408 498108 3460
rect 498160 3448 498166 3460
rect 578602 3448 578608 3460
rect 498160 3420 578608 3448
rect 498160 3408 498166 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 132586 3340 132592 3392
rect 132644 3380 132650 3392
rect 133782 3380 133788 3392
rect 132644 3352 133788 3380
rect 132644 3340 132650 3352
rect 133782 3340 133788 3352
rect 133840 3340 133846 3392
rect 433334 3340 433340 3392
rect 433392 3380 433398 3392
rect 434622 3380 434628 3392
rect 433392 3352 434628 3380
rect 433392 3340 433398 3352
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 451274 3340 451280 3392
rect 451332 3380 451338 3392
rect 452470 3380 452476 3392
rect 451332 3352 452476 3380
rect 451332 3340 451338 3352
rect 452470 3340 452476 3352
rect 452528 3340 452534 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 511994 3340 512000 3392
rect 512052 3380 512058 3392
rect 513190 3380 513196 3392
rect 512052 3352 513196 3380
rect 512052 3340 512058 3352
rect 513190 3340 513196 3352
rect 513248 3340 513254 3392
rect 536834 3340 536840 3392
rect 536892 3380 536898 3392
rect 538122 3380 538128 3392
rect 536892 3352 538128 3380
rect 536892 3340 536898 3352
rect 538122 3340 538128 3352
rect 538180 3340 538186 3392
rect 567194 3340 567200 3392
rect 567252 3380 567258 3392
rect 567838 3380 567844 3392
rect 567252 3352 567844 3380
rect 567252 3340 567258 3352
rect 567838 3340 567844 3352
rect 567896 3340 567902 3392
rect 140774 3000 140780 3052
rect 140832 3040 140838 3052
rect 142062 3040 142068 3052
rect 140832 3012 142068 3040
rect 140832 3000 140838 3012
rect 142062 3000 142068 3012
rect 142120 3000 142126 3052
rect 498194 2796 498200 2848
rect 498252 2836 498258 2848
rect 498252 2808 498976 2836
rect 498252 2796 498258 2808
rect 498948 2780 498976 2808
rect 499574 2796 499580 2848
rect 499632 2836 499638 2848
rect 499632 2808 500172 2836
rect 499632 2796 499638 2808
rect 500144 2780 500172 2808
rect 498930 2728 498936 2780
rect 498988 2728 498994 2780
rect 500126 2728 500132 2780
rect 500184 2728 500190 2780
rect 502334 2048 502340 2100
rect 502392 2088 502398 2100
rect 503622 2088 503628 2100
rect 502392 2060 503628 2088
rect 502392 2048 502398 2060
rect 503622 2048 503628 2060
rect 503680 2048 503686 2100
rect 126974 552 126980 604
rect 127032 592 127038 604
rect 127802 592 127808 604
rect 127032 564 127808 592
rect 127032 552 127038 564
rect 127802 552 127808 564
rect 127860 552 127866 604
rect 131114 552 131120 604
rect 131172 592 131178 604
rect 131390 592 131396 604
rect 131172 564 131396 592
rect 131172 552 131178 564
rect 131390 552 131396 564
rect 131448 552 131454 604
rect 496538 592 496544 604
rect 496499 564 496544 592
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 579614 552 579620 604
rect 579672 592 579678 604
rect 579798 592 579804 604
rect 579672 564 579804 592
rect 579672 552 579678 564
rect 579798 552 579804 564
rect 579856 552 579862 604
<< via1 >>
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 331220 697552 331272 697604
rect 332508 697552 332560 697604
rect 538864 696940 538916 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 694084 72752 694136
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 347780 692792 347832 692844
rect 348884 692792 348936 692844
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 412824 692724 412876 692776
rect 542544 692724 542596 692776
rect 542728 692724 542780 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 429200 684428 429252 684480
rect 429844 684428 429896 684480
rect 558920 684428 558972 684480
rect 559656 684428 559708 684480
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 412640 683068 412692 683120
rect 429200 683068 429252 683120
rect 542360 683068 542412 683120
rect 558920 683068 558972 683120
rect 3792 681708 3844 681760
rect 32404 681708 32456 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 347780 673480 347832 673532
rect 347964 673480 348016 673532
rect 364340 673480 364392 673532
rect 364524 673480 364576 673532
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 494060 673480 494112 673532
rect 494244 673480 494296 673532
rect 536104 673480 536156 673532
rect 580172 673480 580224 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 219072 666544 219124 666596
rect 413100 666544 413152 666596
rect 429660 666544 429712 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 73068 656820 73120 656872
rect 219348 656820 219400 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 284024 654100 284076 654152
rect 284208 654100 284260 654152
rect 347780 654100 347832 654152
rect 347964 654100 348016 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 10324 652740 10376 652792
rect 529204 650020 529256 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 72976 640364 73028 640416
rect 219256 640364 219308 640416
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 72792 640228 72844 640280
rect 219072 640228 219124 640280
rect 72792 637551 72844 637560
rect 72792 637517 72801 637551
rect 72801 637517 72835 637551
rect 72835 637517 72844 637551
rect 72792 637508 72844 637517
rect 219072 637551 219124 637560
rect 219072 637517 219081 637551
rect 219081 637517 219115 637551
rect 219115 637517 219124 637551
rect 219072 637508 219124 637517
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 284024 634788 284076 634840
rect 284208 634788 284260 634840
rect 347780 634788 347832 634840
rect 347964 634788 348016 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 73068 627920 73120 627972
rect 219348 627920 219400 627972
rect 571984 626560 572036 626612
rect 580172 626560 580224 626612
rect 3240 623772 3292 623824
rect 8944 623772 8996 623824
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 284024 615476 284076 615528
rect 284208 615476 284260 615528
rect 347780 615476 347832 615528
rect 347964 615476 348016 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 477500 615476 477552 615528
rect 477684 615476 477736 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 300768 604392 300820 604444
rect 307484 604392 307536 604444
rect 89628 603984 89680 604036
rect 151912 603984 151964 604036
rect 73068 603916 73120 603968
rect 136364 603916 136416 603968
rect 41328 603848 41380 603900
rect 120816 603848 120868 603900
rect 154304 603848 154356 603900
rect 198556 603848 198608 603900
rect 385224 603848 385276 603900
rect 412732 603848 412784 603900
rect 447416 603848 447468 603900
rect 494244 603848 494296 603900
rect 494336 603848 494388 603900
rect 559012 603848 559064 603900
rect 24768 603780 24820 603832
rect 105268 603780 105320 603832
rect 137744 603780 137796 603832
rect 183008 603780 183060 603832
rect 202788 603780 202840 603832
rect 229652 603780 229704 603832
rect 235908 603780 235960 603832
rect 260748 603780 260800 603832
rect 400772 603780 400824 603832
rect 429292 603780 429344 603832
rect 431868 603780 431920 603832
rect 477684 603780 477736 603832
rect 478512 603780 478564 603832
rect 542452 603780 542504 603832
rect 8024 603712 8076 603764
rect 89720 603712 89772 603764
rect 106188 603712 106240 603764
rect 167460 603712 167512 603764
rect 171048 603712 171100 603764
rect 214104 603712 214156 603764
rect 219348 603712 219400 603764
rect 245200 603712 245252 603764
rect 267648 603712 267700 603764
rect 276296 603712 276348 603764
rect 284024 603712 284076 603764
rect 291844 603712 291896 603764
rect 323032 603712 323084 603764
rect 331220 603712 331272 603764
rect 338580 603712 338632 603764
rect 347964 603712 348016 603764
rect 354128 603712 354180 603764
rect 364524 603712 364576 603764
rect 369676 603712 369728 603764
rect 397460 603712 397512 603764
rect 416320 603712 416372 603764
rect 462320 603712 462372 603764
rect 462964 603712 463016 603764
rect 527180 603712 527232 603764
rect 565084 603100 565136 603152
rect 580172 603100 580224 603152
rect 505008 597456 505060 597508
rect 538864 597456 538916 597508
rect 32404 596096 32456 596148
rect 78680 596096 78732 596148
rect 3332 594804 3384 594856
rect 13084 594804 13136 594856
rect 507124 592016 507176 592068
rect 579896 592016 579948 592068
rect 504640 586440 504692 586492
rect 580264 586440 580316 586492
rect 3424 585080 3476 585132
rect 78680 585080 78732 585132
rect 511264 579640 511316 579692
rect 580172 579640 580224 579692
rect 505008 573996 505060 574048
rect 536104 573996 536156 574048
rect 10324 572636 10376 572688
rect 78680 572636 78732 572688
rect 3424 567196 3476 567248
rect 10324 567196 10376 567248
rect 505008 562980 505060 563032
rect 529204 562980 529256 563032
rect 8944 560192 8996 560244
rect 78680 560192 78732 560244
rect 504364 556180 504416 556232
rect 580172 556180 580224 556232
rect 505008 551964 505060 552016
rect 580356 551964 580408 552016
rect 3516 549176 3568 549228
rect 78680 549176 78732 549228
rect 505008 540880 505060 540932
rect 571984 540880 572036 540932
rect 13084 536732 13136 536784
rect 78680 536732 78732 536784
rect 505744 532720 505796 532772
rect 580172 532720 580224 532772
rect 505008 529864 505060 529916
rect 565084 529864 565136 529916
rect 10324 525716 10376 525768
rect 78680 525716 78732 525768
rect 504180 518508 504232 518560
rect 507124 518508 507176 518560
rect 3424 513272 3476 513324
rect 78680 513272 78732 513324
rect 507124 509260 507176 509312
rect 580172 509260 580224 509312
rect 505008 507696 505060 507748
rect 511264 507696 511316 507748
rect 3516 500896 3568 500948
rect 78680 500896 78732 500948
rect 3424 489812 3476 489864
rect 78680 489812 78732 489864
rect 504364 485800 504416 485852
rect 580172 485800 580224 485852
rect 505008 485732 505060 485784
rect 580264 485732 580316 485784
rect 3516 477436 3568 477488
rect 78680 477436 78732 477488
rect 503720 474308 503772 474360
rect 505744 474308 505796 474360
rect 3424 464992 3476 465044
rect 78680 464992 78732 465044
rect 503812 463632 503864 463684
rect 507124 463632 507176 463684
rect 3424 452548 3476 452600
rect 78680 452548 78732 452600
rect 504180 452548 504232 452600
rect 580356 452548 580408 452600
rect 504364 438880 504416 438932
rect 580172 438880 580224 438932
rect 3148 438812 3200 438864
rect 78680 438812 78732 438864
rect 505008 430516 505060 430568
rect 580264 430516 580316 430568
rect 3240 425008 3292 425060
rect 78680 425008 78732 425060
rect 505008 419432 505060 419484
rect 580448 419432 580500 419484
rect 505008 397400 505060 397452
rect 580356 397400 580408 397452
rect 3148 395972 3200 396024
rect 79324 395972 79376 396024
rect 504548 386316 504600 386368
rect 580264 386316 580316 386368
rect 3240 380808 3292 380860
rect 79416 380808 79468 380860
rect 505008 375300 505060 375352
rect 580356 375300 580408 375352
rect 3148 367004 3200 367056
rect 79324 367004 79376 367056
rect 505008 362856 505060 362908
rect 580264 362856 580316 362908
rect 504640 353200 504692 353252
rect 580264 353200 580316 353252
rect 505008 340824 505060 340876
rect 580908 340824 580960 340876
rect 3424 338036 3476 338088
rect 79600 338036 79652 338088
rect 3240 324232 3292 324284
rect 79508 324232 79560 324284
rect 504364 322872 504416 322924
rect 580172 322872 580224 322924
rect 503812 311788 503864 311840
rect 580172 311788 580224 311840
rect 3332 309068 3384 309120
rect 79416 309068 79468 309120
rect 504364 299412 504416 299464
rect 579804 299412 579856 299464
rect 3424 295264 3476 295316
rect 79324 295264 79376 295316
rect 3424 280100 3476 280152
rect 79692 280100 79744 280152
rect 504364 275952 504416 276004
rect 580172 275952 580224 276004
rect 10324 273232 10376 273284
rect 78680 273232 78732 273284
rect 3148 266296 3200 266348
rect 79600 266296 79652 266348
rect 504456 264868 504508 264920
rect 580172 264868 580224 264920
rect 3424 252492 3476 252544
rect 79508 252492 79560 252544
rect 504364 252492 504416 252544
rect 579804 252492 579856 252544
rect 25504 238756 25556 238808
rect 78680 238756 78732 238808
rect 3424 237328 3476 237380
rect 79416 237328 79468 237380
rect 504456 229032 504508 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 79324 223524 79376 223576
rect 504732 217948 504784 218000
rect 580172 217948 580224 218000
rect 3424 208292 3476 208344
rect 10324 208292 10376 208344
rect 504364 205572 504416 205624
rect 579804 205572 579856 205624
rect 24124 202852 24176 202904
rect 78680 202852 78732 202904
rect 3148 194488 3200 194540
rect 79600 194488 79652 194540
rect 504548 182112 504600 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 79508 180752 79560 180804
rect 504640 171028 504692 171080
rect 580172 171028 580224 171080
rect 8944 167016 8996 167068
rect 78680 167016 78732 167068
rect 3516 165520 3568 165572
rect 25504 165520 25556 165572
rect 504456 158652 504508 158704
rect 579804 158652 579856 158704
rect 3148 151716 3200 151768
rect 79416 151716 79468 151768
rect 505008 140768 505060 140820
rect 527824 140768 527876 140820
rect 3240 136552 3292 136604
rect 79324 136552 79376 136604
rect 504364 135192 504416 135244
rect 580172 135192 580224 135244
rect 14464 131112 14516 131164
rect 78680 131112 78732 131164
rect 504824 124108 504876 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 24124 122748 24176 122800
rect 504732 111732 504784 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 79784 108944 79836 108996
rect 504272 106292 504324 106344
rect 571984 106292 572036 106344
rect 84568 100648 84620 100700
rect 85488 100648 85540 100700
rect 88892 100648 88944 100700
rect 89628 100648 89680 100700
rect 94412 100648 94464 100700
rect 95148 100648 95200 100700
rect 95424 100648 95476 100700
rect 96436 100648 96488 100700
rect 99840 100648 99892 100700
rect 100668 100648 100720 100700
rect 100944 100648 100996 100700
rect 102784 100648 102836 100700
rect 105268 100648 105320 100700
rect 106188 100648 106240 100700
rect 106372 100648 106424 100700
rect 107568 100648 107620 100700
rect 156420 100648 156472 100700
rect 157248 100648 157300 100700
rect 228180 100648 228232 100700
rect 229008 100648 229060 100700
rect 229284 100648 229336 100700
rect 230388 100648 230440 100700
rect 233608 100648 233660 100700
rect 234528 100648 234580 100700
rect 243452 100648 243504 100700
rect 244188 100648 244240 100700
rect 321744 100648 321796 100700
rect 322756 100648 322808 100700
rect 327172 100648 327224 100700
rect 329104 100648 329156 100700
rect 331588 100648 331640 100700
rect 332508 100648 332560 100700
rect 337016 100648 337068 100700
rect 338028 100648 338080 100700
rect 338120 100648 338172 100700
rect 339316 100648 339368 100700
rect 392492 100648 392544 100700
rect 393228 100648 393280 100700
rect 397920 100648 397972 100700
rect 398748 100648 398800 100700
rect 408776 100648 408828 100700
rect 409788 100648 409840 100700
rect 418620 100648 418672 100700
rect 419448 100648 419500 100700
rect 424048 100648 424100 100700
rect 424968 100648 425020 100700
rect 425152 100648 425204 100700
rect 427084 100648 427136 100700
rect 459928 100648 459980 100700
rect 460848 100648 460900 100700
rect 461032 100648 461084 100700
rect 462964 100648 463016 100700
rect 476304 100648 476356 100700
rect 478236 100648 478288 100700
rect 480628 100648 480680 100700
rect 481548 100648 481600 100700
rect 481732 100648 481784 100700
rect 482928 100648 482980 100700
rect 91100 100580 91152 100632
rect 92388 100580 92440 100632
rect 240140 100580 240192 100632
rect 241336 100580 241388 100632
rect 326160 100512 326212 100564
rect 326988 100512 327040 100564
rect 153108 100444 153160 100496
rect 153844 100444 153896 100496
rect 295616 100172 295668 100224
rect 296628 100172 296680 100224
rect 301136 100172 301188 100224
rect 302148 100172 302200 100224
rect 211896 100036 211948 100088
rect 231124 100036 231176 100088
rect 286968 100036 287020 100088
rect 323584 100036 323636 100088
rect 325056 100036 325108 100088
rect 337384 100036 337436 100088
rect 353300 100036 353352 100088
rect 362224 100036 362276 100088
rect 385960 100036 386012 100088
rect 411904 100036 411956 100088
rect 414296 100036 414348 100088
rect 438124 100036 438176 100088
rect 492588 100036 492640 100088
rect 560944 100036 560996 100088
rect 85672 99968 85724 100020
rect 97264 99968 97316 100020
rect 117228 99968 117280 100020
rect 161572 99968 161624 100020
rect 162952 99968 163004 100020
rect 211160 99968 211212 100020
rect 231492 99968 231544 100020
rect 287244 99968 287296 100020
rect 329380 99968 329432 100020
rect 393412 99968 393464 100020
rect 430580 99968 430632 100020
rect 502984 99968 503036 100020
rect 224960 99764 225012 99816
rect 226248 99764 226300 99816
rect 409880 99764 409932 99816
rect 411168 99764 411220 99816
rect 419724 99764 419776 99816
rect 420736 99764 420788 99816
rect 239128 99696 239180 99748
rect 240048 99696 240100 99748
rect 332692 99696 332744 99748
rect 333888 99696 333940 99748
rect 393596 99696 393648 99748
rect 394608 99696 394660 99748
rect 465356 99696 465408 99748
rect 466368 99696 466420 99748
rect 89996 99560 90048 99612
rect 91008 99560 91060 99612
rect 296720 99560 296772 99612
rect 298008 99560 298060 99612
rect 394700 99560 394752 99612
rect 395988 99560 396040 99612
rect 107476 99424 107528 99476
rect 113824 99424 113876 99476
rect 110696 99356 110748 99408
rect 111708 99356 111760 99408
rect 115020 99356 115072 99408
rect 115848 99356 115900 99408
rect 116124 99356 116176 99408
rect 117228 99356 117280 99408
rect 120448 99356 120500 99408
rect 121368 99356 121420 99408
rect 121552 99356 121604 99408
rect 122748 99356 122800 99408
rect 125968 99356 126020 99408
rect 126888 99356 126940 99408
rect 126980 99356 127032 99408
rect 129004 99356 129056 99408
rect 130292 99356 130344 99408
rect 131028 99356 131080 99408
rect 131396 99356 131448 99408
rect 132408 99356 132460 99408
rect 132500 99356 132552 99408
rect 133696 99356 133748 99408
rect 135720 99356 135772 99408
rect 136548 99356 136600 99408
rect 136824 99356 136876 99408
rect 138664 99356 138716 99408
rect 141148 99356 141200 99408
rect 142068 99356 142120 99408
rect 142252 99356 142304 99408
rect 143356 99356 143408 99408
rect 146576 99356 146628 99408
rect 147588 99356 147640 99408
rect 152004 99356 152056 99408
rect 157524 99356 157576 99408
rect 158628 99356 158680 99408
rect 161848 99356 161900 99408
rect 162768 99356 162820 99408
rect 166172 99356 166224 99408
rect 166908 99356 166960 99408
rect 167276 99356 167328 99408
rect 168288 99356 168340 99408
rect 168380 99356 168432 99408
rect 169576 99356 169628 99408
rect 171600 99356 171652 99408
rect 172428 99356 172480 99408
rect 172704 99356 172756 99408
rect 173808 99356 173860 99408
rect 177028 99356 177080 99408
rect 177948 99356 178000 99408
rect 178132 99356 178184 99408
rect 179236 99356 179288 99408
rect 182548 99356 182600 99408
rect 183468 99356 183520 99408
rect 183560 99356 183612 99408
rect 185584 99356 185636 99408
rect 187976 99356 188028 99408
rect 153016 99288 153068 99340
rect 188988 99356 189040 99408
rect 189724 99356 189776 99408
rect 192300 99356 192352 99408
rect 193128 99356 193180 99408
rect 193404 99356 193456 99408
rect 194508 99356 194560 99408
rect 197728 99356 197780 99408
rect 198648 99356 198700 99408
rect 202052 99356 202104 99408
rect 202788 99356 202840 99408
rect 203156 99356 203208 99408
rect 204168 99356 204220 99408
rect 204260 99356 204312 99408
rect 205456 99356 205508 99408
rect 207572 99356 207624 99408
rect 208308 99356 208360 99408
rect 208584 99356 208636 99408
rect 209688 99356 209740 99408
rect 213000 99356 213052 99408
rect 213828 99356 213880 99408
rect 214012 99356 214064 99408
rect 215116 99356 215168 99408
rect 218428 99356 218480 99408
rect 219348 99356 219400 99408
rect 220544 99356 220596 99408
rect 221464 99356 221516 99408
rect 223856 99356 223908 99408
rect 224868 99356 224920 99408
rect 244556 99356 244608 99408
rect 245568 99356 245620 99408
rect 248880 99356 248932 99408
rect 249708 99356 249760 99408
rect 249984 99356 250036 99408
rect 250996 99356 251048 99408
rect 254308 99356 254360 99408
rect 255228 99356 255280 99408
rect 255412 99356 255464 99408
rect 256608 99356 256660 99408
rect 259736 99356 259788 99408
rect 260748 99356 260800 99408
rect 260840 99356 260892 99408
rect 262036 99356 262088 99408
rect 265164 99356 265216 99408
rect 266176 99356 266228 99408
rect 269580 99356 269632 99408
rect 270408 99356 270460 99408
rect 275008 99356 275060 99408
rect 275928 99356 275980 99408
rect 276112 99356 276164 99408
rect 277216 99356 277268 99408
rect 279332 99356 279384 99408
rect 280068 99356 280120 99408
rect 280436 99356 280488 99408
rect 281448 99356 281500 99408
rect 284760 99356 284812 99408
rect 285588 99356 285640 99408
rect 285864 99356 285916 99408
rect 286968 99356 287020 99408
rect 290188 99356 290240 99408
rect 291108 99356 291160 99408
rect 291292 99356 291344 99408
rect 292488 99356 292540 99408
rect 305460 99356 305512 99408
rect 306288 99356 306340 99408
rect 306564 99356 306616 99408
rect 309784 99356 309836 99408
rect 310888 99356 310940 99408
rect 311808 99356 311860 99408
rect 311992 99356 312044 99408
rect 313096 99356 313148 99408
rect 315212 99356 315264 99408
rect 315948 99356 316000 99408
rect 316316 99356 316368 99408
rect 317328 99356 317380 99408
rect 320640 99356 320692 99408
rect 321468 99356 321520 99408
rect 341340 99356 341392 99408
rect 342168 99356 342220 99408
rect 343548 99356 343600 99408
rect 345664 99356 345716 99408
rect 346768 99356 346820 99408
rect 347688 99356 347740 99408
rect 347872 99356 347924 99408
rect 348976 99356 349028 99408
rect 352196 99356 352248 99408
rect 353208 99356 353260 99408
rect 356612 99356 356664 99408
rect 357348 99356 357400 99408
rect 357716 99356 357768 99408
rect 358636 99356 358688 99408
rect 362040 99356 362092 99408
rect 362868 99356 362920 99408
rect 363144 99356 363196 99408
rect 364156 99356 364208 99408
rect 367468 99356 367520 99408
rect 368388 99356 368440 99408
rect 368572 99356 368624 99408
rect 369768 99356 369820 99408
rect 372896 99356 372948 99408
rect 373908 99356 373960 99408
rect 374000 99356 374052 99408
rect 375196 99356 375248 99408
rect 377220 99356 377272 99408
rect 378048 99356 378100 99408
rect 378324 99356 378376 99408
rect 380164 99356 380216 99408
rect 382740 99356 382792 99408
rect 383568 99356 383620 99408
rect 383752 99356 383804 99408
rect 384948 99356 385000 99408
rect 388168 99356 388220 99408
rect 389088 99356 389140 99408
rect 399024 99356 399076 99408
rect 400036 99356 400088 99408
rect 403348 99356 403400 99408
rect 404268 99356 404320 99408
rect 404452 99356 404504 99408
rect 405648 99356 405700 99408
rect 428372 99356 428424 99408
rect 429108 99356 429160 99408
rect 429476 99356 429528 99408
rect 430488 99356 430540 99408
rect 433800 99356 433852 99408
rect 434628 99356 434680 99408
rect 434904 99356 434956 99408
rect 435916 99356 435968 99408
rect 439320 99356 439372 99408
rect 440148 99356 440200 99408
rect 444748 99356 444800 99408
rect 445668 99356 445720 99408
rect 445852 99356 445904 99408
rect 447048 99356 447100 99408
rect 450176 99356 450228 99408
rect 451188 99356 451240 99408
rect 451280 99356 451332 99408
rect 452568 99356 452620 99408
rect 454500 99356 454552 99408
rect 455328 99356 455380 99408
rect 455604 99356 455656 99408
rect 456616 99356 456668 99408
rect 466460 99356 466512 99408
rect 467748 99356 467800 99408
rect 469772 99356 469824 99408
rect 470508 99356 470560 99408
rect 470876 99356 470928 99408
rect 471796 99356 471848 99408
rect 475200 99356 475252 99408
rect 476028 99356 476080 99408
rect 486056 99356 486108 99408
rect 487068 99356 487120 99408
rect 487160 99356 487212 99408
rect 488356 99356 488408 99408
rect 490380 99356 490432 99408
rect 491208 99356 491260 99408
rect 491484 99356 491536 99408
rect 492588 99356 492640 99408
rect 495900 99356 495952 99408
rect 496728 99356 496780 99408
rect 496912 99356 496964 99408
rect 498016 99356 498068 99408
rect 501328 99356 501380 99408
rect 502248 99356 502300 99408
rect 188988 99220 189040 99272
rect 147680 98608 147732 98660
rect 194600 98608 194652 98660
rect 198832 98608 198884 98660
rect 251180 98608 251232 98660
rect 270592 98608 270644 98660
rect 329840 98608 329892 98660
rect 342444 98608 342496 98660
rect 408500 98608 408552 98660
rect 440332 98608 440384 98660
rect 514760 98608 514812 98660
rect 111800 97248 111852 97300
rect 155960 97248 156012 97300
rect 234712 97248 234764 97300
rect 289820 97248 289872 97300
rect 317420 97248 317472 97300
rect 380900 97248 380952 97300
rect 443644 97248 443696 97300
rect 518900 97248 518952 97300
rect 395896 96568 395948 96620
rect 219532 95888 219584 95940
rect 273260 95888 273312 95940
rect 281540 95888 281592 95940
rect 340880 95888 340932 95940
rect 370780 95888 370832 95940
rect 438860 95888 438912 95940
rect 446864 95888 446916 95940
rect 521660 95888 521712 95940
rect 389272 94460 389324 94512
rect 459652 94460 459704 94512
rect 478236 94460 478288 94512
rect 554780 94460 554832 94512
rect 3424 93780 3476 93832
rect 79692 93780 79744 93832
rect 368388 93100 368440 93152
rect 434720 93100 434772 93152
rect 480168 93100 480220 93152
rect 557540 93100 557592 93152
rect 354588 91740 354640 91792
rect 420920 91740 420972 91792
rect 435916 91740 435968 91792
rect 509240 91740 509292 91792
rect 364156 90312 364208 90364
rect 430580 90312 430632 90364
rect 441436 90312 441488 90364
rect 516140 90312 516192 90364
rect 148692 89700 148744 89752
rect 148876 89700 148928 89752
rect 225972 89700 226024 89752
rect 226156 89700 226208 89752
rect 235724 89700 235776 89752
rect 235908 89700 235960 89752
rect 297732 89700 297784 89752
rect 297916 89700 297968 89752
rect 462044 89700 462096 89752
rect 462228 89700 462280 89752
rect 419448 88952 419500 89004
rect 491300 88952 491352 89004
rect 498016 88952 498068 89004
rect 574744 88952 574796 89004
rect 504548 88272 504600 88324
rect 580172 88272 580224 88324
rect 351828 87592 351880 87644
rect 416780 87592 416832 87644
rect 395804 87023 395856 87032
rect 395804 86989 395813 87023
rect 395813 86989 395847 87023
rect 395847 86989 395856 87023
rect 395804 86980 395856 86989
rect 410984 86980 411036 87032
rect 411076 86980 411128 87032
rect 152924 86912 152976 86964
rect 342168 86232 342220 86284
rect 407120 86232 407172 86284
rect 462964 86232 463016 86284
rect 536840 86232 536892 86284
rect 339316 84804 339368 84856
rect 402980 84804 403032 84856
rect 467564 84804 467616 84856
rect 545120 84804 545172 84856
rect 322756 83444 322808 83496
rect 385040 83444 385092 83496
rect 491208 83444 491260 83496
rect 569960 83444 570012 83496
rect 188712 82084 188764 82136
rect 188896 82084 188948 82136
rect 328368 82084 328420 82136
rect 391940 82084 391992 82136
rect 410984 82127 411036 82136
rect 410984 82093 410993 82127
rect 410993 82093 411027 82127
rect 411027 82093 411036 82127
rect 410984 82084 411036 82093
rect 433248 82084 433300 82136
rect 506480 82084 506532 82136
rect 315948 80724 316000 80776
rect 378232 80724 378284 80776
rect 375196 80656 375248 80708
rect 443000 80656 443052 80708
rect 452476 80656 452528 80708
rect 528560 80656 528612 80708
rect 395804 80112 395856 80164
rect 462136 80112 462188 80164
rect 395804 79976 395856 80028
rect 462136 79976 462188 80028
rect 3516 79432 3568 79484
rect 8944 79432 8996 79484
rect 302056 79364 302108 79416
rect 364340 79364 364392 79416
rect 364248 79296 364300 79348
rect 431960 79296 432012 79348
rect 456616 79296 456668 79348
rect 531320 79296 531372 79348
rect 299388 77936 299440 77988
rect 360200 77936 360252 77988
rect 361488 77936 361540 77988
rect 427820 77936 427872 77988
rect 459468 77936 459520 77988
rect 535460 77936 535512 77988
rect 410984 77367 411036 77376
rect 410984 77333 410993 77367
rect 410993 77333 411027 77367
rect 411027 77333 411036 77367
rect 410984 77324 411036 77333
rect 152832 77299 152884 77308
rect 152832 77265 152841 77299
rect 152841 77265 152875 77299
rect 152875 77265 152884 77299
rect 152832 77256 152884 77265
rect 148968 77188 149020 77240
rect 188620 77188 188672 77240
rect 225972 77188 226024 77240
rect 235724 77188 235776 77240
rect 297732 77231 297784 77240
rect 297732 77197 297741 77231
rect 297741 77197 297775 77231
rect 297775 77197 297784 77231
rect 297732 77188 297784 77197
rect 378140 77231 378192 77240
rect 378140 77197 378149 77231
rect 378149 77197 378183 77231
rect 378183 77197 378192 77231
rect 378140 77188 378192 77197
rect 504640 77188 504692 77240
rect 580172 77188 580224 77240
rect 296628 76508 296680 76560
rect 356060 76508 356112 76560
rect 358636 76508 358688 76560
rect 425060 76508 425112 76560
rect 430488 76508 430540 76560
rect 502340 76508 502392 76560
rect 260748 75148 260800 75200
rect 317420 75148 317472 75200
rect 318708 75148 318760 75200
rect 382280 75148 382332 75200
rect 426348 75148 426400 75200
rect 499580 75148 499632 75200
rect 256516 73856 256568 73908
rect 313280 73856 313332 73908
rect 313096 73788 313148 73840
rect 374000 73788 374052 73840
rect 423588 73788 423640 73840
rect 495440 73788 495492 73840
rect 246948 72428 247000 72480
rect 303620 72428 303672 72480
rect 309048 72428 309100 72480
rect 371240 72428 371292 72480
rect 420736 72428 420788 72480
rect 492680 72428 492732 72480
rect 280068 71068 280120 71120
rect 339500 71068 339552 71120
rect 224868 71000 224920 71052
rect 278780 71000 278832 71052
rect 335268 71000 335320 71052
rect 400220 71000 400272 71052
rect 409788 71000 409840 71052
rect 480260 71000 480312 71052
rect 153016 70388 153068 70440
rect 410892 70388 410944 70440
rect 152924 70252 152976 70304
rect 410984 70252 411036 70304
rect 230296 69640 230348 69692
rect 285680 69640 285732 69692
rect 286968 69640 287020 69692
rect 346400 69640 346452 69692
rect 405556 69640 405608 69692
rect 477592 69640 477644 69692
rect 215116 68280 215168 68332
rect 267740 68280 267792 68332
rect 273168 68280 273220 68332
rect 331220 68280 331272 68332
rect 332508 68280 332560 68332
rect 396080 68280 396132 68332
rect 402888 68280 402940 68332
rect 473360 68280 473412 68332
rect 378140 67711 378192 67720
rect 378140 67677 378149 67711
rect 378149 67677 378183 67711
rect 378183 67677 378192 67711
rect 378140 67668 378192 67677
rect 148876 67643 148928 67652
rect 148876 67609 148885 67643
rect 148885 67609 148919 67643
rect 148919 67609 148928 67643
rect 148876 67600 148928 67609
rect 188528 67643 188580 67652
rect 188528 67609 188537 67643
rect 188537 67609 188571 67643
rect 188571 67609 188580 67643
rect 188528 67600 188580 67609
rect 225880 67643 225932 67652
rect 225880 67609 225889 67643
rect 225889 67609 225923 67643
rect 225923 67609 225932 67643
rect 225880 67600 225932 67609
rect 235632 67643 235684 67652
rect 235632 67609 235641 67643
rect 235641 67609 235675 67643
rect 235675 67609 235684 67643
rect 235632 67600 235684 67609
rect 297824 67600 297876 67652
rect 378140 67575 378192 67584
rect 378140 67541 378149 67575
rect 378149 67541 378183 67575
rect 378183 67541 378192 67575
rect 378140 67532 378192 67541
rect 499580 67575 499632 67584
rect 499580 67541 499589 67575
rect 499589 67541 499623 67575
rect 499623 67541 499632 67575
rect 499580 67532 499632 67541
rect 237288 66920 237340 66972
rect 292580 66920 292632 66972
rect 395804 66920 395856 66972
rect 466460 66920 466512 66972
rect 184848 66852 184900 66904
rect 236000 66852 236052 66904
rect 292396 66852 292448 66904
rect 353392 66852 353444 66904
rect 466368 66852 466420 66904
rect 542360 66852 542412 66904
rect 371240 66215 371292 66224
rect 371240 66181 371249 66215
rect 371249 66181 371283 66215
rect 371283 66181 371292 66215
rect 371240 66172 371292 66181
rect 393228 65560 393280 65612
rect 462320 65560 462372 65612
rect 182088 65492 182140 65544
rect 231860 65492 231912 65544
rect 234528 65492 234580 65544
rect 288440 65492 288492 65544
rect 289728 65492 289780 65544
rect 349160 65492 349212 65544
rect 462044 65492 462096 65544
rect 538220 65492 538272 65544
rect 3332 64812 3384 64864
rect 79600 64812 79652 64864
rect 527824 64812 527876 64864
rect 579804 64812 579856 64864
rect 179236 64200 179288 64252
rect 227720 64200 227772 64252
rect 227628 64132 227680 64184
rect 281540 64132 281592 64184
rect 282828 64132 282880 64184
rect 342260 64132 342312 64184
rect 383568 64132 383620 64184
rect 451280 64132 451332 64184
rect 452568 64132 452620 64184
rect 527180 64132 527232 64184
rect 172428 62772 172480 62824
rect 220820 62772 220872 62824
rect 221464 62772 221516 62824
rect 274640 62772 274692 62824
rect 277216 62772 277268 62824
rect 335360 62772 335412 62824
rect 376668 62772 376720 62824
rect 444380 62772 444432 62824
rect 447048 62772 447100 62824
rect 520280 62772 520332 62824
rect 211068 61412 211120 61464
rect 263600 61412 263652 61464
rect 410708 61412 410760 61464
rect 410984 61412 411036 61464
rect 158536 61344 158588 61396
rect 207020 61344 207072 61396
rect 263508 61344 263560 61396
rect 321560 61344 321612 61396
rect 347688 61344 347740 61396
rect 412640 61344 412692 61396
rect 413928 61344 413980 61396
rect 485780 61344 485832 61396
rect 148876 60800 148928 60852
rect 297824 60800 297876 60852
rect 148784 60664 148836 60716
rect 297732 60664 297784 60716
rect 217968 60052 218020 60104
rect 270500 60052 270552 60104
rect 169576 59984 169628 60036
rect 218060 59984 218112 60036
rect 270408 59984 270460 60036
rect 328460 59984 328512 60036
rect 369676 59984 369728 60036
rect 437480 59984 437532 60036
rect 440148 59984 440200 60036
rect 513380 59984 513432 60036
rect 155868 58624 155920 58676
rect 202880 58624 202932 58676
rect 208308 58624 208360 58676
rect 260840 58624 260892 58676
rect 314568 58624 314620 58676
rect 376760 58624 376812 58676
rect 379428 58624 379480 58676
rect 448520 58624 448572 58676
rect 449808 58624 449860 58676
rect 524420 58624 524472 58676
rect 333704 57944 333756 57996
rect 333796 57944 333848 57996
rect 378140 57987 378192 57996
rect 378140 57953 378149 57987
rect 378149 57953 378183 57987
rect 378183 57953 378192 57987
rect 378140 57944 378192 57953
rect 499580 57987 499632 57996
rect 499580 57953 499589 57987
rect 499589 57953 499623 57987
rect 499623 57953 499632 57987
rect 499580 57944 499632 57953
rect 353300 57919 353352 57928
rect 353300 57885 353309 57919
rect 353309 57885 353343 57919
rect 353343 57885 353352 57919
rect 353300 57876 353352 57885
rect 495440 57919 495492 57928
rect 495440 57885 495449 57919
rect 495449 57885 495483 57919
rect 495483 57885 495492 57919
rect 495440 57876 495492 57885
rect 378140 57851 378192 57860
rect 378140 57817 378149 57851
rect 378149 57817 378183 57851
rect 378183 57817 378192 57851
rect 378140 57808 378192 57817
rect 205456 57264 205508 57316
rect 256700 57264 256752 57316
rect 306288 57264 306340 57316
rect 367100 57264 367152 57316
rect 152924 57196 152976 57248
rect 200120 57196 200172 57248
rect 253848 57196 253900 57248
rect 310520 57196 310572 57248
rect 367008 57196 367060 57248
rect 433340 57196 433392 57248
rect 436008 57196 436060 57248
rect 510620 57196 510672 57248
rect 371240 56627 371292 56636
rect 371240 56593 371249 56627
rect 371249 56593 371283 56627
rect 371283 56593 371292 56627
rect 371240 56584 371292 56593
rect 410708 56559 410760 56568
rect 410708 56525 410717 56559
rect 410717 56525 410751 56559
rect 410751 56525 410760 56559
rect 410708 56516 410760 56525
rect 201408 55904 201460 55956
rect 252560 55904 252612 55956
rect 148784 55836 148836 55888
rect 195980 55836 196032 55888
rect 250996 55836 251048 55888
rect 306380 55836 306432 55888
rect 307668 55836 307720 55888
rect 369860 55836 369912 55888
rect 373908 55836 373960 55888
rect 441620 55836 441672 55888
rect 442908 55836 442960 55888
rect 517520 55836 517572 55888
rect 194416 54544 194468 54596
rect 245660 54544 245712 54596
rect 350448 54544 350500 54596
rect 416872 54544 416924 54596
rect 146208 54476 146260 54528
rect 193220 54476 193272 54528
rect 244188 54476 244240 54528
rect 299480 54476 299532 54528
rect 416688 54476 416740 54528
rect 488540 54476 488592 54528
rect 191748 53116 191800 53168
rect 242900 53116 242952 53168
rect 143356 53048 143408 53100
rect 189080 53048 189132 53100
rect 241336 53048 241388 53100
rect 296720 53048 296772 53100
rect 297732 53048 297784 53100
rect 358820 53048 358872 53100
rect 360108 53048 360160 53100
rect 426440 53048 426492 53100
rect 458088 53048 458140 53100
rect 534080 53048 534132 53100
rect 139308 51688 139360 51740
rect 184940 51688 184992 51740
rect 188712 51688 188764 51740
rect 238760 51688 238812 51740
rect 242808 51688 242860 51740
rect 298100 51688 298152 51740
rect 340788 51688 340840 51740
rect 405740 51688 405792 51740
rect 455328 51688 455380 51740
rect 529940 51688 529992 51740
rect 3424 51008 3476 51060
rect 79508 51008 79560 51060
rect 410984 50940 411036 50992
rect 235816 50439 235868 50448
rect 235816 50405 235825 50439
rect 235825 50405 235859 50439
rect 235859 50405 235868 50439
rect 235816 50396 235868 50405
rect 136548 50328 136600 50380
rect 182180 50328 182232 50380
rect 209596 50328 209648 50380
rect 262220 50328 262272 50380
rect 275928 50328 275980 50380
rect 333980 50328 334032 50380
rect 338028 50328 338080 50380
rect 401600 50328 401652 50380
rect 431868 50328 431920 50380
rect 505100 50328 505152 50380
rect 133696 49036 133748 49088
rect 178040 49036 178092 49088
rect 175188 48968 175240 49020
rect 224960 48968 225012 49020
rect 225972 48968 226024 49020
rect 280160 48968 280212 49020
rect 292488 48968 292540 49020
rect 351920 48968 351972 49020
rect 357348 48968 357400 49020
rect 423680 48968 423732 49020
rect 427084 48968 427136 49020
rect 498200 48968 498252 49020
rect 353300 48331 353352 48340
rect 353300 48297 353309 48331
rect 353309 48297 353343 48331
rect 353343 48297 353352 48331
rect 353300 48288 353352 48297
rect 378140 48331 378192 48340
rect 378140 48297 378149 48331
rect 378149 48297 378183 48331
rect 378183 48297 378192 48331
rect 378140 48288 378192 48297
rect 495440 48331 495492 48340
rect 495440 48297 495449 48331
rect 495449 48297 495483 48331
rect 495483 48297 495492 48331
rect 495440 48288 495492 48297
rect 333796 48195 333848 48204
rect 333796 48161 333805 48195
rect 333805 48161 333839 48195
rect 333839 48161 333848 48195
rect 333796 48152 333848 48161
rect 164148 47540 164200 47592
rect 212540 47540 212592 47592
rect 213828 47540 213880 47592
rect 266360 47540 266412 47592
rect 271696 47540 271748 47592
rect 331312 47540 331364 47592
rect 398840 47540 398892 47592
rect 400036 47540 400088 47592
rect 469220 47540 469272 47592
rect 473268 47540 473320 47592
rect 550640 47540 550692 47592
rect 371240 46903 371292 46912
rect 371240 46869 371249 46903
rect 371249 46869 371283 46903
rect 371283 46869 371292 46903
rect 371240 46860 371292 46869
rect 129648 46180 129700 46232
rect 175280 46180 175332 46232
rect 197268 46180 197320 46232
rect 248420 46180 248472 46232
rect 269028 46180 269080 46232
rect 327080 46180 327132 46232
rect 329104 46180 329156 46232
rect 390560 46180 390612 46232
rect 429108 46180 429160 46232
rect 502432 46180 502484 46232
rect 235908 45568 235960 45620
rect 169668 44820 169720 44872
rect 218152 44820 218204 44872
rect 262036 44820 262088 44872
rect 318800 44820 318852 44872
rect 324228 44820 324280 44872
rect 387800 44820 387852 44872
rect 422208 44820 422260 44872
rect 494060 44820 494112 44872
rect 126888 43392 126940 43444
rect 171140 43392 171192 43444
rect 194508 43392 194560 43444
rect 244280 43392 244332 43444
rect 245476 43392 245528 43444
rect 302240 43392 302292 43444
rect 304908 43392 304960 43444
rect 365720 43392 365772 43444
rect 415308 43392 415360 43444
rect 487160 43392 487212 43444
rect 488356 43392 488408 43444
rect 565820 43392 565872 43444
rect 122656 42100 122708 42152
rect 167000 42100 167052 42152
rect 348976 42100 349028 42152
rect 414020 42100 414072 42152
rect 165528 42032 165580 42084
rect 213920 42032 213972 42084
rect 229008 42032 229060 42084
rect 282920 42032 282972 42084
rect 295248 42032 295300 42084
rect 356152 42032 356204 42084
rect 412548 42032 412600 42084
rect 484400 42032 484452 42084
rect 493968 42032 494020 42084
rect 572720 42032 572772 42084
rect 235816 41420 235868 41472
rect 504456 41352 504508 41404
rect 580172 41352 580224 41404
rect 345664 40740 345716 40792
rect 408592 40740 408644 40792
rect 119988 40672 120040 40724
rect 164240 40672 164292 40724
rect 173716 40672 173768 40724
rect 223580 40672 223632 40724
rect 230388 40672 230440 40724
rect 284300 40672 284352 40724
rect 285588 40672 285640 40724
rect 345020 40672 345072 40724
rect 408408 40672 408460 40724
rect 478880 40672 478932 40724
rect 115848 39312 115900 39364
rect 158720 39312 158772 39364
rect 162768 39312 162820 39364
rect 209780 39312 209832 39364
rect 215208 39312 215260 39364
rect 269120 39312 269172 39364
rect 291108 39312 291160 39364
rect 350540 39312 350592 39364
rect 365628 39312 365680 39364
rect 433432 39312 433484 39364
rect 438768 39312 438820 39364
rect 512000 39312 512052 39364
rect 353300 38564 353352 38616
rect 353392 38564 353444 38616
rect 378140 38607 378192 38616
rect 378140 38573 378149 38607
rect 378149 38573 378183 38607
rect 378183 38573 378192 38607
rect 378140 38564 378192 38573
rect 495440 38607 495492 38616
rect 495440 38573 495449 38607
rect 495449 38573 495483 38607
rect 495483 38573 495492 38607
rect 495440 38564 495492 38573
rect 108948 37884 109000 37936
rect 151820 37884 151872 37936
rect 158628 37884 158680 37936
rect 205640 37884 205692 37936
rect 206928 37884 206980 37936
rect 259460 37884 259512 37936
rect 262128 37884 262180 37936
rect 320180 37884 320232 37936
rect 331128 37884 331180 37936
rect 394700 37884 394752 37936
rect 405648 37884 405700 37936
rect 476120 37884 476172 37936
rect 477408 37884 477460 37936
rect 554872 37884 554924 37936
rect 371240 37315 371292 37324
rect 371240 37281 371249 37315
rect 371249 37281 371283 37315
rect 371283 37281 371292 37315
rect 371240 37272 371292 37281
rect 154488 36592 154540 36644
rect 201500 36592 201552 36644
rect 106188 36524 106240 36576
rect 149060 36524 149112 36576
rect 198648 36524 198700 36576
rect 249800 36524 249852 36576
rect 251088 36524 251140 36576
rect 307760 36524 307812 36576
rect 311808 36524 311860 36576
rect 374092 36524 374144 36576
rect 401508 36524 401560 36576
rect 471980 36524 472032 36576
rect 484308 36524 484360 36576
rect 563152 36524 563204 36576
rect 3424 35844 3476 35896
rect 14464 35844 14516 35896
rect 410892 35887 410944 35896
rect 410892 35853 410901 35887
rect 410901 35853 410935 35887
rect 410935 35853 410944 35887
rect 410892 35844 410944 35853
rect 102048 35164 102100 35216
rect 144920 35164 144972 35216
rect 151728 35164 151780 35216
rect 198740 35164 198792 35216
rect 199936 35164 199988 35216
rect 252652 35164 252704 35216
rect 259368 35164 259420 35216
rect 316040 35164 316092 35216
rect 321468 35164 321520 35216
rect 383660 35164 383712 35216
rect 398748 35164 398800 35216
rect 467932 35164 467984 35216
rect 481548 35164 481600 35216
rect 558920 35164 558972 35216
rect 144828 33804 144880 33856
rect 191840 33804 191892 33856
rect 99288 33736 99340 33788
rect 140780 33736 140832 33788
rect 190368 33736 190420 33788
rect 241520 33736 241572 33788
rect 277308 33736 277360 33788
rect 336740 33736 336792 33788
rect 337384 33736 337436 33788
rect 389180 33736 389232 33788
rect 395988 33736 396040 33788
rect 465080 33736 465132 33788
rect 474648 33736 474700 33788
rect 552020 33736 552072 33788
rect 142068 32444 142120 32496
rect 187700 32444 187752 32496
rect 249708 32444 249760 32496
rect 305000 32444 305052 32496
rect 96436 32376 96488 32428
rect 138020 32376 138072 32428
rect 187608 32376 187660 32428
rect 237380 32376 237432 32428
rect 302148 32376 302200 32428
rect 362960 32376 363012 32428
rect 391848 32376 391900 32428
rect 460940 32376 460992 32428
rect 471796 32376 471848 32428
rect 547880 32376 547932 32428
rect 137928 31016 137980 31068
rect 183560 31016 183612 31068
rect 185584 31016 185636 31068
rect 234620 31016 234672 31068
rect 240048 31016 240100 31068
rect 295340 31016 295392 31068
rect 313188 31016 313240 31068
rect 375380 31016 375432 31068
rect 389088 31016 389140 31068
rect 458180 31016 458232 31068
rect 464988 31016 465040 31068
rect 540980 31016 541032 31068
rect 504364 30268 504416 30320
rect 580172 30268 580224 30320
rect 135168 29656 135220 29708
rect 180800 29656 180852 29708
rect 92296 29588 92348 29640
rect 133880 29588 133932 29640
rect 180708 29588 180760 29640
rect 230480 29588 230532 29640
rect 291200 29588 291252 29640
rect 310428 29588 310480 29640
rect 372620 29588 372672 29640
rect 380164 29588 380216 29640
rect 447140 29588 447192 29640
rect 378140 29087 378192 29096
rect 378140 29053 378149 29087
rect 378149 29053 378183 29087
rect 378183 29053 378192 29087
rect 378140 29044 378192 29053
rect 495440 29019 495492 29028
rect 495440 28985 495449 29019
rect 495449 28985 495483 29019
rect 495483 28985 495492 29019
rect 495440 28976 495492 28985
rect 378140 28908 378192 28960
rect 378232 28908 378284 28960
rect 89628 28228 89680 28280
rect 131120 28228 131172 28280
rect 132408 28228 132460 28280
rect 176660 28228 176712 28280
rect 177948 28228 178000 28280
rect 227812 28228 227864 28280
rect 233148 28228 233200 28280
rect 287152 28228 287204 28280
rect 288348 28228 288400 28280
rect 347780 28228 347832 28280
rect 375288 28228 375340 28280
rect 443092 28228 443144 28280
rect 448428 28228 448480 28280
rect 523040 28228 523092 28280
rect 353300 27548 353352 27600
rect 353852 27548 353904 27600
rect 371240 27591 371292 27600
rect 371240 27557 371249 27591
rect 371249 27557 371283 27591
rect 371283 27557 371292 27591
rect 371240 27548 371292 27557
rect 128268 26936 128320 26988
rect 173900 26936 173952 26988
rect 171048 26868 171100 26920
rect 219440 26868 219492 26920
rect 223488 26868 223540 26920
rect 277400 26868 277452 26920
rect 278688 26868 278740 26920
rect 338120 26868 338172 26920
rect 372528 26868 372580 26920
rect 440240 26868 440292 26920
rect 445668 26868 445720 26920
rect 520372 26868 520424 26920
rect 410984 26256 411036 26308
rect 125508 25576 125560 25628
rect 169760 25576 169812 25628
rect 216588 25576 216640 25628
rect 270592 25576 270644 25628
rect 168288 25508 168340 25560
rect 216680 25508 216732 25560
rect 266176 25508 266228 25560
rect 322940 25508 322992 25560
rect 362868 25508 362920 25560
rect 429200 25508 429252 25560
rect 482836 25508 482888 25560
rect 561680 25508 561732 25560
rect 202788 24148 202840 24200
rect 253940 24148 253992 24200
rect 122748 24080 122800 24132
rect 167092 24080 167144 24132
rect 252468 24080 252520 24132
rect 309140 24080 309192 24132
rect 349068 24080 349120 24132
rect 415400 24080 415452 24132
rect 470508 24080 470560 24132
rect 546592 24080 546644 24132
rect 161388 22788 161440 22840
rect 209872 22788 209924 22840
rect 118608 22720 118660 22772
rect 162860 22720 162912 22772
rect 204168 22720 204220 22772
rect 255320 22720 255372 22772
rect 256608 22720 256660 22772
rect 313372 22720 313424 22772
rect 333888 22720 333940 22772
rect 397552 22720 397604 22772
rect 453948 22720 454000 22772
rect 528652 22720 528704 22772
rect 410984 22108 411036 22160
rect 3148 22040 3200 22092
rect 79416 22040 79468 22092
rect 226248 21428 226300 21480
rect 278872 21428 278924 21480
rect 322848 21428 322900 21480
rect 386420 21428 386472 21480
rect 114468 21360 114520 21412
rect 158812 21360 158864 21412
rect 166908 21360 166960 21412
rect 215300 21360 215352 21412
rect 266268 21360 266320 21412
rect 324320 21360 324372 21412
rect 384856 21360 384908 21412
rect 454040 21360 454092 21412
rect 467748 21360 467800 21412
rect 543740 21360 543792 21412
rect 111708 19932 111760 19984
rect 154580 19932 154632 19984
rect 157248 19932 157300 19984
rect 204260 19932 204312 19984
rect 205548 19932 205600 19984
rect 258080 19932 258132 19984
rect 293868 19932 293920 19984
rect 354680 19932 354732 19984
rect 355968 19932 356020 19984
rect 422300 19932 422352 19984
rect 463608 19932 463660 19984
rect 539600 19932 539652 19984
rect 369860 19295 369912 19304
rect 369860 19261 369869 19295
rect 369869 19261 369903 19295
rect 369903 19261 369912 19295
rect 369860 19252 369912 19261
rect 378140 19295 378192 19304
rect 378140 19261 378149 19295
rect 378149 19261 378183 19295
rect 378183 19261 378192 19295
rect 378140 19252 378192 19261
rect 389180 19252 389232 19304
rect 389364 19252 389416 19304
rect 397460 19295 397512 19304
rect 397460 19261 397469 19295
rect 397469 19261 397503 19295
rect 397503 19261 397512 19295
rect 397460 19252 397512 19261
rect 408592 19252 408644 19304
rect 409696 19252 409748 19304
rect 414020 19252 414072 19304
rect 414480 19252 414532 19304
rect 415400 19295 415452 19304
rect 415400 19261 415409 19295
rect 415409 19261 415443 19295
rect 415443 19261 415452 19295
rect 415400 19252 415452 19261
rect 495440 19252 495492 19304
rect 495624 19252 495676 19304
rect 561680 19295 561732 19304
rect 561680 19261 561689 19295
rect 561689 19261 561723 19295
rect 561723 19261 561732 19295
rect 561680 19252 561732 19261
rect 113824 18572 113876 18624
rect 150532 18572 150584 18624
rect 153844 18572 153896 18624
rect 201592 18572 201644 18624
rect 222108 18572 222160 18624
rect 276020 18572 276072 18624
rect 284208 18572 284260 18624
rect 343640 18572 343692 18624
rect 346308 18572 346360 18624
rect 411904 18572 411956 18624
rect 455420 18572 455472 18624
rect 456708 18572 456760 18624
rect 532700 18572 532752 18624
rect 412088 18504 412140 18556
rect 371240 18003 371292 18012
rect 371240 17969 371249 18003
rect 371249 17969 371283 18003
rect 371283 17969 371292 18003
rect 371240 17960 371292 17969
rect 571984 17892 572036 17944
rect 579804 17892 579856 17944
rect 281448 17280 281500 17332
rect 339592 17280 339644 17332
rect 104808 17212 104860 17264
rect 147680 17212 147732 17264
rect 150348 17212 150400 17264
rect 197360 17212 197412 17264
rect 209688 17212 209740 17264
rect 262312 17212 262364 17264
rect 339408 17212 339460 17264
rect 404360 17212 404412 17264
rect 451188 17212 451240 17264
rect 525800 17212 525852 17264
rect 102784 15852 102836 15904
rect 143540 15852 143592 15904
rect 147588 15852 147640 15904
rect 193312 15852 193364 15904
rect 195888 15852 195940 15904
rect 247040 15852 247092 15904
rect 267648 15852 267700 15904
rect 325700 15852 325752 15904
rect 326988 15852 327040 15904
rect 390652 15852 390704 15904
rect 437388 15852 437440 15904
rect 512092 15852 512144 15904
rect 320088 14492 320140 14544
rect 382372 14492 382424 14544
rect 97908 14424 97960 14476
rect 140872 14424 140924 14476
rect 143448 14424 143500 14476
rect 190460 14424 190512 14476
rect 193128 14424 193180 14476
rect 244372 14424 244424 14476
rect 257988 14424 258040 14476
rect 314660 14424 314712 14476
rect 382188 14424 382240 14476
rect 451372 14424 451424 14476
rect 460848 14424 460900 14476
rect 536932 14424 536984 14476
rect 97264 13064 97316 13116
rect 126980 13064 127032 13116
rect 140688 13064 140740 13116
rect 186320 13064 186372 13116
rect 189724 13064 189776 13116
rect 240140 13064 240192 13116
rect 255228 13064 255280 13116
rect 311900 13064 311952 13116
rect 317328 13064 317380 13116
rect 379520 13064 379572 13116
rect 434628 13064 434680 13116
rect 507860 13064 507912 13116
rect 354680 12452 354732 12504
rect 371240 12452 371292 12504
rect 372620 12452 372672 12504
rect 394700 12452 394752 12504
rect 350540 12384 350592 12436
rect 351368 12384 351420 12436
rect 351920 12384 351972 12436
rect 352564 12384 352616 12436
rect 358820 12384 358872 12436
rect 359740 12384 359792 12436
rect 354956 12316 355008 12368
rect 371608 12316 371660 12368
rect 375380 12384 375432 12436
rect 376392 12384 376444 12436
rect 376760 12384 376812 12436
rect 377588 12384 377640 12436
rect 391940 12384 391992 12436
rect 393044 12384 393096 12436
rect 393412 12384 393464 12436
rect 394240 12384 394292 12436
rect 372804 12316 372856 12368
rect 396080 12384 396132 12436
rect 396632 12384 396684 12436
rect 412640 12384 412692 12436
rect 413284 12384 413336 12436
rect 554872 12384 554924 12436
rect 555976 12384 556028 12436
rect 557540 12384 557592 12436
rect 558368 12384 558420 12436
rect 558920 12384 558972 12436
rect 559564 12384 559616 12436
rect 395436 12316 395488 12368
rect 427728 11772 427780 11824
rect 501236 11772 501288 11824
rect 92388 11704 92440 11756
rect 132592 11704 132644 11756
rect 133788 11704 133840 11756
rect 179420 11704 179472 11756
rect 183468 11704 183520 11756
rect 233240 11704 233292 11756
rect 241428 11704 241480 11756
rect 296812 11704 296864 11756
rect 300768 11704 300820 11756
rect 361580 11704 361632 11756
rect 362224 11704 362276 11756
rect 419540 11704 419592 11756
rect 500868 11704 500920 11756
rect 581092 11704 581144 11756
rect 309784 10344 309836 10396
rect 368480 10344 368532 10396
rect 95148 10276 95200 10328
rect 136640 10276 136692 10328
rect 138664 10276 138716 10328
rect 183652 10276 183704 10328
rect 186228 10276 186280 10328
rect 236092 10276 236144 10328
rect 248328 10276 248380 10328
rect 305092 10276 305144 10328
rect 344928 10276 344980 10328
rect 410800 10276 410852 10328
rect 424968 10276 425020 10328
rect 497740 10276 497792 10328
rect 499488 10276 499540 10328
rect 579620 10276 579672 10328
rect 370412 9664 370464 9716
rect 378784 9664 378836 9716
rect 397828 9664 397880 9716
rect 415676 9664 415728 9716
rect 561956 9664 562008 9716
rect 353760 9596 353812 9648
rect 354956 9596 355008 9648
rect 389456 9596 389508 9648
rect 395436 9596 395488 9648
rect 495440 9596 495492 9648
rect 353760 9460 353812 9512
rect 354956 9460 355008 9512
rect 389456 9460 389508 9512
rect 395436 9460 395488 9512
rect 88248 8916 88300 8968
rect 130200 8916 130252 8968
rect 131028 8916 131080 8968
rect 176568 8916 176620 8968
rect 179328 8916 179380 8968
rect 230112 8916 230164 8968
rect 245568 8916 245620 8968
rect 301412 8916 301464 8968
rect 303528 8916 303580 8968
rect 365812 8916 365864 8968
rect 369768 8916 369820 8968
rect 437020 8916 437072 8968
rect 438124 8916 438176 8968
rect 486976 8916 487028 8968
rect 487068 8916 487120 8968
rect 565544 8916 565596 8968
rect 410892 8415 410944 8424
rect 410892 8381 410901 8415
rect 410901 8381 410935 8415
rect 410935 8381 410944 8415
rect 410892 8372 410944 8381
rect 3424 8236 3476 8288
rect 79324 8236 79376 8288
rect 410892 8279 410944 8288
rect 410892 8245 410901 8279
rect 410901 8245 410935 8279
rect 410935 8245 410944 8279
rect 410892 8236 410944 8245
rect 86868 7624 86920 7676
rect 128912 7624 128964 7676
rect 358728 7624 358780 7676
rect 426348 7624 426400 7676
rect 124128 7556 124180 7608
rect 169392 7556 169444 7608
rect 176384 7556 176436 7608
rect 226524 7556 226576 7608
rect 238668 7556 238720 7608
rect 294328 7556 294380 7608
rect 298008 7556 298060 7608
rect 356060 7556 356112 7608
rect 357348 7556 357400 7608
rect 374000 7556 374052 7608
rect 375196 7556 375248 7608
rect 390560 7556 390612 7608
rect 391848 7556 391900 7608
rect 416780 7556 416832 7608
rect 417976 7556 418028 7608
rect 420828 7556 420880 7608
rect 494152 7556 494204 7608
rect 496728 7556 496780 7608
rect 576216 7556 576268 7608
rect 358544 7488 358596 7540
rect 121368 6196 121420 6248
rect 165896 6196 165948 6248
rect 160008 6128 160060 6180
rect 208676 6128 208728 6180
rect 219348 6128 219400 6180
rect 272892 6128 272944 6180
rect 274548 6128 274600 6180
rect 333612 6128 333664 6180
rect 336648 6128 336700 6180
rect 401324 6128 401376 6180
rect 483480 6128 483532 6180
rect 489828 6128 489880 6180
rect 569040 6128 569092 6180
rect 502984 5448 503036 5500
rect 504824 5448 504876 5500
rect 231124 4836 231176 4888
rect 265808 4836 265860 4888
rect 353208 4836 353260 4888
rect 85488 4768 85540 4820
rect 126612 4768 126664 4820
rect 129004 4768 129056 4820
rect 172980 4768 173032 4820
rect 173808 4768 173860 4820
rect 222936 4768 222988 4820
rect 264888 4768 264940 4820
rect 322848 4768 322900 4820
rect 323584 4768 323636 4820
rect 347872 4768 347924 4820
rect 419172 4836 419224 4888
rect 418068 4768 418120 4820
rect 490564 4768 490616 4820
rect 560944 4768 560996 4820
rect 572628 4768 572680 4820
rect 520280 4156 520332 4208
rect 521476 4156 521528 4208
rect 528652 4156 528704 4208
rect 529848 4156 529900 4208
rect 384948 4088 385000 4140
rect 453672 4088 453724 4140
rect 471888 4088 471940 4140
rect 550088 4088 550140 4140
rect 378048 4020 378100 4072
rect 446588 4020 446640 4072
rect 476028 4020 476080 4072
rect 553584 4020 553636 4072
rect 91008 3952 91060 4004
rect 132500 3952 132552 4004
rect 394608 3952 394660 4004
rect 464436 3952 464488 4004
rect 478788 3952 478840 4004
rect 557172 3952 557224 4004
rect 574744 3952 574796 4004
rect 577412 3952 577464 4004
rect 93768 3884 93820 3936
rect 136088 3884 136140 3936
rect 390468 3884 390520 3936
rect 460848 3884 460900 3936
rect 482928 3884 482980 3936
rect 560760 3884 560812 3936
rect 100668 3816 100720 3868
rect 143264 3816 143316 3868
rect 387708 3816 387760 3868
rect 457260 3816 457312 3868
rect 485688 3816 485740 3868
rect 564348 3816 564400 3868
rect 96528 3748 96580 3800
rect 139676 3748 139728 3800
rect 380808 3748 380860 3800
rect 450176 3748 450228 3800
rect 469128 3748 469180 3800
rect 546500 3748 546552 3800
rect 103428 3680 103480 3732
rect 146852 3680 146904 3732
rect 397368 3680 397420 3732
rect 467840 3680 467892 3732
rect 492588 3680 492640 3732
rect 107568 3612 107620 3664
rect 150440 3612 150492 3664
rect 404268 3612 404320 3664
rect 475108 3612 475160 3664
rect 488448 3612 488500 3664
rect 110328 3544 110380 3596
rect 153936 3544 153988 3596
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 218152 3544 218204 3596
rect 219348 3544 219400 3596
rect 227720 3544 227772 3596
rect 228916 3544 228968 3596
rect 262220 3544 262272 3596
rect 263416 3544 263468 3596
rect 270500 3544 270552 3596
rect 271696 3544 271748 3596
rect 278872 3544 278924 3596
rect 280068 3544 280120 3596
rect 331220 3544 331272 3596
rect 332416 3544 332468 3596
rect 365720 3544 365772 3596
rect 366916 3544 366968 3596
rect 382372 3544 382424 3596
rect 383568 3544 383620 3596
rect 400128 3544 400180 3596
rect 471520 3544 471572 3596
rect 495256 3544 495308 3596
rect 502248 3680 502300 3732
rect 582196 3680 582248 3732
rect 567200 3612 567252 3664
rect 572 3476 624 3528
rect 81440 3476 81492 3528
rect 117228 3476 117280 3528
rect 1676 3408 1728 3460
rect 82820 3408 82872 3460
rect 113088 3408 113140 3460
rect 157524 3408 157576 3460
rect 158720 3476 158772 3528
rect 159916 3476 159968 3528
rect 167000 3476 167052 3528
rect 168196 3476 168248 3528
rect 183560 3476 183612 3528
rect 184848 3476 184900 3528
rect 209780 3476 209832 3528
rect 211068 3476 211120 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 252560 3476 252612 3528
rect 253848 3476 253900 3528
rect 287152 3476 287204 3528
rect 288348 3476 288400 3528
rect 305000 3476 305052 3528
rect 306196 3476 306248 3528
rect 313280 3476 313332 3528
rect 314568 3476 314620 3528
rect 347780 3476 347832 3528
rect 349068 3476 349120 3528
rect 411168 3476 411220 3528
rect 482284 3476 482336 3528
rect 494060 3476 494112 3528
rect 495348 3476 495400 3528
rect 571432 3544 571484 3596
rect 575020 3476 575072 3528
rect 161112 3408 161164 3460
rect 407028 3408 407080 3460
rect 478696 3408 478748 3460
rect 498108 3408 498160 3460
rect 578608 3408 578660 3460
rect 132592 3340 132644 3392
rect 133788 3340 133840 3392
rect 433340 3340 433392 3392
rect 434628 3340 434680 3392
rect 451280 3340 451332 3392
rect 452476 3340 452528 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 512000 3340 512052 3392
rect 513196 3340 513248 3392
rect 536840 3340 536892 3392
rect 538128 3340 538180 3392
rect 567200 3340 567252 3392
rect 567844 3340 567896 3392
rect 140780 3000 140832 3052
rect 142068 3000 142120 3052
rect 498200 2796 498252 2848
rect 499580 2796 499632 2848
rect 498936 2728 498988 2780
rect 500132 2728 500184 2780
rect 502340 2048 502392 2100
rect 503628 2048 503680 2100
rect 126980 552 127032 604
rect 127808 552 127860 604
rect 131120 552 131172 604
rect 131396 552 131448 604
rect 496544 595 496596 604
rect 496544 561 496553 595
rect 496553 561 496587 595
rect 496587 561 496596 595
rect 496544 552 496596 561
rect 579620 552 579672 604
rect 579804 552 579856 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3790 682272 3846 682281
rect 3790 682207 3846 682216
rect 3804 681766 3832 682207
rect 3792 681760 3844 681766
rect 3792 681702 3844 681708
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3238 624880 3294 624889
rect 3238 624815 3294 624824
rect 3252 623830 3280 624815
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 3436 585138 3464 667927
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 10324 652792 10376 652798
rect 10324 652734 10376 652740
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 8944 623824 8996 623830
rect 8944 623766 8996 623772
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 3514 610464 3570 610473
rect 3514 610399 3570 610408
rect 3424 585132 3476 585138
rect 3424 585074 3476 585080
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 513330 3464 553007
rect 3528 549234 3556 610399
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 603770 8064 605798
rect 8024 603764 8076 603770
rect 8024 603706 8076 603712
rect 8956 560250 8984 623766
rect 10336 572694 10364 652734
rect 24780 603838 24808 699654
rect 32404 681760 32456 681766
rect 32404 681702 32456 681708
rect 24768 603832 24820 603838
rect 24768 603774 24820 603780
rect 32416 596154 32444 681702
rect 41340 603906 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 73068 627972 73120 627978
rect 73068 627914 73120 627920
rect 73080 603974 73108 627914
rect 89640 604042 89668 699654
rect 89628 604036 89680 604042
rect 89628 603978 89680 603984
rect 73068 603968 73120 603974
rect 73068 603910 73120 603916
rect 41328 603900 41380 603906
rect 41328 603842 41380 603848
rect 105268 603832 105320 603838
rect 105268 603774 105320 603780
rect 89720 603764 89772 603770
rect 89720 603706 89772 603712
rect 89732 601868 89760 603706
rect 105280 601868 105308 603774
rect 106200 603770 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 136364 603968 136416 603974
rect 136364 603910 136416 603916
rect 120816 603900 120868 603906
rect 120816 603842 120868 603848
rect 106188 603764 106240 603770
rect 106188 603706 106240 603712
rect 120828 601868 120856 603842
rect 136376 601868 136404 603910
rect 137756 603838 137784 605798
rect 151912 604036 151964 604042
rect 151912 603978 151964 603984
rect 137744 603832 137796 603838
rect 137744 603774 137796 603780
rect 151924 601868 151952 603978
rect 154316 603906 154344 605798
rect 154304 603900 154356 603906
rect 154304 603842 154356 603848
rect 171060 603770 171088 700198
rect 198556 603900 198608 603906
rect 198556 603842 198608 603848
rect 183008 603832 183060 603838
rect 183008 603774 183060 603780
rect 167460 603764 167512 603770
rect 167460 603706 167512 603712
rect 171048 603764 171100 603770
rect 171048 603706 171100 603712
rect 167472 601868 167500 603706
rect 183020 601868 183048 603774
rect 198568 601868 198596 603842
rect 202800 603838 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219348 627972 219400 627978
rect 219348 627914 219400 627920
rect 202788 603832 202840 603838
rect 202788 603774 202840 603780
rect 219360 603770 219388 627914
rect 235920 603838 235948 699654
rect 229652 603832 229704 603838
rect 229652 603774 229704 603780
rect 235908 603832 235960 603838
rect 235908 603774 235960 603780
rect 260748 603832 260800 603838
rect 260748 603774 260800 603780
rect 214104 603764 214156 603770
rect 214104 603706 214156 603712
rect 219348 603764 219400 603770
rect 219348 603706 219400 603712
rect 214116 601868 214144 603706
rect 229664 601868 229692 603774
rect 245200 603764 245252 603770
rect 245200 603706 245252 603712
rect 245212 601868 245240 603706
rect 260760 601868 260788 603774
rect 267660 603770 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654158 284064 663734
rect 284024 654152 284076 654158
rect 284024 654094 284076 654100
rect 284208 654152 284260 654158
rect 284208 654094 284260 654100
rect 284220 644450 284248 654094
rect 284036 644422 284248 644450
rect 284036 634846 284064 644422
rect 284024 634840 284076 634846
rect 284024 634782 284076 634788
rect 284208 634840 284260 634846
rect 284208 634782 284260 634788
rect 284220 625138 284248 634782
rect 284036 625110 284248 625138
rect 284036 615534 284064 625110
rect 284024 615528 284076 615534
rect 284024 615470 284076 615476
rect 284208 615528 284260 615534
rect 284208 615470 284260 615476
rect 284220 605826 284248 615470
rect 284036 605798 284248 605826
rect 284036 603770 284064 605798
rect 300780 604450 300808 699654
rect 332520 697610 332548 703520
rect 348804 703474 348832 703520
rect 364996 703474 365024 703520
rect 348804 703446 348924 703474
rect 364996 703446 365116 703474
rect 331220 697604 331272 697610
rect 331220 697546 331272 697552
rect 332508 697604 332560 697610
rect 332508 697546 332560 697552
rect 300768 604444 300820 604450
rect 300768 604386 300820 604392
rect 307484 604444 307536 604450
rect 307484 604386 307536 604392
rect 267648 603764 267700 603770
rect 267648 603706 267700 603712
rect 276296 603764 276348 603770
rect 276296 603706 276348 603712
rect 284024 603764 284076 603770
rect 284024 603706 284076 603712
rect 291844 603764 291896 603770
rect 291844 603706 291896 603712
rect 276308 601868 276336 603706
rect 291856 601868 291884 603706
rect 307496 601868 307524 604386
rect 331232 603770 331260 697546
rect 348896 692850 348924 703446
rect 365088 692850 365116 703446
rect 347780 692844 347832 692850
rect 347780 692786 347832 692792
rect 348884 692844 348936 692850
rect 348884 692786 348936 692792
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 347792 683074 347820 692786
rect 364352 683074 364380 692786
rect 347792 683046 348004 683074
rect 364352 683046 364564 683074
rect 347976 673538 348004 683046
rect 364536 673538 364564 683046
rect 347780 673532 347832 673538
rect 347780 673474 347832 673480
rect 347964 673532 348016 673538
rect 347964 673474 348016 673480
rect 364340 673532 364392 673538
rect 364340 673474 364392 673480
rect 364524 673532 364576 673538
rect 364524 673474 364576 673480
rect 347792 663762 347820 673474
rect 364352 663762 364380 673474
rect 347792 663734 348004 663762
rect 364352 663734 364564 663762
rect 347976 654158 348004 663734
rect 364536 654158 364564 663734
rect 347780 654152 347832 654158
rect 347780 654094 347832 654100
rect 347964 654152 348016 654158
rect 347964 654094 348016 654100
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 347792 644450 347820 654094
rect 364352 644450 364380 654094
rect 347792 644422 348004 644450
rect 364352 644422 364564 644450
rect 347976 634846 348004 644422
rect 364536 634846 364564 644422
rect 347780 634840 347832 634846
rect 347780 634782 347832 634788
rect 347964 634840 348016 634846
rect 347964 634782 348016 634788
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 347792 625138 347820 634782
rect 364352 625138 364380 634782
rect 347792 625110 348004 625138
rect 364352 625110 364564 625138
rect 347976 615534 348004 625110
rect 364536 615534 364564 625110
rect 347780 615528 347832 615534
rect 347780 615470 347832 615476
rect 347964 615528 348016 615534
rect 347964 615470 348016 615476
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 347792 605826 347820 615470
rect 364352 605826 364380 615470
rect 347792 605798 348004 605826
rect 364352 605798 364564 605826
rect 347976 603770 348004 605798
rect 364536 603770 364564 605798
rect 385224 603900 385276 603906
rect 385224 603842 385276 603848
rect 323032 603764 323084 603770
rect 323032 603706 323084 603712
rect 331220 603764 331272 603770
rect 331220 603706 331272 603712
rect 338580 603764 338632 603770
rect 338580 603706 338632 603712
rect 347964 603764 348016 603770
rect 347964 603706 348016 603712
rect 354128 603764 354180 603770
rect 354128 603706 354180 603712
rect 364524 603764 364576 603770
rect 364524 603706 364576 603712
rect 369676 603764 369728 603770
rect 369676 603706 369728 603712
rect 323044 601868 323072 603706
rect 338592 601868 338620 603706
rect 354140 601868 354168 603706
rect 369688 601868 369716 603706
rect 385236 601868 385264 603842
rect 397472 603770 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 413756 698290 413784 703446
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 429856 684486 429884 703520
rect 429200 684480 429252 684486
rect 429200 684422 429252 684428
rect 429844 684480 429896 684486
rect 429844 684422 429896 684428
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 429212 683126 429240 684422
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 429200 683120 429252 683126
rect 429200 683062 429252 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 413112 659682 413140 666538
rect 429672 659682 429700 666538
rect 412928 659654 413140 659682
rect 429488 659654 429700 659682
rect 412928 647290 412956 659654
rect 429488 647290 429516 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 412836 640422 412864 647226
rect 429396 640422 429424 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 412928 630698 412956 640358
rect 429488 630698 429516 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 412744 630578 412772 630634
rect 429304 630578 429332 630634
rect 412744 630550 412864 630578
rect 429304 630550 429424 630578
rect 412836 621058 412864 630550
rect 429396 621058 429424 630550
rect 412836 621030 412956 621058
rect 429396 621030 429516 621058
rect 412928 611386 412956 621030
rect 429488 611386 429516 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 412744 603906 412772 611322
rect 412732 603900 412784 603906
rect 412732 603842 412784 603848
rect 429304 603838 429332 611322
rect 447416 603900 447468 603906
rect 447416 603842 447468 603848
rect 400772 603832 400824 603838
rect 400772 603774 400824 603780
rect 429292 603832 429344 603838
rect 429292 603774 429344 603780
rect 431868 603832 431920 603838
rect 431868 603774 431920 603780
rect 397460 603764 397512 603770
rect 397460 603706 397512 603712
rect 400784 601868 400812 603774
rect 416320 603764 416372 603770
rect 416320 603706 416372 603712
rect 416332 601868 416360 603706
rect 431880 601868 431908 603774
rect 447428 601868 447456 603842
rect 462332 603770 462360 703520
rect 478524 703474 478552 703520
rect 494808 703474 494836 703520
rect 478524 703446 478644 703474
rect 494808 703446 494928 703474
rect 478616 692850 478644 703446
rect 494900 692850 494928 703446
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 477512 683074 477540 692786
rect 494072 683074 494100 692786
rect 477512 683046 477724 683074
rect 494072 683046 494284 683074
rect 477696 673538 477724 683046
rect 494256 673538 494284 683046
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 494060 673532 494112 673538
rect 494060 673474 494112 673480
rect 494244 673532 494296 673538
rect 494244 673474 494296 673480
rect 477512 663762 477540 673474
rect 494072 663762 494100 673474
rect 477512 663734 477724 663762
rect 494072 663734 494284 663762
rect 477696 654158 477724 663734
rect 494256 654158 494284 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 477512 644450 477540 654094
rect 494072 644450 494100 654094
rect 477512 644422 477724 644450
rect 494072 644422 494284 644450
rect 477696 634846 477724 644422
rect 494256 634846 494284 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 477512 625138 477540 634782
rect 494072 625138 494100 634782
rect 477512 625110 477724 625138
rect 494072 625110 494284 625138
rect 477696 615534 477724 625110
rect 494256 615534 494284 625110
rect 477500 615528 477552 615534
rect 477500 615470 477552 615476
rect 477684 615528 477736 615534
rect 477684 615470 477736 615476
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 477512 605826 477540 615470
rect 494072 605826 494100 615470
rect 477512 605798 477724 605826
rect 494072 605798 494284 605826
rect 477696 603838 477724 605798
rect 494256 603906 494284 605798
rect 494244 603900 494296 603906
rect 494244 603842 494296 603848
rect 494336 603900 494388 603906
rect 494336 603842 494388 603848
rect 477684 603832 477736 603838
rect 477684 603774 477736 603780
rect 478512 603832 478564 603838
rect 478512 603774 478564 603780
rect 462320 603764 462372 603770
rect 462320 603706 462372 603712
rect 462964 603764 463016 603770
rect 462964 603706 463016 603712
rect 462976 601868 463004 603706
rect 478524 601868 478552 603774
rect 494348 601882 494376 603842
rect 527192 603770 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 538864 696992 538916 696998
rect 538864 696934 538916 696940
rect 536104 673532 536156 673538
rect 536104 673474 536156 673480
rect 529204 650072 529256 650078
rect 529204 650014 529256 650020
rect 527180 603764 527232 603770
rect 527180 603706 527232 603712
rect 494086 601854 494376 601882
rect 505008 597508 505060 597514
rect 505008 597450 505060 597456
rect 505020 596329 505048 597450
rect 505006 596320 505062 596329
rect 505006 596255 505062 596264
rect 32404 596148 32456 596154
rect 32404 596090 32456 596096
rect 78680 596148 78732 596154
rect 78680 596090 78732 596096
rect 78692 595921 78720 596090
rect 78678 595912 78734 595921
rect 78678 595847 78734 595856
rect 13084 594856 13136 594862
rect 13084 594798 13136 594804
rect 10324 572688 10376 572694
rect 10324 572630 10376 572636
rect 10324 567248 10376 567254
rect 10324 567190 10376 567196
rect 8944 560244 8996 560250
rect 8944 560186 8996 560192
rect 3516 549228 3568 549234
rect 3516 549170 3568 549176
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3424 513324 3476 513330
rect 3424 513266 3476 513272
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 3436 489870 3464 509895
rect 3528 500954 3556 538591
rect 10336 525774 10364 567190
rect 13096 536790 13124 594798
rect 507124 592068 507176 592074
rect 507124 592010 507176 592016
rect 504640 586492 504692 586498
rect 504640 586434 504692 586440
rect 504652 585177 504680 586434
rect 504638 585168 504694 585177
rect 78680 585132 78732 585138
rect 504638 585103 504694 585112
rect 78680 585074 78732 585080
rect 78692 583953 78720 585074
rect 78678 583944 78734 583953
rect 78678 583879 78734 583888
rect 505008 574048 505060 574054
rect 505006 574016 505008 574025
rect 505060 574016 505062 574025
rect 505006 573951 505062 573960
rect 78680 572688 78732 572694
rect 78680 572630 78732 572636
rect 78692 572121 78720 572630
rect 78678 572112 78734 572121
rect 78678 572047 78734 572056
rect 505008 563032 505060 563038
rect 505006 563000 505008 563009
rect 505060 563000 505062 563009
rect 505006 562935 505062 562944
rect 78680 560244 78732 560250
rect 78680 560186 78732 560192
rect 78692 560153 78720 560186
rect 78678 560144 78734 560153
rect 78678 560079 78734 560088
rect 504364 556232 504416 556238
rect 504364 556174 504416 556180
rect 78680 549228 78732 549234
rect 78680 549170 78732 549176
rect 78692 548321 78720 549170
rect 78678 548312 78734 548321
rect 78678 548247 78734 548256
rect 13084 536784 13136 536790
rect 13084 536726 13136 536732
rect 78680 536784 78732 536790
rect 78680 536726 78732 536732
rect 78692 536353 78720 536726
rect 78678 536344 78734 536353
rect 78678 536279 78734 536288
rect 10324 525768 10376 525774
rect 10324 525710 10376 525716
rect 78680 525768 78732 525774
rect 78680 525710 78732 525716
rect 78692 524521 78720 525710
rect 78678 524512 78734 524521
rect 78678 524447 78734 524456
rect 504180 518560 504232 518566
rect 504178 518528 504180 518537
rect 504232 518528 504234 518537
rect 504178 518463 504234 518472
rect 78680 513324 78732 513330
rect 78680 513266 78732 513272
rect 78692 512553 78720 513266
rect 78678 512544 78734 512553
rect 78678 512479 78734 512488
rect 3516 500948 3568 500954
rect 3516 500890 3568 500896
rect 78680 500948 78732 500954
rect 78680 500890 78732 500896
rect 78692 500721 78720 500890
rect 78678 500712 78734 500721
rect 78678 500647 78734 500656
rect 504376 496369 504404 556174
rect 505008 552016 505060 552022
rect 505008 551958 505060 551964
rect 505020 551857 505048 551958
rect 505006 551848 505062 551857
rect 505006 551783 505062 551792
rect 505008 540932 505060 540938
rect 505008 540874 505060 540880
rect 505020 540705 505048 540874
rect 505006 540696 505062 540705
rect 505006 540631 505062 540640
rect 505744 532772 505796 532778
rect 505744 532714 505796 532720
rect 505008 529916 505060 529922
rect 505008 529858 505060 529864
rect 505020 529689 505048 529858
rect 505006 529680 505062 529689
rect 505006 529615 505062 529624
rect 505008 507748 505060 507754
rect 505008 507690 505060 507696
rect 505020 507385 505048 507690
rect 505006 507376 505062 507385
rect 505006 507311 505062 507320
rect 504362 496360 504418 496369
rect 504362 496295 504418 496304
rect 3514 495544 3570 495553
rect 3514 495479 3570 495488
rect 3424 489864 3476 489870
rect 3424 489806 3476 489812
rect 3422 481128 3478 481137
rect 3422 481063 3478 481072
rect 3436 465050 3464 481063
rect 3528 477494 3556 495479
rect 78680 489864 78732 489870
rect 78680 489806 78732 489812
rect 78692 488753 78720 489806
rect 78678 488744 78734 488753
rect 78678 488679 78734 488688
rect 504364 485852 504416 485858
rect 504364 485794 504416 485800
rect 3516 477488 3568 477494
rect 3516 477430 3568 477436
rect 78680 477488 78732 477494
rect 78680 477430 78732 477436
rect 78692 476921 78720 477430
rect 78678 476912 78734 476921
rect 78678 476847 78734 476856
rect 503720 474360 503772 474366
rect 503720 474302 503772 474308
rect 503732 474065 503760 474302
rect 503718 474056 503774 474065
rect 503718 473991 503774 474000
rect 3424 465044 3476 465050
rect 3424 464986 3476 464992
rect 78680 465044 78732 465050
rect 78680 464986 78732 464992
rect 78692 464953 78720 464986
rect 78678 464944 78734 464953
rect 78678 464879 78734 464888
rect 503812 463684 503864 463690
rect 503812 463626 503864 463632
rect 503824 463049 503852 463626
rect 503810 463040 503866 463049
rect 503810 462975 503866 462984
rect 78678 453112 78734 453121
rect 78678 453047 78734 453056
rect 78692 452606 78720 453047
rect 3424 452600 3476 452606
rect 3424 452542 3476 452548
rect 78680 452600 78732 452606
rect 78680 452542 78732 452548
rect 504180 452600 504232 452606
rect 504180 452542 504232 452548
rect 3436 452441 3464 452542
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 504192 451897 504220 452542
rect 504178 451888 504234 451897
rect 504178 451823 504234 451832
rect 78678 441144 78734 441153
rect 78678 441079 78734 441088
rect 78692 438870 78720 441079
rect 504376 440745 504404 485794
rect 505008 485784 505060 485790
rect 505008 485726 505060 485732
rect 505020 485217 505048 485726
rect 505006 485208 505062 485217
rect 505006 485143 505062 485152
rect 505756 474366 505784 532714
rect 507136 518566 507164 592010
rect 511264 579692 511316 579698
rect 511264 579634 511316 579640
rect 507124 518560 507176 518566
rect 507124 518502 507176 518508
rect 507124 509312 507176 509318
rect 507124 509254 507176 509260
rect 505744 474360 505796 474366
rect 505744 474302 505796 474308
rect 507136 463690 507164 509254
rect 511276 507754 511304 579634
rect 529216 563038 529244 650014
rect 536116 574054 536144 673474
rect 538876 597514 538904 696934
rect 542740 694142 542768 698226
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 692782 542584 694078
rect 542544 692776 542596 692782
rect 542544 692718 542596 692724
rect 542728 692776 542780 692782
rect 542728 692718 542780 692724
rect 542740 683233 542768 692718
rect 559668 684486 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 558920 684480 558972 684486
rect 558920 684422 558972 684428
rect 559656 684480 559708 684486
rect 559656 684422 559708 684428
rect 542358 683224 542414 683233
rect 542358 683159 542414 683168
rect 542726 683224 542782 683233
rect 542726 683159 542782 683168
rect 542372 683126 542400 683159
rect 558932 683126 558960 684422
rect 542360 683120 542412 683126
rect 542360 683062 542412 683068
rect 558920 683120 558972 683126
rect 558920 683062 558972 683068
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 542832 659682 542860 666538
rect 559392 659682 559420 666538
rect 542648 659654 542860 659682
rect 559208 659654 559420 659682
rect 542648 647290 542676 659654
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 542556 640422 542584 647226
rect 559116 640422 559144 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 542648 630698 542676 640358
rect 559208 630698 559236 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 542464 630578 542492 630634
rect 559024 630578 559052 630634
rect 542464 630550 542584 630578
rect 559024 630550 559144 630578
rect 542556 621058 542584 630550
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 571984 626612 572036 626618
rect 571984 626554 572036 626560
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 559116 621030 559236 621058
rect 542648 611386 542676 621030
rect 559208 611386 559236 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 542464 603838 542492 611322
rect 559024 603906 559052 611322
rect 559012 603900 559064 603906
rect 559012 603842 559064 603848
rect 542452 603832 542504 603838
rect 542452 603774 542504 603780
rect 565084 603152 565136 603158
rect 565084 603094 565136 603100
rect 538864 597508 538916 597514
rect 538864 597450 538916 597456
rect 536104 574048 536156 574054
rect 536104 573990 536156 573996
rect 529204 563032 529256 563038
rect 529204 562974 529256 562980
rect 565096 529922 565124 603094
rect 571996 540938 572024 626554
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 579894 592512 579950 592521
rect 579894 592447 579950 592456
rect 579908 592074 579936 592447
rect 579896 592068 579948 592074
rect 579896 592010 579948 592016
rect 580276 586498 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580264 586492 580316 586498
rect 580264 586434 580316 586440
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580368 552022 580396 639367
rect 580356 552016 580408 552022
rect 580356 551958 580408 551964
rect 580262 545592 580318 545601
rect 580262 545527 580318 545536
rect 571984 540932 572036 540938
rect 571984 540874 572036 540880
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 565084 529916 565136 529922
rect 565084 529858 565136 529864
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 511264 507748 511316 507754
rect 511264 507690 511316 507696
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580276 485790 580304 545527
rect 580354 498672 580410 498681
rect 580354 498607 580410 498616
rect 580264 485784 580316 485790
rect 580264 485726 580316 485732
rect 507124 463684 507176 463690
rect 507124 463626 507176 463632
rect 580262 463448 580318 463457
rect 580262 463383 580318 463392
rect 504362 440736 504418 440745
rect 504362 440671 504418 440680
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 504364 438932 504416 438938
rect 504364 438874 504416 438880
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 78680 438864 78732 438870
rect 78680 438806 78732 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 78678 429312 78734 429321
rect 78678 429247 78734 429256
rect 78692 425066 78720 429247
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 78680 425060 78732 425066
rect 78680 425002 78732 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 79322 417344 79378 417353
rect 79322 417279 79378 417288
rect 79336 396030 79364 417279
rect 504376 407425 504404 438874
rect 580276 430574 580304 463383
rect 580368 452606 580396 498607
rect 580356 452600 580408 452606
rect 580356 452542 580408 452548
rect 580446 451752 580502 451761
rect 580446 451687 580502 451696
rect 505008 430568 505060 430574
rect 505008 430510 505060 430516
rect 580264 430568 580316 430574
rect 580264 430510 580316 430516
rect 505020 429593 505048 430510
rect 505006 429584 505062 429593
rect 505006 429519 505062 429528
rect 580460 419490 580488 451687
rect 505008 419484 505060 419490
rect 505008 419426 505060 419432
rect 580448 419484 580500 419490
rect 580448 419426 580500 419432
rect 505020 418577 505048 419426
rect 505006 418568 505062 418577
rect 505006 418503 505062 418512
rect 580354 416528 580410 416537
rect 580354 416463 580410 416472
rect 504362 407416 504418 407425
rect 504362 407351 504418 407360
rect 79414 405512 79470 405521
rect 79414 405447 79470 405456
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 79324 396024 79376 396030
rect 79324 395966 79376 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 79322 393544 79378 393553
rect 79322 393479 79378 393488
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 79336 367062 79364 393479
rect 79428 380866 79456 405447
rect 580262 404832 580318 404841
rect 580262 404767 580318 404776
rect 505008 397452 505060 397458
rect 505008 397394 505060 397400
rect 505020 396273 505048 397394
rect 505006 396264 505062 396273
rect 505006 396199 505062 396208
rect 580276 386374 580304 404767
rect 580368 397458 580396 416463
rect 580356 397452 580408 397458
rect 580356 397394 580408 397400
rect 580354 393000 580410 393009
rect 580354 392935 580410 392944
rect 504548 386368 504600 386374
rect 504548 386310 504600 386316
rect 580264 386368 580316 386374
rect 580264 386310 580316 386316
rect 504560 385257 504588 386310
rect 504546 385248 504602 385257
rect 504546 385183 504602 385192
rect 79598 381712 79654 381721
rect 79598 381647 79654 381656
rect 79416 380860 79468 380866
rect 79416 380802 79468 380808
rect 79506 369744 79562 369753
rect 79506 369679 79562 369688
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 79324 367056 79376 367062
rect 79324 366998 79376 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 79414 357912 79470 357921
rect 79414 357847 79470 357856
rect 79322 345944 79378 345953
rect 79322 345879 79378 345888
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 79336 295322 79364 345879
rect 79428 309126 79456 357847
rect 79520 324290 79548 369679
rect 79612 338094 79640 381647
rect 580368 375358 580396 392935
rect 505008 375352 505060 375358
rect 505008 375294 505060 375300
rect 580356 375352 580408 375358
rect 580356 375294 580408 375300
rect 505020 374105 505048 375294
rect 505006 374096 505062 374105
rect 505006 374031 505062 374040
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 505006 362944 505062 362953
rect 580276 362914 580304 369543
rect 505006 362879 505008 362888
rect 505060 362879 505062 362888
rect 580264 362908 580316 362914
rect 505008 362850 505060 362856
rect 580264 362850 580316 362856
rect 580262 357912 580318 357921
rect 580262 357847 580318 357856
rect 580276 353258 580304 357847
rect 504640 353252 504692 353258
rect 504640 353194 504692 353200
rect 580264 353252 580316 353258
rect 580264 353194 580316 353200
rect 504652 351937 504680 353194
rect 504638 351928 504694 351937
rect 504638 351863 504694 351872
rect 580906 346080 580962 346089
rect 580906 346015 580962 346024
rect 580920 340882 580948 346015
rect 505008 340876 505060 340882
rect 505008 340818 505060 340824
rect 580908 340876 580960 340882
rect 580908 340818 580960 340824
rect 505020 340785 505048 340818
rect 505006 340776 505062 340785
rect 505006 340711 505062 340720
rect 79600 338088 79652 338094
rect 79600 338030 79652 338036
rect 79690 333976 79746 333985
rect 79690 333911 79746 333920
rect 79508 324284 79560 324290
rect 79508 324226 79560 324232
rect 79598 322144 79654 322153
rect 79598 322079 79654 322088
rect 79506 310176 79562 310185
rect 79506 310111 79562 310120
rect 79416 309120 79468 309126
rect 79416 309062 79468 309068
rect 79414 298344 79470 298353
rect 79414 298279 79470 298288
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 79324 295316 79376 295322
rect 79324 295258 79376 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 79322 286376 79378 286385
rect 79322 286311 79378 286320
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 78678 274544 78734 274553
rect 78678 274479 78734 274488
rect 78692 273290 78720 274479
rect 10324 273284 10376 273290
rect 10324 273226 10376 273232
rect 78680 273284 78732 273290
rect 78680 273226 78732 273232
rect 3148 266348 3200 266354
rect 3148 266290 3200 266296
rect 3160 265713 3188 266290
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 10336 208350 10364 273226
rect 25504 238808 25556 238814
rect 78680 238808 78732 238814
rect 25504 238750 25556 238756
rect 78678 238776 78680 238785
rect 78732 238776 78734 238785
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 10324 208344 10376 208350
rect 10324 208286 10376 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 24124 202904 24176 202910
rect 24124 202846 24176 202852
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 8944 167068 8996 167074
rect 8944 167010 8996 167016
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 8956 79490 8984 167010
rect 14464 131164 14516 131170
rect 14464 131106 14516 131112
rect 3516 79484 3568 79490
rect 3516 79426 3568 79432
rect 8944 79484 8996 79490
rect 8944 79426 8996 79432
rect 3528 78985 3556 79426
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 14476 35902 14504 131106
rect 24136 122806 24164 202846
rect 25516 165578 25544 238750
rect 78678 238711 78734 238720
rect 79336 223582 79364 286311
rect 79428 237386 79456 298279
rect 79520 252550 79548 310111
rect 79612 266354 79640 322079
rect 79704 280158 79732 333911
rect 504362 329624 504418 329633
rect 504362 329559 504418 329568
rect 504376 322930 504404 329559
rect 504364 322924 504416 322930
rect 504364 322866 504416 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 503810 318608 503866 318617
rect 503810 318543 503866 318552
rect 503824 311846 503852 318543
rect 503812 311840 503864 311846
rect 503812 311782 503864 311788
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 504362 307456 504418 307465
rect 504362 307391 504418 307400
rect 504376 299470 504404 307391
rect 504364 299464 504416 299470
rect 504364 299406 504416 299412
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 504362 296304 504418 296313
rect 504362 296239 504418 296248
rect 79692 280152 79744 280158
rect 79692 280094 79744 280100
rect 504376 276010 504404 296239
rect 504454 285288 504510 285297
rect 504454 285223 504510 285232
rect 504364 276004 504416 276010
rect 504364 275946 504416 275952
rect 504362 274136 504418 274145
rect 504362 274071 504418 274080
rect 79600 266348 79652 266354
rect 79600 266290 79652 266296
rect 79598 262576 79654 262585
rect 79598 262511 79654 262520
rect 79508 252544 79560 252550
rect 79508 252486 79560 252492
rect 79506 250744 79562 250753
rect 79506 250679 79562 250688
rect 79416 237380 79468 237386
rect 79416 237322 79468 237328
rect 79414 226944 79470 226953
rect 79414 226879 79470 226888
rect 79324 223576 79376 223582
rect 79324 223518 79376 223524
rect 79322 214976 79378 214985
rect 79322 214911 79378 214920
rect 78678 203144 78734 203153
rect 78678 203079 78734 203088
rect 78692 202910 78720 203079
rect 78680 202904 78732 202910
rect 78680 202846 78732 202852
rect 78678 167376 78734 167385
rect 78678 167311 78734 167320
rect 78692 167074 78720 167311
rect 78680 167068 78732 167074
rect 78680 167010 78732 167016
rect 25504 165572 25556 165578
rect 25504 165514 25556 165520
rect 79336 136610 79364 214911
rect 79428 151774 79456 226879
rect 79520 180810 79548 250679
rect 79612 194546 79640 262511
rect 504376 252550 504404 274071
rect 504468 264926 504496 285223
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 504456 264920 504508 264926
rect 504456 264862 504508 264868
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 504454 262984 504510 262993
rect 504454 262919 504510 262928
rect 504364 252544 504416 252550
rect 504364 252486 504416 252492
rect 504362 240816 504418 240825
rect 504362 240751 504418 240760
rect 504376 205630 504404 240751
rect 504468 229090 504496 262919
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 504730 251832 504786 251841
rect 504730 251767 504786 251776
rect 504546 229664 504602 229673
rect 504546 229599 504602 229608
rect 504456 229084 504508 229090
rect 504456 229026 504508 229032
rect 504454 207496 504510 207505
rect 504454 207431 504510 207440
rect 504364 205624 504416 205630
rect 504364 205566 504416 205572
rect 504362 196344 504418 196353
rect 504362 196279 504418 196288
rect 79600 194540 79652 194546
rect 79600 194482 79652 194488
rect 79782 191176 79838 191185
rect 79782 191111 79838 191120
rect 79508 180804 79560 180810
rect 79508 180746 79560 180752
rect 79690 179344 79746 179353
rect 79690 179279 79746 179288
rect 79598 155544 79654 155553
rect 79598 155479 79654 155488
rect 79416 151768 79468 151774
rect 79416 151710 79468 151716
rect 79506 143576 79562 143585
rect 79506 143511 79562 143520
rect 79324 136604 79376 136610
rect 79324 136546 79376 136552
rect 78678 131744 78734 131753
rect 78678 131679 78734 131688
rect 78692 131170 78720 131679
rect 78680 131164 78732 131170
rect 78680 131106 78732 131112
rect 24124 122800 24176 122806
rect 24124 122742 24176 122748
rect 79414 119776 79470 119785
rect 79414 119711 79470 119720
rect 79322 107944 79378 107953
rect 79322 107879 79378 107888
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 14464 35896 14516 35902
rect 3476 35864 3478 35873
rect 14464 35838 14516 35844
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 79336 8294 79364 107879
rect 79428 22098 79456 119711
rect 79520 51066 79548 143511
rect 79612 64870 79640 155479
rect 79704 93838 79732 179279
rect 79796 109002 79824 191111
rect 504376 135250 504404 196279
rect 504468 158710 504496 207431
rect 504560 182170 504588 229599
rect 504638 218512 504694 218521
rect 504638 218447 504694 218456
rect 504548 182164 504600 182170
rect 504548 182106 504600 182112
rect 504652 171086 504680 218447
rect 504744 218006 504772 251767
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 504732 218000 504784 218006
rect 504732 217942 504784 217948
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 504822 185192 504878 185201
rect 504822 185127 504878 185136
rect 504730 174176 504786 174185
rect 504730 174111 504786 174120
rect 504640 171080 504692 171086
rect 504640 171022 504692 171028
rect 504546 163024 504602 163033
rect 504546 162959 504602 162968
rect 504456 158704 504508 158710
rect 504456 158646 504508 158652
rect 504364 135244 504416 135250
rect 504364 135186 504416 135192
rect 504454 129704 504510 129713
rect 504454 129639 504510 129648
rect 504362 118552 504418 118561
rect 504362 118487 504418 118496
rect 79784 108996 79836 109002
rect 79784 108938 79836 108944
rect 504270 107536 504326 107545
rect 504270 107471 504326 107480
rect 504284 106350 504312 107471
rect 504272 106344 504324 106350
rect 504272 106286 504324 106292
rect 426282 102326 426480 102354
rect 92230 102190 92428 102218
rect 101982 102190 102180 102218
rect 148810 102190 149008 102218
rect 235842 102190 236040 102218
rect 81452 102054 82478 102082
rect 82832 102054 83490 102082
rect 79692 93832 79744 93838
rect 79692 93774 79744 93780
rect 79600 64864 79652 64870
rect 79600 64806 79652 64812
rect 79508 51060 79560 51066
rect 79508 51002 79560 51008
rect 79416 22092 79468 22098
rect 79416 22034 79468 22040
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 79324 8288 79376 8294
rect 79324 8230 79376 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 81452 3534 81480 102054
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 81440 3528 81492 3534
rect 81440 3470 81492 3476
rect 584 480 612 3470
rect 82832 3466 82860 102054
rect 84580 100706 84608 102068
rect 84568 100700 84620 100706
rect 84568 100642 84620 100648
rect 85488 100700 85540 100706
rect 85488 100642 85540 100648
rect 85500 4826 85528 100642
rect 85684 100026 85712 102068
rect 86696 102054 86802 102082
rect 87906 102054 88288 102082
rect 85672 100020 85724 100026
rect 85672 99962 85724 99968
rect 86696 96665 86724 102054
rect 86682 96656 86738 96665
rect 86682 96591 86738 96600
rect 86866 96656 86922 96665
rect 86866 96591 86922 96600
rect 86880 7682 86908 96591
rect 88260 8974 88288 102054
rect 88904 100706 88932 102068
rect 88892 100700 88944 100706
rect 88892 100642 88944 100648
rect 89628 100700 89680 100706
rect 89628 100642 89680 100648
rect 89640 28286 89668 100642
rect 90008 99618 90036 102068
rect 91112 100638 91140 102068
rect 92400 100722 92428 102190
rect 93334 102054 93808 102082
rect 92308 100694 92428 100722
rect 91100 100632 91152 100638
rect 91100 100574 91152 100580
rect 89996 99612 90048 99618
rect 89996 99554 90048 99560
rect 91008 99612 91060 99618
rect 91008 99554 91060 99560
rect 89628 28280 89680 28286
rect 89628 28222 89680 28228
rect 88248 8968 88300 8974
rect 88248 8910 88300 8916
rect 86868 7676 86920 7682
rect 86868 7618 86920 7624
rect 85488 4820 85540 4826
rect 85488 4762 85540 4768
rect 91020 4010 91048 99554
rect 92308 29646 92336 100694
rect 92388 100632 92440 100638
rect 92388 100574 92440 100580
rect 92296 29640 92348 29646
rect 92296 29582 92348 29588
rect 92400 11762 92428 100574
rect 92388 11756 92440 11762
rect 92388 11698 92440 11704
rect 91008 4004 91060 4010
rect 91008 3946 91060 3952
rect 93780 3942 93808 102054
rect 94424 100706 94452 102068
rect 95436 100706 95464 102068
rect 94412 100700 94464 100706
rect 94412 100642 94464 100648
rect 95148 100700 95200 100706
rect 95148 100642 95200 100648
rect 95424 100700 95476 100706
rect 95424 100642 95476 100648
rect 96436 100700 96488 100706
rect 96436 100642 96488 100648
rect 95160 10334 95188 100642
rect 96448 32434 96476 100642
rect 96436 32428 96488 32434
rect 96436 32370 96488 32376
rect 95148 10328 95200 10334
rect 95148 10270 95200 10276
rect 93768 3936 93820 3942
rect 93768 3878 93820 3884
rect 96540 3806 96568 102068
rect 97658 102054 97948 102082
rect 98762 102054 99328 102082
rect 97264 100020 97316 100026
rect 97264 99962 97316 99968
rect 97276 13122 97304 99962
rect 97920 14482 97948 102054
rect 99300 33794 99328 102054
rect 99852 100706 99880 102068
rect 100956 100706 100984 102068
rect 99840 100700 99892 100706
rect 99840 100642 99892 100648
rect 100668 100700 100720 100706
rect 100668 100642 100720 100648
rect 100944 100700 100996 100706
rect 100944 100642 100996 100648
rect 99288 33788 99340 33794
rect 99288 33730 99340 33736
rect 97908 14476 97960 14482
rect 97908 14418 97960 14424
rect 97264 13116 97316 13122
rect 97264 13058 97316 13064
rect 100680 3874 100708 100642
rect 102152 99362 102180 102190
rect 103086 102054 103468 102082
rect 104190 102054 104848 102082
rect 102784 100700 102836 100706
rect 102784 100642 102836 100648
rect 102060 99334 102180 99362
rect 102060 35222 102088 99334
rect 102048 35216 102100 35222
rect 102048 35158 102100 35164
rect 102796 15910 102824 100642
rect 102784 15904 102836 15910
rect 102784 15846 102836 15852
rect 100668 3868 100720 3874
rect 100668 3810 100720 3816
rect 96528 3800 96580 3806
rect 96528 3742 96580 3748
rect 103440 3738 103468 102054
rect 104820 17270 104848 102054
rect 105280 100706 105308 102068
rect 106384 100706 106412 102068
rect 105268 100700 105320 100706
rect 105268 100642 105320 100648
rect 106188 100700 106240 100706
rect 106188 100642 106240 100648
rect 106372 100700 106424 100706
rect 106372 100642 106424 100648
rect 106200 36582 106228 100642
rect 107488 99482 107516 102068
rect 108514 102054 108988 102082
rect 109618 102054 110368 102082
rect 107568 100700 107620 100706
rect 107568 100642 107620 100648
rect 107476 99476 107528 99482
rect 107476 99418 107528 99424
rect 106188 36576 106240 36582
rect 106188 36518 106240 36524
rect 104808 17264 104860 17270
rect 104808 17206 104860 17212
rect 103428 3732 103480 3738
rect 103428 3674 103480 3680
rect 107580 3670 107608 100642
rect 108960 37942 108988 102054
rect 108948 37936 109000 37942
rect 108948 37878 109000 37884
rect 107568 3664 107620 3670
rect 107568 3606 107620 3612
rect 110340 3602 110368 102054
rect 110708 99414 110736 102068
rect 110696 99408 110748 99414
rect 110696 99350 110748 99356
rect 111708 99408 111760 99414
rect 111708 99350 111760 99356
rect 111720 19990 111748 99350
rect 111812 97306 111840 102068
rect 112930 102054 113128 102082
rect 113942 102054 114508 102082
rect 111800 97300 111852 97306
rect 111800 97242 111852 97248
rect 111708 19984 111760 19990
rect 111708 19926 111760 19932
rect 110328 3596 110380 3602
rect 110328 3538 110380 3544
rect 113100 3466 113128 102054
rect 113824 99476 113876 99482
rect 113824 99418 113876 99424
rect 113836 18630 113864 99418
rect 114480 21418 114508 102054
rect 115032 99414 115060 102068
rect 116136 99414 116164 102068
rect 117240 100026 117268 102068
rect 118358 102054 118648 102082
rect 119462 102054 120028 102082
rect 117228 100020 117280 100026
rect 117228 99962 117280 99968
rect 115020 99408 115072 99414
rect 115020 99350 115072 99356
rect 115848 99408 115900 99414
rect 115848 99350 115900 99356
rect 116124 99408 116176 99414
rect 116124 99350 116176 99356
rect 117228 99408 117280 99414
rect 117228 99350 117280 99356
rect 115860 39370 115888 99350
rect 115848 39364 115900 39370
rect 115848 39306 115900 39312
rect 114468 21412 114520 21418
rect 114468 21354 114520 21360
rect 113824 18624 113876 18630
rect 113824 18566 113876 18572
rect 117240 3534 117268 99350
rect 118620 22778 118648 102054
rect 120000 40730 120028 102054
rect 120460 99414 120488 102068
rect 121564 99414 121592 102068
rect 120448 99408 120500 99414
rect 120448 99350 120500 99356
rect 121368 99408 121420 99414
rect 121368 99350 121420 99356
rect 121552 99408 121604 99414
rect 121552 99350 121604 99356
rect 119988 40724 120040 40730
rect 119988 40666 120040 40672
rect 118608 22772 118660 22778
rect 118608 22714 118660 22720
rect 121380 6254 121408 99350
rect 122668 42158 122696 102068
rect 123786 102054 124168 102082
rect 124890 102054 125548 102082
rect 122748 99408 122800 99414
rect 122748 99350 122800 99356
rect 122656 42152 122708 42158
rect 122656 42094 122708 42100
rect 122760 24138 122788 99350
rect 122748 24132 122800 24138
rect 122748 24074 122800 24080
rect 124140 7614 124168 102054
rect 125520 25634 125548 102054
rect 125980 99414 126008 102068
rect 126992 99414 127020 102068
rect 128110 102054 128308 102082
rect 129214 102054 129688 102082
rect 125968 99408 126020 99414
rect 125968 99350 126020 99356
rect 126888 99408 126940 99414
rect 126888 99350 126940 99356
rect 126980 99408 127032 99414
rect 126980 99350 127032 99356
rect 126900 43450 126928 99350
rect 126888 43444 126940 43450
rect 126888 43386 126940 43392
rect 128280 26994 128308 102054
rect 129004 99408 129056 99414
rect 129004 99350 129056 99356
rect 128268 26988 128320 26994
rect 128268 26930 128320 26936
rect 125508 25628 125560 25634
rect 125508 25570 125560 25576
rect 126980 13116 127032 13122
rect 126980 13058 127032 13064
rect 124128 7608 124180 7614
rect 124128 7550 124180 7556
rect 121368 6248 121420 6254
rect 121368 6190 121420 6196
rect 126612 4820 126664 4826
rect 126612 4762 126664 4768
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 82820 3460 82872 3466
rect 82820 3402 82872 3408
rect 113088 3460 113140 3466
rect 113088 3402 113140 3408
rect 1688 480 1716 3402
rect 126624 480 126652 4762
rect 126992 610 127020 13058
rect 128912 7676 128964 7682
rect 128912 7618 128964 7624
rect 128924 3482 128952 7618
rect 129016 4826 129044 99350
rect 129660 46238 129688 102054
rect 130304 99414 130332 102068
rect 131408 99414 131436 102068
rect 132512 99414 132540 102068
rect 133538 102054 133828 102082
rect 134642 102054 135208 102082
rect 130292 99408 130344 99414
rect 130292 99350 130344 99356
rect 131028 99408 131080 99414
rect 131028 99350 131080 99356
rect 131396 99408 131448 99414
rect 131396 99350 131448 99356
rect 132408 99408 132460 99414
rect 132408 99350 132460 99356
rect 132500 99408 132552 99414
rect 132500 99350 132552 99356
rect 133696 99408 133748 99414
rect 133696 99350 133748 99356
rect 129648 46232 129700 46238
rect 129648 46174 129700 46180
rect 131040 8974 131068 99350
rect 132420 28286 132448 99350
rect 133708 49094 133736 99350
rect 133696 49088 133748 49094
rect 133696 49030 133748 49036
rect 131120 28280 131172 28286
rect 131120 28222 131172 28228
rect 132408 28280 132460 28286
rect 132408 28222 132460 28228
rect 130200 8968 130252 8974
rect 130200 8910 130252 8916
rect 131028 8968 131080 8974
rect 131028 8910 131080 8916
rect 129004 4820 129056 4826
rect 129004 4762 129056 4768
rect 128924 3454 129044 3482
rect 126980 604 127032 610
rect 126980 546 127032 552
rect 127808 604 127860 610
rect 127808 546 127860 552
rect 127820 480 127848 546
rect 129016 480 129044 3454
rect 130212 480 130240 8910
rect 131132 610 131160 28222
rect 133800 11762 133828 102054
rect 135180 29714 135208 102054
rect 135732 99414 135760 102068
rect 136836 99414 136864 102068
rect 135720 99408 135772 99414
rect 135720 99350 135772 99356
rect 136548 99408 136600 99414
rect 136548 99350 136600 99356
rect 136824 99408 136876 99414
rect 136824 99350 136876 99356
rect 136560 50386 136588 99350
rect 136548 50380 136600 50386
rect 136548 50322 136600 50328
rect 137940 31074 137968 102068
rect 138966 102054 139348 102082
rect 140070 102054 140728 102082
rect 138664 99408 138716 99414
rect 138664 99350 138716 99356
rect 138020 32428 138072 32434
rect 138020 32370 138072 32376
rect 137928 31068 137980 31074
rect 137928 31010 137980 31016
rect 135168 29708 135220 29714
rect 135168 29650 135220 29656
rect 133880 29640 133932 29646
rect 133880 29582 133932 29588
rect 132592 11756 132644 11762
rect 132592 11698 132644 11704
rect 133788 11756 133840 11762
rect 133788 11698 133840 11704
rect 132500 4004 132552 4010
rect 132500 3946 132552 3952
rect 132512 3210 132540 3946
rect 132604 3398 132632 11698
rect 133892 3482 133920 29582
rect 136640 10328 136692 10334
rect 136640 10270 136692 10276
rect 136088 3936 136140 3942
rect 136088 3878 136140 3884
rect 133892 3454 134932 3482
rect 132592 3392 132644 3398
rect 132592 3334 132644 3340
rect 133788 3392 133840 3398
rect 133788 3334 133840 3340
rect 132512 3182 132632 3210
rect 131120 604 131172 610
rect 131120 546 131172 552
rect 131396 604 131448 610
rect 131396 546 131448 552
rect 131408 480 131436 546
rect 132604 480 132632 3182
rect 133800 480 133828 3334
rect 134904 480 134932 3454
rect 136100 480 136128 3878
rect 136652 3482 136680 10270
rect 138032 3482 138060 32370
rect 138676 10334 138704 99350
rect 139320 51746 139348 102054
rect 139308 51740 139360 51746
rect 139308 51682 139360 51688
rect 140700 13122 140728 102054
rect 141160 99414 141188 102068
rect 142264 99414 142292 102068
rect 143368 99498 143396 102068
rect 144486 102054 144868 102082
rect 145498 102054 146248 102082
rect 143368 99470 143488 99498
rect 141148 99408 141200 99414
rect 141148 99350 141200 99356
rect 142068 99408 142120 99414
rect 142068 99350 142120 99356
rect 142252 99408 142304 99414
rect 142252 99350 142304 99356
rect 143356 99408 143408 99414
rect 143356 99350 143408 99356
rect 140780 33788 140832 33794
rect 140780 33730 140832 33736
rect 140688 13116 140740 13122
rect 140688 13058 140740 13064
rect 138664 10328 138716 10334
rect 138664 10270 138716 10276
rect 139676 3800 139728 3806
rect 139676 3742 139728 3748
rect 136652 3454 137324 3482
rect 138032 3454 138520 3482
rect 137296 480 137324 3454
rect 138492 480 138520 3454
rect 139688 480 139716 3742
rect 140792 3058 140820 33730
rect 142080 32502 142108 99350
rect 143368 53106 143396 99350
rect 143356 53100 143408 53106
rect 143356 53042 143408 53048
rect 142068 32496 142120 32502
rect 142068 32438 142120 32444
rect 143460 14482 143488 99470
rect 144840 33862 144868 102054
rect 146220 54534 146248 102054
rect 146588 99414 146616 102068
rect 146576 99408 146628 99414
rect 146576 99350 146628 99356
rect 147588 99408 147640 99414
rect 147588 99350 147640 99356
rect 146208 54528 146260 54534
rect 146208 54470 146260 54476
rect 144920 35216 144972 35222
rect 144920 35158 144972 35164
rect 144828 33856 144880 33862
rect 144828 33798 144880 33804
rect 143540 15904 143592 15910
rect 143540 15846 143592 15852
rect 140872 14476 140924 14482
rect 140872 14418 140924 14424
rect 143448 14476 143500 14482
rect 143448 14418 143500 14424
rect 140780 3052 140832 3058
rect 140780 2994 140832 3000
rect 140884 480 140912 14418
rect 143264 3868 143316 3874
rect 143264 3810 143316 3816
rect 142068 3052 142120 3058
rect 142068 2994 142120 3000
rect 142080 480 142108 2994
rect 143276 480 143304 3810
rect 143552 3482 143580 15846
rect 144932 3482 144960 35158
rect 147600 15910 147628 99350
rect 147692 98666 147720 102068
rect 147680 98660 147732 98666
rect 147680 98602 147732 98608
rect 148980 96642 149008 102190
rect 149914 102054 150388 102082
rect 151018 102054 151768 102082
rect 148888 96614 149008 96642
rect 148888 89758 148916 96614
rect 148692 89752 148744 89758
rect 148876 89752 148928 89758
rect 148744 89700 148876 89706
rect 148692 89694 148928 89700
rect 148704 89678 148916 89694
rect 148888 77330 148916 89678
rect 148888 77302 149008 77330
rect 148980 77246 149008 77302
rect 148968 77240 149020 77246
rect 148968 77182 149020 77188
rect 148876 67652 148928 67658
rect 148876 67594 148928 67600
rect 148888 60858 148916 67594
rect 148876 60852 148928 60858
rect 148876 60794 148928 60800
rect 148784 60716 148836 60722
rect 148784 60658 148836 60664
rect 148796 55894 148824 60658
rect 148784 55888 148836 55894
rect 148784 55830 148836 55836
rect 149060 36576 149112 36582
rect 149060 36518 149112 36524
rect 147680 17264 147732 17270
rect 147680 17206 147732 17212
rect 147588 15904 147640 15910
rect 147588 15846 147640 15852
rect 146852 3732 146904 3738
rect 146852 3674 146904 3680
rect 143552 3454 144500 3482
rect 144932 3454 145696 3482
rect 144472 480 144500 3454
rect 145668 480 145696 3454
rect 146864 480 146892 3674
rect 147692 3482 147720 17206
rect 149072 3482 149100 36518
rect 150360 17270 150388 102054
rect 151740 35222 151768 102054
rect 152016 99414 152044 102068
rect 153120 100502 153148 102068
rect 154238 102054 154528 102082
rect 155342 102054 155908 102082
rect 153108 100496 153160 100502
rect 153108 100438 153160 100444
rect 153844 100496 153896 100502
rect 153844 100438 153896 100444
rect 152004 99408 152056 99414
rect 152004 99350 152056 99356
rect 153016 99340 153068 99346
rect 153016 99282 153068 99288
rect 153028 89706 153056 99282
rect 152936 89678 153056 89706
rect 152936 86970 152964 89678
rect 152924 86964 152976 86970
rect 152924 86906 152976 86912
rect 152832 77308 152884 77314
rect 152832 77250 152884 77256
rect 152844 77217 152872 77250
rect 152830 77208 152886 77217
rect 152830 77143 152886 77152
rect 153014 77208 153070 77217
rect 153014 77143 153070 77152
rect 153028 70446 153056 77143
rect 153016 70440 153068 70446
rect 153016 70382 153068 70388
rect 152924 70304 152976 70310
rect 152924 70246 152976 70252
rect 152936 57254 152964 70246
rect 152924 57248 152976 57254
rect 152924 57190 152976 57196
rect 151820 37936 151872 37942
rect 151820 37878 151872 37884
rect 151728 35216 151780 35222
rect 151728 35158 151780 35164
rect 150532 18624 150584 18630
rect 150532 18566 150584 18572
rect 150348 17264 150400 17270
rect 150348 17206 150400 17212
rect 150440 3664 150492 3670
rect 150440 3606 150492 3612
rect 147692 3454 148088 3482
rect 149072 3454 149284 3482
rect 148060 480 148088 3454
rect 149256 480 149284 3454
rect 150452 480 150480 3606
rect 150544 3482 150572 18566
rect 150544 3454 151584 3482
rect 151556 480 151584 3454
rect 151832 3346 151860 37878
rect 153856 18630 153884 100438
rect 154500 36650 154528 102054
rect 155880 58682 155908 102054
rect 156432 100706 156460 102068
rect 156420 100700 156472 100706
rect 156420 100642 156472 100648
rect 157248 100700 157300 100706
rect 157248 100642 157300 100648
rect 155960 97300 156012 97306
rect 155960 97242 156012 97248
rect 155868 58676 155920 58682
rect 155868 58618 155920 58624
rect 154488 36644 154540 36650
rect 154488 36586 154540 36592
rect 154580 19984 154632 19990
rect 154580 19926 154632 19932
rect 153844 18624 153896 18630
rect 153844 18566 153896 18572
rect 153936 3596 153988 3602
rect 153936 3538 153988 3544
rect 151832 3318 152780 3346
rect 152752 480 152780 3318
rect 153948 480 153976 3538
rect 154592 3346 154620 19926
rect 155972 3346 156000 97242
rect 157260 19990 157288 100642
rect 157536 99414 157564 102068
rect 157524 99408 157576 99414
rect 157524 99350 157576 99356
rect 158548 61402 158576 102068
rect 159666 102054 160048 102082
rect 160770 102054 161428 102082
rect 158628 99408 158680 99414
rect 158628 99350 158680 99356
rect 158536 61396 158588 61402
rect 158536 61338 158588 61344
rect 158640 37942 158668 99350
rect 158720 39364 158772 39370
rect 158720 39306 158772 39312
rect 158628 37936 158680 37942
rect 158628 37878 158680 37884
rect 157248 19984 157300 19990
rect 157248 19926 157300 19932
rect 158732 3534 158760 39306
rect 158812 21412 158864 21418
rect 158812 21354 158864 21360
rect 158720 3528 158772 3534
rect 158720 3470 158772 3476
rect 157524 3460 157576 3466
rect 157524 3402 157576 3408
rect 154592 3318 155172 3346
rect 155972 3318 156368 3346
rect 155144 480 155172 3318
rect 156340 480 156368 3318
rect 157536 480 157564 3402
rect 158824 1442 158852 21354
rect 160020 6186 160048 102054
rect 161400 22846 161428 102054
rect 161572 100020 161624 100026
rect 161572 99962 161624 99968
rect 161388 22840 161440 22846
rect 161388 22782 161440 22788
rect 160008 6180 160060 6186
rect 160008 6122 160060 6128
rect 159916 3528 159968 3534
rect 159916 3470 159968 3476
rect 161584 3482 161612 99962
rect 161860 99414 161888 102068
rect 162964 100026 162992 102068
rect 163990 102054 164188 102082
rect 165094 102054 165568 102082
rect 162952 100020 163004 100026
rect 162952 99962 163004 99968
rect 161848 99408 161900 99414
rect 161848 99350 161900 99356
rect 162768 99408 162820 99414
rect 162768 99350 162820 99356
rect 162780 39370 162808 99350
rect 164160 47598 164188 102054
rect 164148 47592 164200 47598
rect 164148 47534 164200 47540
rect 165540 42090 165568 102054
rect 166184 99414 166212 102068
rect 167288 99414 167316 102068
rect 168392 99414 168420 102068
rect 169510 102054 169708 102082
rect 170522 102054 171088 102082
rect 166172 99408 166224 99414
rect 166172 99350 166224 99356
rect 166908 99408 166960 99414
rect 166908 99350 166960 99356
rect 167276 99408 167328 99414
rect 167276 99350 167328 99356
rect 168288 99408 168340 99414
rect 168288 99350 168340 99356
rect 168380 99408 168432 99414
rect 168380 99350 168432 99356
rect 169576 99408 169628 99414
rect 169576 99350 169628 99356
rect 165528 42084 165580 42090
rect 165528 42026 165580 42032
rect 164240 40724 164292 40730
rect 164240 40666 164292 40672
rect 162768 39364 162820 39370
rect 162768 39306 162820 39312
rect 162860 22772 162912 22778
rect 162860 22714 162912 22720
rect 162872 3482 162900 22714
rect 164252 3482 164280 40666
rect 166920 21418 166948 99350
rect 167000 42152 167052 42158
rect 167000 42094 167052 42100
rect 166908 21412 166960 21418
rect 166908 21354 166960 21360
rect 165896 6248 165948 6254
rect 165896 6190 165948 6196
rect 158732 1414 158852 1442
rect 158732 480 158760 1414
rect 159928 480 159956 3470
rect 161112 3460 161164 3466
rect 161584 3454 162348 3482
rect 162872 3454 163544 3482
rect 164252 3454 164740 3482
rect 161112 3402 161164 3408
rect 161124 480 161152 3402
rect 162320 480 162348 3454
rect 163516 480 163544 3454
rect 164712 480 164740 3454
rect 165908 480 165936 6190
rect 167012 3534 167040 42094
rect 168300 25566 168328 99350
rect 169588 60042 169616 99350
rect 169576 60036 169628 60042
rect 169576 59978 169628 59984
rect 169680 44878 169708 102054
rect 169668 44872 169720 44878
rect 169668 44814 169720 44820
rect 171060 26926 171088 102054
rect 171612 99414 171640 102068
rect 172716 99414 172744 102068
rect 173728 102054 173834 102082
rect 174938 102054 175228 102082
rect 176042 102054 176608 102082
rect 171600 99408 171652 99414
rect 171600 99350 171652 99356
rect 172428 99408 172480 99414
rect 172428 99350 172480 99356
rect 172704 99408 172756 99414
rect 172704 99350 172756 99356
rect 172440 62830 172468 99350
rect 172428 62824 172480 62830
rect 172428 62766 172480 62772
rect 171140 43444 171192 43450
rect 171140 43386 171192 43392
rect 171048 26920 171100 26926
rect 171048 26862 171100 26868
rect 169760 25628 169812 25634
rect 169760 25570 169812 25576
rect 168288 25560 168340 25566
rect 168288 25502 168340 25508
rect 167092 24132 167144 24138
rect 167092 24074 167144 24080
rect 167000 3528 167052 3534
rect 167000 3470 167052 3476
rect 167104 480 167132 24074
rect 169392 7608 169444 7614
rect 169392 7550 169444 7556
rect 168196 3528 168248 3534
rect 168196 3470 168248 3476
rect 168208 480 168236 3470
rect 169404 480 169432 7550
rect 169772 3482 169800 25570
rect 171152 3482 171180 43386
rect 173728 40730 173756 102054
rect 173808 99408 173860 99414
rect 173808 99350 173860 99356
rect 173716 40724 173768 40730
rect 173716 40666 173768 40672
rect 173820 4826 173848 99350
rect 175200 49026 175228 102054
rect 175188 49020 175240 49026
rect 175188 48962 175240 48968
rect 175280 46232 175332 46238
rect 175280 46174 175332 46180
rect 173900 26988 173952 26994
rect 173900 26930 173952 26936
rect 172980 4820 173032 4826
rect 172980 4762 173032 4768
rect 173808 4820 173860 4826
rect 173808 4762 173860 4768
rect 169772 3454 170628 3482
rect 171152 3454 171824 3482
rect 170600 480 170628 3454
rect 171796 480 171824 3454
rect 172992 480 173020 4762
rect 173912 3482 173940 26930
rect 175292 3482 175320 46174
rect 176580 12050 176608 102054
rect 177040 99414 177068 102068
rect 178144 99414 178172 102068
rect 179248 99498 179276 102068
rect 180366 102054 180748 102082
rect 181470 102054 182128 102082
rect 179248 99470 179368 99498
rect 177028 99408 177080 99414
rect 177028 99350 177080 99356
rect 177948 99408 178000 99414
rect 177948 99350 178000 99356
rect 178132 99408 178184 99414
rect 178132 99350 178184 99356
rect 179236 99408 179288 99414
rect 179236 99350 179288 99356
rect 177960 28286 177988 99350
rect 179248 64258 179276 99350
rect 179236 64252 179288 64258
rect 179236 64194 179288 64200
rect 178040 49088 178092 49094
rect 178040 49030 178092 49036
rect 176660 28280 176712 28286
rect 176660 28222 176712 28228
rect 177948 28280 178000 28286
rect 177948 28222 178000 28228
rect 176396 12022 176608 12050
rect 176396 7614 176424 12022
rect 176568 8968 176620 8974
rect 176568 8910 176620 8916
rect 176384 7608 176436 7614
rect 176384 7550 176436 7556
rect 173912 3454 174216 3482
rect 175292 3454 175412 3482
rect 174188 480 174216 3454
rect 175384 480 175412 3454
rect 176580 480 176608 8910
rect 176672 3482 176700 28222
rect 178052 3482 178080 49030
rect 179340 8974 179368 99470
rect 180720 29646 180748 102054
rect 182100 65550 182128 102054
rect 182560 99414 182588 102068
rect 183572 99414 183600 102068
rect 184690 102054 184888 102082
rect 185794 102054 186268 102082
rect 186898 102054 187648 102082
rect 182548 99408 182600 99414
rect 182548 99350 182600 99356
rect 183468 99408 183520 99414
rect 183468 99350 183520 99356
rect 183560 99408 183612 99414
rect 183560 99350 183612 99356
rect 182088 65544 182140 65550
rect 182088 65486 182140 65492
rect 182180 50380 182232 50386
rect 182180 50322 182232 50328
rect 180800 29708 180852 29714
rect 180800 29650 180852 29656
rect 180708 29640 180760 29646
rect 180708 29582 180760 29588
rect 179420 11756 179472 11762
rect 179420 11698 179472 11704
rect 179328 8968 179380 8974
rect 179328 8910 179380 8916
rect 179432 3482 179460 11698
rect 180812 3482 180840 29650
rect 182192 3482 182220 50322
rect 183480 11762 183508 99350
rect 184860 66910 184888 102054
rect 185584 99408 185636 99414
rect 185584 99350 185636 99356
rect 184848 66904 184900 66910
rect 184848 66846 184900 66852
rect 184940 51740 184992 51746
rect 184940 51682 184992 51688
rect 183560 31068 183612 31074
rect 183560 31010 183612 31016
rect 183468 11756 183520 11762
rect 183468 11698 183520 11704
rect 183572 3534 183600 31010
rect 183652 10328 183704 10334
rect 183652 10270 183704 10276
rect 183560 3528 183612 3534
rect 176672 3454 177804 3482
rect 178052 3454 179000 3482
rect 179432 3454 180196 3482
rect 180812 3454 181392 3482
rect 182192 3454 182588 3482
rect 183560 3470 183612 3476
rect 183664 3482 183692 10270
rect 184848 3528 184900 3534
rect 183664 3454 183784 3482
rect 184848 3470 184900 3476
rect 184952 3482 184980 51682
rect 185596 31074 185624 99350
rect 185584 31068 185636 31074
rect 185584 31010 185636 31016
rect 186240 10334 186268 102054
rect 187620 32434 187648 102054
rect 187988 99414 188016 102068
rect 189000 99414 189028 102068
rect 190118 102054 190408 102082
rect 191222 102054 191788 102082
rect 187976 99408 188028 99414
rect 187976 99350 188028 99356
rect 188988 99408 189040 99414
rect 188988 99350 189040 99356
rect 189724 99408 189776 99414
rect 189724 99350 189776 99356
rect 188988 99272 189040 99278
rect 188988 99214 189040 99220
rect 189000 93786 189028 99214
rect 188908 93758 189028 93786
rect 188908 89706 188936 93758
rect 188724 89678 188936 89706
rect 188724 82142 188752 89678
rect 188712 82136 188764 82142
rect 188712 82078 188764 82084
rect 188896 82136 188948 82142
rect 188896 82078 188948 82084
rect 188908 77353 188936 82078
rect 188710 77344 188766 77353
rect 188632 77302 188710 77330
rect 188632 77246 188660 77302
rect 188710 77279 188766 77288
rect 188894 77344 188950 77353
rect 188894 77279 188950 77288
rect 188620 77240 188672 77246
rect 188620 77182 188672 77188
rect 188528 67652 188580 67658
rect 188528 67594 188580 67600
rect 188540 60738 188568 67594
rect 188540 60710 188752 60738
rect 188724 51746 188752 60710
rect 189080 53100 189132 53106
rect 189080 53042 189132 53048
rect 188712 51740 188764 51746
rect 188712 51682 188764 51688
rect 187700 32496 187752 32502
rect 187700 32438 187752 32444
rect 187608 32428 187660 32434
rect 187608 32370 187660 32376
rect 186320 13116 186372 13122
rect 186320 13058 186372 13064
rect 186228 10328 186280 10334
rect 186228 10270 186280 10276
rect 186332 3482 186360 13058
rect 187712 3482 187740 32438
rect 189092 3482 189120 53042
rect 189736 13122 189764 99350
rect 190380 33794 190408 102054
rect 191760 53174 191788 102054
rect 192312 99414 192340 102068
rect 193416 99414 193444 102068
rect 194428 102054 194534 102082
rect 195546 102054 195928 102082
rect 196650 102054 197308 102082
rect 192300 99408 192352 99414
rect 192300 99350 192352 99356
rect 193128 99408 193180 99414
rect 193128 99350 193180 99356
rect 193404 99408 193456 99414
rect 193404 99350 193456 99356
rect 191748 53168 191800 53174
rect 191748 53110 191800 53116
rect 191840 33856 191892 33862
rect 191840 33798 191892 33804
rect 190368 33788 190420 33794
rect 190368 33730 190420 33736
rect 190460 14476 190512 14482
rect 190460 14418 190512 14424
rect 189724 13116 189776 13122
rect 189724 13058 189776 13064
rect 190472 3482 190500 14418
rect 191852 3482 191880 33798
rect 193140 14482 193168 99350
rect 194428 54602 194456 102054
rect 194508 99408 194560 99414
rect 194508 99350 194560 99356
rect 194416 54596 194468 54602
rect 194416 54538 194468 54544
rect 193220 54528 193272 54534
rect 193220 54470 193272 54476
rect 193128 14476 193180 14482
rect 193128 14418 193180 14424
rect 177776 480 177804 3454
rect 178972 480 179000 3454
rect 180168 480 180196 3454
rect 181364 480 181392 3454
rect 182560 480 182588 3454
rect 183756 480 183784 3454
rect 184860 480 184888 3470
rect 184952 3454 186084 3482
rect 186332 3454 187280 3482
rect 187712 3454 188476 3482
rect 189092 3454 189672 3482
rect 190472 3454 190868 3482
rect 191852 3454 192064 3482
rect 186056 480 186084 3454
rect 187252 480 187280 3454
rect 188448 480 188476 3454
rect 189644 480 189672 3454
rect 190840 480 190868 3454
rect 192036 480 192064 3454
rect 193232 480 193260 54470
rect 194520 43450 194548 99350
rect 194600 98660 194652 98666
rect 194600 98602 194652 98608
rect 194508 43444 194560 43450
rect 194508 43386 194560 43392
rect 193312 15904 193364 15910
rect 193312 15846 193364 15852
rect 193324 3482 193352 15846
rect 194612 3482 194640 98602
rect 195900 15910 195928 102054
rect 195980 55888 196032 55894
rect 195980 55830 196032 55836
rect 195888 15904 195940 15910
rect 195888 15846 195940 15852
rect 195992 3482 196020 55830
rect 197280 46238 197308 102054
rect 197740 99414 197768 102068
rect 197728 99408 197780 99414
rect 197728 99350 197780 99356
rect 198648 99408 198700 99414
rect 198648 99350 198700 99356
rect 197268 46232 197320 46238
rect 197268 46174 197320 46180
rect 198660 36582 198688 99350
rect 198844 98666 198872 102068
rect 198832 98660 198884 98666
rect 198832 98602 198884 98608
rect 198648 36576 198700 36582
rect 198648 36518 198700 36524
rect 199948 35222 199976 102068
rect 201066 102054 201448 102082
rect 200120 57248 200172 57254
rect 200120 57190 200172 57196
rect 198740 35216 198792 35222
rect 198740 35158 198792 35164
rect 199936 35216 199988 35222
rect 199936 35158 199988 35164
rect 197360 17264 197412 17270
rect 197360 17206 197412 17212
rect 197372 3482 197400 17206
rect 198752 3482 198780 35158
rect 200132 3482 200160 57190
rect 201420 55962 201448 102054
rect 202064 99414 202092 102068
rect 203168 99414 203196 102068
rect 204272 99414 204300 102068
rect 205390 102054 205588 102082
rect 206494 102054 206968 102082
rect 202052 99408 202104 99414
rect 202052 99350 202104 99356
rect 202788 99408 202840 99414
rect 202788 99350 202840 99356
rect 203156 99408 203208 99414
rect 203156 99350 203208 99356
rect 204168 99408 204220 99414
rect 204168 99350 204220 99356
rect 204260 99408 204312 99414
rect 204260 99350 204312 99356
rect 205456 99408 205508 99414
rect 205456 99350 205508 99356
rect 201408 55956 201460 55962
rect 201408 55898 201460 55904
rect 201500 36644 201552 36650
rect 201500 36586 201552 36592
rect 201512 3602 201540 36586
rect 202800 24206 202828 99350
rect 202880 58676 202932 58682
rect 202880 58618 202932 58624
rect 202788 24200 202840 24206
rect 202788 24142 202840 24148
rect 201592 18624 201644 18630
rect 201592 18566 201644 18572
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 201604 3482 201632 18566
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 193324 3454 194456 3482
rect 194612 3454 195652 3482
rect 195992 3454 196848 3482
rect 197372 3454 198044 3482
rect 198752 3454 199240 3482
rect 200132 3454 200436 3482
rect 194428 480 194456 3454
rect 195624 480 195652 3454
rect 196820 480 196848 3454
rect 198016 480 198044 3454
rect 199212 480 199240 3454
rect 200408 480 200436 3454
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202708 480 202736 3538
rect 202892 3482 202920 58618
rect 204180 22778 204208 99350
rect 205468 57322 205496 99350
rect 205456 57316 205508 57322
rect 205456 57258 205508 57264
rect 204168 22772 204220 22778
rect 204168 22714 204220 22720
rect 205560 19990 205588 102054
rect 206940 37942 206968 102054
rect 207584 99414 207612 102068
rect 208596 99414 208624 102068
rect 209608 102054 209714 102082
rect 210818 102054 211108 102082
rect 207572 99408 207624 99414
rect 207572 99350 207624 99356
rect 208308 99408 208360 99414
rect 208308 99350 208360 99356
rect 208584 99408 208636 99414
rect 208584 99350 208636 99356
rect 207020 61396 207072 61402
rect 207020 61338 207072 61344
rect 205640 37936 205692 37942
rect 205640 37878 205692 37884
rect 206928 37936 206980 37942
rect 206928 37878 206980 37884
rect 204260 19984 204312 19990
rect 204260 19926 204312 19932
rect 205548 19984 205600 19990
rect 205548 19926 205600 19932
rect 204272 3482 204300 19926
rect 205652 3482 205680 37878
rect 207032 3482 207060 61338
rect 208320 58682 208348 99350
rect 208308 58676 208360 58682
rect 208308 58618 208360 58624
rect 209608 50386 209636 102054
rect 209688 99408 209740 99414
rect 209688 99350 209740 99356
rect 209596 50380 209648 50386
rect 209596 50322 209648 50328
rect 209700 17270 209728 99350
rect 211080 61470 211108 102054
rect 211908 100094 211936 102068
rect 211896 100088 211948 100094
rect 211896 100030 211948 100036
rect 211160 100020 211212 100026
rect 211160 99962 211212 99968
rect 211068 61464 211120 61470
rect 211068 61406 211120 61412
rect 209780 39364 209832 39370
rect 209780 39306 209832 39312
rect 209688 17264 209740 17270
rect 209688 17206 209740 17212
rect 208676 6180 208728 6186
rect 208676 6122 208728 6128
rect 202892 3454 203932 3482
rect 204272 3454 205128 3482
rect 205652 3454 206324 3482
rect 207032 3454 207520 3482
rect 203904 480 203932 3454
rect 205100 480 205128 3454
rect 206296 480 206324 3454
rect 207492 480 207520 3454
rect 208688 480 208716 6122
rect 209792 3534 209820 39306
rect 209872 22840 209924 22846
rect 209872 22782 209924 22788
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 209884 480 209912 22782
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 211172 3482 211200 99962
rect 213012 99414 213040 102068
rect 214024 99414 214052 102068
rect 215128 99498 215156 102068
rect 216246 102054 216628 102082
rect 217350 102054 218008 102082
rect 215128 99470 215248 99498
rect 213000 99408 213052 99414
rect 213000 99350 213052 99356
rect 213828 99408 213880 99414
rect 213828 99350 213880 99356
rect 214012 99408 214064 99414
rect 214012 99350 214064 99356
rect 215116 99408 215168 99414
rect 215116 99350 215168 99356
rect 213840 47598 213868 99350
rect 215128 68338 215156 99350
rect 215116 68332 215168 68338
rect 215116 68274 215168 68280
rect 212540 47592 212592 47598
rect 212540 47534 212592 47540
rect 213828 47592 213880 47598
rect 213828 47534 213880 47540
rect 212552 3482 212580 47534
rect 213920 42084 213972 42090
rect 213920 42026 213972 42032
rect 213932 3482 213960 42026
rect 215220 39370 215248 99470
rect 215208 39364 215260 39370
rect 215208 39306 215260 39312
rect 216600 25634 216628 102054
rect 217980 60110 218008 102054
rect 218440 99414 218468 102068
rect 218428 99408 218480 99414
rect 218428 99350 218480 99356
rect 219348 99408 219400 99414
rect 219348 99350 219400 99356
rect 217968 60104 218020 60110
rect 217968 60046 218020 60052
rect 218060 60036 218112 60042
rect 218060 59978 218112 59984
rect 216588 25628 216640 25634
rect 216588 25570 216640 25576
rect 216680 25560 216732 25566
rect 216680 25502 216732 25508
rect 215300 21412 215352 21418
rect 215300 21354 215352 21360
rect 215312 3482 215340 21354
rect 216692 3482 216720 25502
rect 218072 3482 218100 59978
rect 218152 44872 218204 44878
rect 218152 44814 218204 44820
rect 218164 3602 218192 44814
rect 219360 6186 219388 99350
rect 219544 95946 219572 102068
rect 220556 99414 220584 102068
rect 221674 102054 222148 102082
rect 222778 102054 223528 102082
rect 220544 99408 220596 99414
rect 220544 99350 220596 99356
rect 221464 99408 221516 99414
rect 221464 99350 221516 99356
rect 219532 95940 219584 95946
rect 219532 95882 219584 95888
rect 221476 62830 221504 99350
rect 220820 62824 220872 62830
rect 220820 62766 220872 62772
rect 221464 62824 221516 62830
rect 221464 62766 221516 62772
rect 219440 26920 219492 26926
rect 219440 26862 219492 26868
rect 219348 6180 219400 6186
rect 219348 6122 219400 6128
rect 218152 3596 218204 3602
rect 218152 3538 218204 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 211080 480 211108 3470
rect 211172 3454 212304 3482
rect 212552 3454 213500 3482
rect 213932 3454 214696 3482
rect 215312 3454 215892 3482
rect 216692 3454 217088 3482
rect 218072 3454 218192 3482
rect 212276 480 212304 3454
rect 213472 480 213500 3454
rect 214668 480 214696 3454
rect 215864 480 215892 3454
rect 217060 480 217088 3454
rect 218164 480 218192 3454
rect 219360 480 219388 3538
rect 219452 3482 219480 26862
rect 220832 3482 220860 62766
rect 222120 18630 222148 102054
rect 223500 26926 223528 102054
rect 223868 99414 223896 102068
rect 224972 99822 225000 102068
rect 225984 102054 226090 102082
rect 227102 102054 227668 102082
rect 224960 99816 225012 99822
rect 224960 99758 225012 99764
rect 223856 99408 223908 99414
rect 223856 99350 223908 99356
rect 224868 99408 224920 99414
rect 224868 99350 224920 99356
rect 224880 71058 224908 99350
rect 225984 96665 226012 102054
rect 226248 99816 226300 99822
rect 226248 99758 226300 99764
rect 225970 96656 226026 96665
rect 225970 96591 226026 96600
rect 226154 96656 226210 96665
rect 226154 96591 226210 96600
rect 226168 89758 226196 96591
rect 225972 89752 226024 89758
rect 225972 89694 226024 89700
rect 226156 89752 226208 89758
rect 226156 89694 226208 89700
rect 225984 77246 226012 89694
rect 225972 77240 226024 77246
rect 225972 77182 226024 77188
rect 224868 71052 224920 71058
rect 224868 70994 224920 71000
rect 225880 67652 225932 67658
rect 225880 67594 225932 67600
rect 225892 60738 225920 67594
rect 225892 60710 226104 60738
rect 226076 51082 226104 60710
rect 225984 51054 226104 51082
rect 225984 49026 226012 51054
rect 224960 49020 225012 49026
rect 224960 48962 225012 48968
rect 225972 49020 226024 49026
rect 225972 48962 226024 48968
rect 223580 40724 223632 40730
rect 223580 40666 223632 40672
rect 223488 26920 223540 26926
rect 223488 26862 223540 26868
rect 222108 18624 222160 18630
rect 222108 18566 222160 18572
rect 222936 4820 222988 4826
rect 222936 4762 222988 4768
rect 219452 3454 220584 3482
rect 220832 3454 221780 3482
rect 220556 480 220584 3454
rect 221752 480 221780 3454
rect 222948 480 222976 4762
rect 223592 3482 223620 40666
rect 224972 3482 225000 48962
rect 226260 21486 226288 99758
rect 227640 64190 227668 102054
rect 228192 100706 228220 102068
rect 229296 100706 229324 102068
rect 230308 102054 230414 102082
rect 228180 100700 228232 100706
rect 228180 100642 228232 100648
rect 229008 100700 229060 100706
rect 229008 100642 229060 100648
rect 229284 100700 229336 100706
rect 229284 100642 229336 100648
rect 227720 64252 227772 64258
rect 227720 64194 227772 64200
rect 227628 64184 227680 64190
rect 227628 64126 227680 64132
rect 226248 21480 226300 21486
rect 226248 21422 226300 21428
rect 226524 7608 226576 7614
rect 226524 7550 226576 7556
rect 223592 3454 224172 3482
rect 224972 3454 225368 3482
rect 224144 480 224172 3454
rect 225340 480 225368 3454
rect 226536 480 226564 7550
rect 227732 3602 227760 64194
rect 229020 42090 229048 100642
rect 230308 69698 230336 102054
rect 230388 100700 230440 100706
rect 230388 100642 230440 100648
rect 230296 69692 230348 69698
rect 230296 69634 230348 69640
rect 229008 42084 229060 42090
rect 229008 42026 229060 42032
rect 230400 40730 230428 100642
rect 231124 100088 231176 100094
rect 231124 100030 231176 100036
rect 230388 40724 230440 40730
rect 230388 40666 230440 40672
rect 230480 29640 230532 29646
rect 230480 29582 230532 29588
rect 227812 28280 227864 28286
rect 227812 28222 227864 28228
rect 227720 3596 227772 3602
rect 227720 3538 227772 3544
rect 227824 3482 227852 28222
rect 230112 8968 230164 8974
rect 230112 8910 230164 8916
rect 228916 3596 228968 3602
rect 228916 3538 228968 3544
rect 227732 3454 227852 3482
rect 227732 480 227760 3454
rect 228928 480 228956 3538
rect 230124 480 230152 8910
rect 230492 3618 230520 29582
rect 231136 4894 231164 100030
rect 231504 100026 231532 102068
rect 232622 102054 233188 102082
rect 231492 100020 231544 100026
rect 231492 99962 231544 99968
rect 231860 65544 231912 65550
rect 231860 65486 231912 65492
rect 231124 4888 231176 4894
rect 231124 4830 231176 4836
rect 230492 3590 231348 3618
rect 231320 480 231348 3590
rect 231872 3482 231900 65486
rect 233160 28286 233188 102054
rect 233620 100706 233648 102068
rect 233608 100700 233660 100706
rect 233608 100642 233660 100648
rect 234528 100700 234580 100706
rect 234528 100642 234580 100648
rect 234540 65550 234568 100642
rect 234724 97306 234752 102068
rect 234712 97300 234764 97306
rect 234712 97242 234764 97248
rect 236012 96642 236040 102190
rect 328104 102190 328302 102218
rect 395830 102190 396028 102218
rect 411010 102190 411208 102218
rect 236946 102054 237328 102082
rect 238050 102054 238708 102082
rect 235920 96614 236040 96642
rect 235920 89758 235948 96614
rect 235724 89752 235776 89758
rect 235724 89694 235776 89700
rect 235908 89752 235960 89758
rect 235908 89694 235960 89700
rect 235736 77246 235764 89694
rect 235724 77240 235776 77246
rect 235724 77182 235776 77188
rect 235632 67652 235684 67658
rect 235632 67594 235684 67600
rect 234528 65544 234580 65550
rect 234528 65486 234580 65492
rect 235644 60738 235672 67594
rect 237300 66978 237328 102054
rect 237288 66972 237340 66978
rect 237288 66914 237340 66920
rect 236000 66904 236052 66910
rect 236000 66846 236052 66852
rect 235644 60710 235856 60738
rect 235828 50454 235856 60710
rect 235816 50448 235868 50454
rect 235816 50390 235868 50396
rect 235908 45620 235960 45626
rect 235908 45562 235960 45568
rect 235920 45506 235948 45562
rect 235828 45478 235948 45506
rect 235828 41478 235856 45478
rect 235816 41472 235868 41478
rect 235816 41414 235868 41420
rect 234620 31068 234672 31074
rect 234620 31010 234672 31016
rect 233148 28280 233200 28286
rect 233148 28222 233200 28228
rect 233240 11756 233292 11762
rect 233240 11698 233292 11704
rect 233252 3482 233280 11698
rect 234632 3482 234660 31010
rect 231872 3454 232544 3482
rect 233252 3454 233740 3482
rect 234632 3454 234844 3482
rect 232516 480 232544 3454
rect 233712 480 233740 3454
rect 234816 480 234844 3454
rect 236012 480 236040 66846
rect 237380 32428 237432 32434
rect 237380 32370 237432 32376
rect 236092 10328 236144 10334
rect 236092 10270 236144 10276
rect 236104 3482 236132 10270
rect 237392 3482 237420 32370
rect 238680 7614 238708 102054
rect 239140 99754 239168 102068
rect 240152 100638 240180 102068
rect 241270 102054 241468 102082
rect 242374 102054 242848 102082
rect 240140 100632 240192 100638
rect 240140 100574 240192 100580
rect 241336 100632 241388 100638
rect 241336 100574 241388 100580
rect 239128 99748 239180 99754
rect 239128 99690 239180 99696
rect 240048 99748 240100 99754
rect 240048 99690 240100 99696
rect 238760 51740 238812 51746
rect 238760 51682 238812 51688
rect 238668 7608 238720 7614
rect 238668 7550 238720 7556
rect 238772 3482 238800 51682
rect 240060 31074 240088 99690
rect 241348 53106 241376 100574
rect 241336 53100 241388 53106
rect 241336 53042 241388 53048
rect 240048 31068 240100 31074
rect 240048 31010 240100 31016
rect 240140 13116 240192 13122
rect 240140 13058 240192 13064
rect 240152 3482 240180 13058
rect 241440 11762 241468 102054
rect 242820 51746 242848 102054
rect 243464 100706 243492 102068
rect 243452 100700 243504 100706
rect 243452 100642 243504 100648
rect 244188 100700 244240 100706
rect 244188 100642 244240 100648
rect 244200 54534 244228 100642
rect 244568 99414 244596 102068
rect 245488 102054 245594 102082
rect 246698 102054 246988 102082
rect 247802 102054 248368 102082
rect 244556 99408 244608 99414
rect 244556 99350 244608 99356
rect 244188 54528 244240 54534
rect 244188 54470 244240 54476
rect 242900 53168 242952 53174
rect 242900 53110 242952 53116
rect 242808 51740 242860 51746
rect 242808 51682 242860 51688
rect 241520 33788 241572 33794
rect 241520 33730 241572 33736
rect 241428 11756 241480 11762
rect 241428 11698 241480 11704
rect 241532 3482 241560 33730
rect 242912 3482 242940 53110
rect 245488 43450 245516 102054
rect 245568 99408 245620 99414
rect 245568 99350 245620 99356
rect 244280 43444 244332 43450
rect 244280 43386 244332 43392
rect 245476 43444 245528 43450
rect 245476 43386 245528 43392
rect 244292 3534 244320 43386
rect 244372 14476 244424 14482
rect 244372 14418 244424 14424
rect 244280 3528 244332 3534
rect 236104 3454 237236 3482
rect 237392 3454 238432 3482
rect 238772 3454 239628 3482
rect 240152 3454 240824 3482
rect 241532 3454 242020 3482
rect 242912 3454 243216 3482
rect 244280 3470 244332 3476
rect 237208 480 237236 3454
rect 238404 480 238432 3454
rect 239600 480 239628 3454
rect 240796 480 240824 3454
rect 241992 480 242020 3454
rect 243188 480 243216 3454
rect 244384 480 244412 14418
rect 245580 8974 245608 99350
rect 246960 72486 246988 102054
rect 246948 72480 247000 72486
rect 246948 72422 247000 72428
rect 245660 54596 245712 54602
rect 245660 54538 245712 54544
rect 245568 8968 245620 8974
rect 245568 8910 245620 8916
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245672 3482 245700 54538
rect 247040 15904 247092 15910
rect 247040 15846 247092 15852
rect 247052 3482 247080 15846
rect 248340 10334 248368 102054
rect 248892 99414 248920 102068
rect 249996 99414 250024 102068
rect 248880 99408 248932 99414
rect 248880 99350 248932 99356
rect 249708 99408 249760 99414
rect 249708 99350 249760 99356
rect 249984 99408 250036 99414
rect 249984 99350 250036 99356
rect 250996 99408 251048 99414
rect 250996 99350 251048 99356
rect 248420 46232 248472 46238
rect 248420 46174 248472 46180
rect 248328 10328 248380 10334
rect 248328 10270 248380 10276
rect 248432 3482 248460 46174
rect 249720 32502 249748 99350
rect 251008 55894 251036 99350
rect 250996 55888 251048 55894
rect 250996 55830 251048 55836
rect 251100 36582 251128 102068
rect 252126 102054 252508 102082
rect 253230 102054 253888 102082
rect 251180 98660 251232 98666
rect 251180 98602 251232 98608
rect 249800 36576 249852 36582
rect 249800 36518 249852 36524
rect 251088 36576 251140 36582
rect 251088 36518 251140 36524
rect 249708 32496 249760 32502
rect 249708 32438 249760 32444
rect 249812 3482 249840 36518
rect 251192 3482 251220 98602
rect 252480 24138 252508 102054
rect 253860 57254 253888 102054
rect 254320 99414 254348 102068
rect 255424 99414 255452 102068
rect 254308 99408 254360 99414
rect 254308 99350 254360 99356
rect 255228 99408 255280 99414
rect 255228 99350 255280 99356
rect 255412 99408 255464 99414
rect 255412 99350 255464 99356
rect 253848 57248 253900 57254
rect 253848 57190 253900 57196
rect 252560 55956 252612 55962
rect 252560 55898 252612 55904
rect 252468 24132 252520 24138
rect 252468 24074 252520 24080
rect 252572 3534 252600 55898
rect 252652 35216 252704 35222
rect 252652 35158 252704 35164
rect 252560 3528 252612 3534
rect 245580 480 245608 3470
rect 245672 3454 246804 3482
rect 247052 3454 248000 3482
rect 248432 3454 249196 3482
rect 249812 3454 250392 3482
rect 251192 3454 251496 3482
rect 252560 3470 252612 3476
rect 246776 480 246804 3454
rect 247972 480 248000 3454
rect 249168 480 249196 3454
rect 250364 480 250392 3454
rect 251468 480 251496 3454
rect 252664 480 252692 35158
rect 253940 24200 253992 24206
rect 253940 24142 253992 24148
rect 253848 3528 253900 3534
rect 253848 3470 253900 3476
rect 253952 3482 253980 24142
rect 255240 13122 255268 99350
rect 256528 73914 256556 102068
rect 257646 102054 258028 102082
rect 258658 102054 259408 102082
rect 256608 99408 256660 99414
rect 256608 99350 256660 99356
rect 256516 73908 256568 73914
rect 256516 73850 256568 73856
rect 256620 22778 256648 99350
rect 256700 57316 256752 57322
rect 256700 57258 256752 57264
rect 255320 22772 255372 22778
rect 255320 22714 255372 22720
rect 256608 22772 256660 22778
rect 256608 22714 256660 22720
rect 255228 13116 255280 13122
rect 255228 13058 255280 13064
rect 255332 3482 255360 22714
rect 256712 3482 256740 57258
rect 258000 14482 258028 102054
rect 259380 35222 259408 102054
rect 259748 99414 259776 102068
rect 260852 99414 260880 102068
rect 261970 102054 262168 102082
rect 263074 102054 263548 102082
rect 264178 102054 264928 102082
rect 259736 99408 259788 99414
rect 259736 99350 259788 99356
rect 260748 99408 260800 99414
rect 260748 99350 260800 99356
rect 260840 99408 260892 99414
rect 260840 99350 260892 99356
rect 262036 99408 262088 99414
rect 262036 99350 262088 99356
rect 260760 75206 260788 99350
rect 260748 75200 260800 75206
rect 260748 75142 260800 75148
rect 260840 58676 260892 58682
rect 260840 58618 260892 58624
rect 259460 37936 259512 37942
rect 259460 37878 259512 37884
rect 259368 35216 259420 35222
rect 259368 35158 259420 35164
rect 258080 19984 258132 19990
rect 258080 19926 258132 19932
rect 257988 14476 258040 14482
rect 257988 14418 258040 14424
rect 258092 3482 258120 19926
rect 259472 3482 259500 37878
rect 260852 3482 260880 58618
rect 262048 44878 262076 99350
rect 262036 44872 262088 44878
rect 262036 44814 262088 44820
rect 262140 37942 262168 102054
rect 263520 61402 263548 102054
rect 263600 61464 263652 61470
rect 263600 61406 263652 61412
rect 263508 61396 263560 61402
rect 263508 61338 263560 61344
rect 262220 50380 262272 50386
rect 262220 50322 262272 50328
rect 262128 37936 262180 37942
rect 262128 37878 262180 37884
rect 262232 3602 262260 50322
rect 262312 17264 262364 17270
rect 262312 17206 262364 17212
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 262324 3482 262352 17206
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 253860 480 253888 3470
rect 253952 3454 255084 3482
rect 255332 3454 256280 3482
rect 256712 3454 257476 3482
rect 258092 3454 258672 3482
rect 259472 3454 259868 3482
rect 260852 3454 261064 3482
rect 255056 480 255084 3454
rect 256252 480 256280 3454
rect 257448 480 257476 3454
rect 258644 480 258672 3454
rect 259840 480 259868 3454
rect 261036 480 261064 3454
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3538
rect 263612 3482 263640 61406
rect 264900 4826 264928 102054
rect 265176 99414 265204 102068
rect 265164 99408 265216 99414
rect 265164 99350 265216 99356
rect 266176 99408 266228 99414
rect 266176 99350 266228 99356
rect 266188 25566 266216 99350
rect 266176 25560 266228 25566
rect 266176 25502 266228 25508
rect 266280 21418 266308 102068
rect 267398 102054 267688 102082
rect 268502 102054 269068 102082
rect 266360 47592 266412 47598
rect 266360 47534 266412 47540
rect 266268 21412 266320 21418
rect 266268 21354 266320 21360
rect 265808 4888 265860 4894
rect 265808 4830 265860 4836
rect 264888 4820 264940 4826
rect 264888 4762 264940 4768
rect 263612 3454 264652 3482
rect 264624 480 264652 3454
rect 265820 480 265848 4830
rect 266372 3482 266400 47534
rect 267660 15910 267688 102054
rect 267740 68332 267792 68338
rect 267740 68274 267792 68280
rect 267648 15904 267700 15910
rect 267648 15846 267700 15852
rect 267752 3482 267780 68274
rect 269040 46238 269068 102054
rect 269592 99414 269620 102068
rect 269580 99408 269632 99414
rect 269580 99350 269632 99356
rect 270408 99408 270460 99414
rect 270408 99350 270460 99356
rect 270420 60042 270448 99350
rect 270604 98666 270632 102068
rect 270592 98660 270644 98666
rect 270592 98602 270644 98608
rect 270500 60104 270552 60110
rect 270500 60046 270552 60052
rect 270408 60036 270460 60042
rect 270408 59978 270460 59984
rect 269028 46232 269080 46238
rect 269028 46174 269080 46180
rect 269120 39364 269172 39370
rect 269120 39306 269172 39312
rect 269132 3482 269160 39306
rect 270512 3602 270540 60046
rect 271708 47598 271736 102068
rect 272826 102054 273208 102082
rect 273930 102054 274588 102082
rect 273180 68338 273208 102054
rect 273260 95940 273312 95946
rect 273260 95882 273312 95888
rect 273168 68332 273220 68338
rect 273168 68274 273220 68280
rect 271696 47592 271748 47598
rect 271696 47534 271748 47540
rect 270592 25628 270644 25634
rect 270592 25570 270644 25576
rect 270500 3596 270552 3602
rect 270500 3538 270552 3544
rect 270604 3482 270632 25570
rect 272892 6180 272944 6186
rect 272892 6122 272944 6128
rect 271696 3596 271748 3602
rect 271696 3538 271748 3544
rect 266372 3454 267044 3482
rect 267752 3454 268148 3482
rect 269132 3454 269344 3482
rect 267016 480 267044 3454
rect 268120 480 268148 3454
rect 269316 480 269344 3454
rect 270512 3454 270632 3482
rect 270512 480 270540 3454
rect 271708 480 271736 3538
rect 272904 480 272932 6122
rect 273272 3482 273300 95882
rect 274560 6186 274588 102054
rect 275020 99414 275048 102068
rect 276124 99414 276152 102068
rect 277150 102054 277348 102082
rect 278254 102054 278728 102082
rect 275008 99408 275060 99414
rect 275008 99350 275060 99356
rect 275928 99408 275980 99414
rect 275928 99350 275980 99356
rect 276112 99408 276164 99414
rect 276112 99350 276164 99356
rect 277216 99408 277268 99414
rect 277216 99350 277268 99356
rect 274640 62824 274692 62830
rect 274640 62766 274692 62772
rect 274548 6180 274600 6186
rect 274548 6122 274600 6128
rect 274652 3482 274680 62766
rect 275940 50386 275968 99350
rect 277228 62830 277256 99350
rect 277216 62824 277268 62830
rect 277216 62766 277268 62772
rect 275928 50380 275980 50386
rect 275928 50322 275980 50328
rect 277320 33794 277348 102054
rect 277308 33788 277360 33794
rect 277308 33730 277360 33736
rect 278700 26926 278728 102054
rect 279344 99414 279372 102068
rect 280448 99414 280476 102068
rect 279332 99408 279384 99414
rect 279332 99350 279384 99356
rect 280068 99408 280120 99414
rect 280068 99350 280120 99356
rect 280436 99408 280488 99414
rect 280436 99350 280488 99356
rect 281448 99408 281500 99414
rect 281448 99350 281500 99356
rect 280080 71126 280108 99350
rect 280068 71120 280120 71126
rect 280068 71062 280120 71068
rect 278780 71052 278832 71058
rect 278780 70994 278832 71000
rect 277400 26920 277452 26926
rect 277400 26862 277452 26868
rect 278688 26920 278740 26926
rect 278688 26862 278740 26868
rect 276020 18624 276072 18630
rect 276020 18566 276072 18572
rect 276032 3482 276060 18566
rect 277412 3482 277440 26862
rect 278792 3482 278820 70994
rect 280160 49020 280212 49026
rect 280160 48962 280212 48968
rect 278872 21480 278924 21486
rect 278872 21422 278924 21428
rect 278884 3602 278912 21422
rect 278872 3596 278924 3602
rect 278872 3538 278924 3544
rect 280068 3596 280120 3602
rect 280068 3538 280120 3544
rect 273272 3454 274128 3482
rect 274652 3454 275324 3482
rect 276032 3454 276520 3482
rect 277412 3454 277716 3482
rect 278792 3454 278912 3482
rect 274100 480 274128 3454
rect 275296 480 275324 3454
rect 276492 480 276520 3454
rect 277688 480 277716 3454
rect 278884 480 278912 3454
rect 280080 480 280108 3538
rect 280172 3482 280200 48962
rect 281460 17338 281488 99350
rect 281552 95946 281580 102068
rect 282670 102054 282868 102082
rect 283682 102054 284248 102082
rect 281540 95940 281592 95946
rect 281540 95882 281592 95888
rect 282840 64190 282868 102054
rect 281540 64184 281592 64190
rect 281540 64126 281592 64132
rect 282828 64184 282880 64190
rect 282828 64126 282880 64132
rect 281448 17332 281500 17338
rect 281448 17274 281500 17280
rect 281552 3482 281580 64126
rect 282920 42084 282972 42090
rect 282920 42026 282972 42032
rect 282932 3482 282960 42026
rect 284220 18630 284248 102054
rect 284772 99414 284800 102068
rect 285876 99414 285904 102068
rect 286980 100094 287008 102068
rect 288098 102054 288388 102082
rect 289202 102054 289768 102082
rect 286968 100088 287020 100094
rect 286968 100030 287020 100036
rect 287244 100020 287296 100026
rect 287244 99962 287296 99968
rect 284760 99408 284812 99414
rect 284760 99350 284812 99356
rect 285588 99408 285640 99414
rect 285588 99350 285640 99356
rect 285864 99408 285916 99414
rect 285864 99350 285916 99356
rect 286968 99408 287020 99414
rect 286968 99350 287020 99356
rect 285600 40730 285628 99350
rect 286980 69698 287008 99350
rect 285680 69692 285732 69698
rect 285680 69634 285732 69640
rect 286968 69692 287020 69698
rect 286968 69634 287020 69640
rect 284300 40724 284352 40730
rect 284300 40666 284352 40672
rect 285588 40724 285640 40730
rect 285588 40666 285640 40672
rect 284208 18624 284260 18630
rect 284208 18566 284260 18572
rect 284312 3482 284340 40666
rect 285692 3482 285720 69634
rect 287152 28280 287204 28286
rect 287152 28222 287204 28228
rect 287164 3534 287192 28222
rect 287152 3528 287204 3534
rect 280172 3454 281304 3482
rect 281552 3454 282500 3482
rect 282932 3454 283696 3482
rect 284312 3454 284800 3482
rect 285692 3454 285996 3482
rect 287152 3470 287204 3476
rect 281276 480 281304 3454
rect 282472 480 282500 3454
rect 283668 480 283696 3454
rect 284772 480 284800 3454
rect 285968 480 285996 3454
rect 287256 1442 287284 99962
rect 288360 28286 288388 102054
rect 289740 65550 289768 102054
rect 290200 99414 290228 102068
rect 291304 99414 291332 102068
rect 290188 99408 290240 99414
rect 290188 99350 290240 99356
rect 291108 99408 291160 99414
rect 291108 99350 291160 99356
rect 291292 99408 291344 99414
rect 291292 99350 291344 99356
rect 289820 97300 289872 97306
rect 289820 97242 289872 97248
rect 288440 65544 288492 65550
rect 288440 65486 288492 65492
rect 289728 65544 289780 65550
rect 289728 65486 289780 65492
rect 288348 28280 288400 28286
rect 288348 28222 288400 28228
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288452 3482 288480 65486
rect 289832 3482 289860 97242
rect 291120 39370 291148 99350
rect 292408 66910 292436 102068
rect 293526 102054 293908 102082
rect 294630 102054 295288 102082
rect 292488 99408 292540 99414
rect 292488 99350 292540 99356
rect 292396 66904 292448 66910
rect 292396 66846 292448 66852
rect 292500 49026 292528 99350
rect 292580 66972 292632 66978
rect 292580 66914 292632 66920
rect 292488 49020 292540 49026
rect 292488 48962 292540 48968
rect 291108 39364 291160 39370
rect 291108 39306 291160 39312
rect 291200 29640 291252 29646
rect 291200 29582 291252 29588
rect 291212 3482 291240 29582
rect 292592 3482 292620 66914
rect 293880 19990 293908 102054
rect 295260 42090 295288 102054
rect 295628 100230 295656 102068
rect 295616 100224 295668 100230
rect 295616 100166 295668 100172
rect 296628 100224 296680 100230
rect 296628 100166 296680 100172
rect 296640 76566 296668 100166
rect 296732 99618 296760 102068
rect 297744 102054 297850 102082
rect 298954 102054 299428 102082
rect 300058 102054 300808 102082
rect 296720 99612 296772 99618
rect 296720 99554 296772 99560
rect 297744 96665 297772 102054
rect 298008 99612 298060 99618
rect 298008 99554 298060 99560
rect 297730 96656 297786 96665
rect 297730 96591 297786 96600
rect 297914 96656 297970 96665
rect 297914 96591 297970 96600
rect 297928 89758 297956 96591
rect 297732 89752 297784 89758
rect 297732 89694 297784 89700
rect 297916 89752 297968 89758
rect 297916 89694 297968 89700
rect 297744 77246 297772 89694
rect 297732 77240 297784 77246
rect 297732 77182 297784 77188
rect 296628 76560 296680 76566
rect 296628 76502 296680 76508
rect 297824 67652 297876 67658
rect 297824 67594 297876 67600
rect 297836 60858 297864 67594
rect 297824 60852 297876 60858
rect 297824 60794 297876 60800
rect 297732 60716 297784 60722
rect 297732 60658 297784 60664
rect 297744 53106 297772 60658
rect 296720 53100 296772 53106
rect 296720 53042 296772 53048
rect 297732 53100 297784 53106
rect 297732 53042 297784 53048
rect 295248 42084 295300 42090
rect 295248 42026 295300 42032
rect 295340 31068 295392 31074
rect 295340 31010 295392 31016
rect 293868 19984 293920 19990
rect 293868 19926 293920 19932
rect 294328 7608 294380 7614
rect 294328 7550 294380 7556
rect 287164 1414 287284 1442
rect 287164 480 287192 1414
rect 288360 480 288388 3470
rect 288452 3454 289584 3482
rect 289832 3454 290780 3482
rect 291212 3454 291976 3482
rect 292592 3454 293172 3482
rect 289556 480 289584 3454
rect 290752 480 290780 3454
rect 291948 480 291976 3454
rect 293144 480 293172 3454
rect 294340 480 294368 7550
rect 295352 3482 295380 31010
rect 295352 3454 295564 3482
rect 295536 480 295564 3454
rect 296732 480 296760 53042
rect 296812 11756 296864 11762
rect 296812 11698 296864 11704
rect 296824 3482 296852 11698
rect 298020 7614 298048 99554
rect 299400 77994 299428 102054
rect 299388 77988 299440 77994
rect 299388 77930 299440 77936
rect 299480 54528 299532 54534
rect 299480 54470 299532 54476
rect 298100 51740 298152 51746
rect 298100 51682 298152 51688
rect 298008 7608 298060 7614
rect 298008 7550 298060 7556
rect 298112 3482 298140 51682
rect 299492 3482 299520 54470
rect 300780 11762 300808 102054
rect 301148 100230 301176 102068
rect 302068 102054 302174 102082
rect 303278 102054 303568 102082
rect 304382 102054 304948 102082
rect 301136 100224 301188 100230
rect 301136 100166 301188 100172
rect 302068 79422 302096 102054
rect 302148 100224 302200 100230
rect 302148 100166 302200 100172
rect 302056 79416 302108 79422
rect 302056 79358 302108 79364
rect 302160 32434 302188 100166
rect 302240 43444 302292 43450
rect 302240 43386 302292 43392
rect 302148 32428 302200 32434
rect 302148 32370 302200 32376
rect 300768 11756 300820 11762
rect 300768 11698 300820 11704
rect 301412 8968 301464 8974
rect 301412 8910 301464 8916
rect 296824 3454 297956 3482
rect 298112 3454 299152 3482
rect 299492 3454 300348 3482
rect 297928 480 297956 3454
rect 299124 480 299152 3454
rect 300320 480 300348 3454
rect 301424 480 301452 8910
rect 302252 3482 302280 43386
rect 303540 8974 303568 102054
rect 303620 72480 303672 72486
rect 303620 72422 303672 72428
rect 303528 8968 303580 8974
rect 303528 8910 303580 8916
rect 303632 3482 303660 72422
rect 304920 43450 304948 102054
rect 305472 99414 305500 102068
rect 306576 99414 306604 102068
rect 305460 99408 305512 99414
rect 305460 99350 305512 99356
rect 306288 99408 306340 99414
rect 306288 99350 306340 99356
rect 306564 99408 306616 99414
rect 306564 99350 306616 99356
rect 306300 57322 306328 99350
rect 306288 57316 306340 57322
rect 306288 57258 306340 57264
rect 307680 55894 307708 102068
rect 308706 102054 309088 102082
rect 309810 102054 310468 102082
rect 309060 72486 309088 102054
rect 309784 99408 309836 99414
rect 309784 99350 309836 99356
rect 309048 72480 309100 72486
rect 309048 72422 309100 72428
rect 306380 55888 306432 55894
rect 306380 55830 306432 55836
rect 307668 55888 307720 55894
rect 307668 55830 307720 55836
rect 304908 43444 304960 43450
rect 304908 43386 304960 43392
rect 305000 32496 305052 32502
rect 305000 32438 305052 32444
rect 305012 3534 305040 32438
rect 305092 10328 305144 10334
rect 305092 10270 305144 10276
rect 305000 3528 305052 3534
rect 302252 3454 302648 3482
rect 303632 3454 303844 3482
rect 305000 3470 305052 3476
rect 302620 480 302648 3454
rect 303816 480 303844 3454
rect 305104 1442 305132 10270
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 306392 3482 306420 55830
rect 307760 36576 307812 36582
rect 307760 36518 307812 36524
rect 307772 3482 307800 36518
rect 309140 24132 309192 24138
rect 309140 24074 309192 24080
rect 309152 3482 309180 24074
rect 309796 10402 309824 99350
rect 310440 29646 310468 102054
rect 310900 99414 310928 102068
rect 312004 99414 312032 102068
rect 313108 99498 313136 102068
rect 314226 102054 314608 102082
rect 313108 99470 313228 99498
rect 310888 99408 310940 99414
rect 310888 99350 310940 99356
rect 311808 99408 311860 99414
rect 311808 99350 311860 99356
rect 311992 99408 312044 99414
rect 311992 99350 312044 99356
rect 313096 99408 313148 99414
rect 313096 99350 313148 99356
rect 310520 57248 310572 57254
rect 310520 57190 310572 57196
rect 310428 29640 310480 29646
rect 310428 29582 310480 29588
rect 309784 10396 309836 10402
rect 309784 10338 309836 10344
rect 310532 3482 310560 57190
rect 311820 36582 311848 99350
rect 313108 73846 313136 99350
rect 313096 73840 313148 73846
rect 313096 73782 313148 73788
rect 311808 36576 311860 36582
rect 311808 36518 311860 36524
rect 313200 31074 313228 99470
rect 313280 73908 313332 73914
rect 313280 73850 313332 73856
rect 313188 31068 313240 31074
rect 313188 31010 313240 31016
rect 311900 13116 311952 13122
rect 311900 13058 311952 13064
rect 311912 3482 311940 13058
rect 313292 3534 313320 73850
rect 314580 58682 314608 102054
rect 315224 99414 315252 102068
rect 316328 99414 316356 102068
rect 315212 99408 315264 99414
rect 315212 99350 315264 99356
rect 315948 99408 316000 99414
rect 315948 99350 316000 99356
rect 316316 99408 316368 99414
rect 316316 99350 316368 99356
rect 317328 99408 317380 99414
rect 317328 99350 317380 99356
rect 315960 80782 315988 99350
rect 315948 80776 316000 80782
rect 315948 80718 316000 80724
rect 314568 58676 314620 58682
rect 314568 58618 314620 58624
rect 316040 35216 316092 35222
rect 316040 35158 316092 35164
rect 313372 22772 313424 22778
rect 313372 22714 313424 22720
rect 313280 3528 313332 3534
rect 305012 1414 305132 1442
rect 305012 480 305040 1414
rect 306208 480 306236 3470
rect 306392 3454 307432 3482
rect 307772 3454 308628 3482
rect 309152 3454 309824 3482
rect 310532 3454 311020 3482
rect 311912 3454 312216 3482
rect 313280 3470 313332 3476
rect 307404 480 307432 3454
rect 308600 480 308628 3454
rect 309796 480 309824 3454
rect 310992 480 311020 3454
rect 312188 480 312216 3454
rect 313384 480 313412 22714
rect 314660 14476 314712 14482
rect 314660 14418 314712 14424
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 314672 3482 314700 14418
rect 314580 480 314608 3470
rect 314672 3454 315804 3482
rect 315776 480 315804 3454
rect 316052 3346 316080 35158
rect 317340 13122 317368 99350
rect 317432 97306 317460 102068
rect 318550 102054 318748 102082
rect 319654 102054 320128 102082
rect 317420 97300 317472 97306
rect 317420 97242 317472 97248
rect 318720 75206 318748 102054
rect 317420 75200 317472 75206
rect 317420 75142 317472 75148
rect 318708 75200 318760 75206
rect 318708 75142 318760 75148
rect 317328 13116 317380 13122
rect 317328 13058 317380 13064
rect 317432 3346 317460 75142
rect 318800 44872 318852 44878
rect 318800 44814 318852 44820
rect 318812 3346 318840 44814
rect 320100 14550 320128 102054
rect 320652 99414 320680 102068
rect 321756 100706 321784 102068
rect 321744 100700 321796 100706
rect 321744 100642 321796 100648
rect 322756 100700 322808 100706
rect 322756 100642 322808 100648
rect 320640 99408 320692 99414
rect 320640 99350 320692 99356
rect 321468 99408 321520 99414
rect 321468 99350 321520 99356
rect 320180 37936 320232 37942
rect 320180 37878 320232 37884
rect 320088 14544 320140 14550
rect 320088 14486 320140 14492
rect 320192 3346 320220 37878
rect 321480 35222 321508 99350
rect 322768 83502 322796 100642
rect 322756 83496 322808 83502
rect 322756 83438 322808 83444
rect 321560 61396 321612 61402
rect 321560 61338 321612 61344
rect 321468 35216 321520 35222
rect 321468 35158 321520 35164
rect 321572 3482 321600 61338
rect 322860 21486 322888 102068
rect 323978 102054 324268 102082
rect 323584 100088 323636 100094
rect 323584 100030 323636 100036
rect 322940 25560 322992 25566
rect 322940 25502 322992 25508
rect 322848 21480 322900 21486
rect 322848 21422 322900 21428
rect 322848 4820 322900 4826
rect 322848 4762 322900 4768
rect 321572 3454 321692 3482
rect 316052 3318 317000 3346
rect 317432 3318 318104 3346
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 316972 480 317000 3318
rect 318076 480 318104 3318
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 3454
rect 322860 480 322888 4762
rect 322952 3346 322980 25502
rect 323596 4826 323624 100030
rect 324240 44878 324268 102054
rect 325068 100094 325096 102068
rect 326172 100570 326200 102068
rect 327184 100706 327212 102068
rect 327172 100700 327224 100706
rect 327172 100642 327224 100648
rect 326160 100564 326212 100570
rect 326160 100506 326212 100512
rect 326988 100564 327040 100570
rect 326988 100506 327040 100512
rect 325056 100088 325108 100094
rect 325056 100030 325108 100036
rect 324228 44872 324280 44878
rect 324228 44814 324280 44820
rect 324320 21412 324372 21418
rect 324320 21354 324372 21360
rect 323584 4820 323636 4826
rect 323584 4762 323636 4768
rect 324332 3346 324360 21354
rect 327000 15910 327028 100506
rect 328104 96665 328132 102190
rect 329104 100700 329156 100706
rect 329104 100642 329156 100648
rect 328090 96656 328146 96665
rect 328090 96591 328146 96600
rect 328366 96656 328422 96665
rect 328366 96591 328422 96600
rect 328380 82142 328408 96591
rect 328368 82136 328420 82142
rect 328368 82078 328420 82084
rect 328460 60036 328512 60042
rect 328460 59978 328512 59984
rect 327080 46232 327132 46238
rect 327080 46174 327132 46180
rect 325700 15904 325752 15910
rect 325700 15846 325752 15852
rect 326988 15904 327040 15910
rect 326988 15846 327040 15852
rect 325712 3482 325740 15846
rect 327092 3482 327120 46174
rect 328472 3482 328500 59978
rect 329116 46238 329144 100642
rect 329392 100026 329420 102068
rect 330510 102054 331168 102082
rect 329380 100020 329432 100026
rect 329380 99962 329432 99968
rect 329840 98660 329892 98666
rect 329840 98602 329892 98608
rect 329104 46232 329156 46238
rect 329104 46174 329156 46180
rect 329852 3482 329880 98602
rect 331140 37942 331168 102054
rect 331600 100706 331628 102068
rect 331588 100700 331640 100706
rect 331588 100642 331640 100648
rect 332508 100700 332560 100706
rect 332508 100642 332560 100648
rect 332520 68338 332548 100642
rect 332704 99754 332732 102068
rect 333624 102054 333730 102082
rect 334834 102054 335308 102082
rect 335938 102054 336688 102082
rect 332692 99748 332744 99754
rect 332692 99690 332744 99696
rect 333624 96665 333652 102054
rect 333888 99748 333940 99754
rect 333888 99690 333940 99696
rect 333610 96656 333666 96665
rect 333610 96591 333666 96600
rect 333794 96656 333850 96665
rect 333794 96591 333850 96600
rect 331220 68332 331272 68338
rect 331220 68274 331272 68280
rect 332508 68332 332560 68338
rect 332508 68274 332560 68280
rect 331128 37936 331180 37942
rect 331128 37878 331180 37884
rect 331232 3602 331260 68274
rect 333808 67538 333836 96591
rect 333716 67510 333836 67538
rect 333716 58002 333744 67510
rect 333704 57996 333756 58002
rect 333704 57938 333756 57944
rect 333796 57996 333848 58002
rect 333796 57938 333848 57944
rect 333808 48210 333836 57938
rect 333796 48204 333848 48210
rect 333796 48146 333848 48152
rect 331312 47592 331364 47598
rect 331312 47534 331364 47540
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 331324 3482 331352 47534
rect 333900 22778 333928 99690
rect 335280 71058 335308 102054
rect 335268 71052 335320 71058
rect 335268 70994 335320 71000
rect 335360 62824 335412 62830
rect 335360 62766 335412 62772
rect 333980 50380 334032 50386
rect 333980 50322 334032 50328
rect 333888 22772 333940 22778
rect 333888 22714 333940 22720
rect 333612 6180 333664 6186
rect 333612 6122 333664 6128
rect 332416 3596 332468 3602
rect 332416 3538 332468 3544
rect 325712 3454 326476 3482
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 329852 3454 330064 3482
rect 322952 3318 324084 3346
rect 324332 3318 325280 3346
rect 324056 480 324084 3318
rect 325252 480 325280 3318
rect 326448 480 326476 3454
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330036 480 330064 3454
rect 331232 3454 331352 3482
rect 331232 480 331260 3454
rect 332428 480 332456 3538
rect 333624 480 333652 6122
rect 333992 3482 334020 50322
rect 335372 3482 335400 62766
rect 336660 6186 336688 102054
rect 337028 100706 337056 102068
rect 338132 100706 338160 102068
rect 339250 102054 339448 102082
rect 340262 102054 340828 102082
rect 337016 100700 337068 100706
rect 337016 100642 337068 100648
rect 338028 100700 338080 100706
rect 338028 100642 338080 100648
rect 338120 100700 338172 100706
rect 338120 100642 338172 100648
rect 339316 100700 339368 100706
rect 339316 100642 339368 100648
rect 337384 100088 337436 100094
rect 337384 100030 337436 100036
rect 337396 33794 337424 100030
rect 338040 50386 338068 100642
rect 339328 84862 339356 100642
rect 339316 84856 339368 84862
rect 339316 84798 339368 84804
rect 338028 50380 338080 50386
rect 338028 50322 338080 50328
rect 336740 33788 336792 33794
rect 336740 33730 336792 33736
rect 337384 33788 337436 33794
rect 337384 33730 337436 33736
rect 336648 6180 336700 6186
rect 336648 6122 336700 6128
rect 336752 3482 336780 33730
rect 338120 26920 338172 26926
rect 338120 26862 338172 26868
rect 338132 3482 338160 26862
rect 339420 17270 339448 102054
rect 339500 71120 339552 71126
rect 339500 71062 339552 71068
rect 339408 17264 339460 17270
rect 339408 17206 339460 17212
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339512 480 339540 71062
rect 340800 51746 340828 102054
rect 341352 99414 341380 102068
rect 341340 99408 341392 99414
rect 341340 99350 341392 99356
rect 342168 99408 342220 99414
rect 342168 99350 342220 99356
rect 340880 95940 340932 95946
rect 340880 95882 340932 95888
rect 340788 51740 340840 51746
rect 340788 51682 340840 51688
rect 339592 17332 339644 17338
rect 339592 17274 339644 17280
rect 339604 3482 339632 17274
rect 340892 3482 340920 95882
rect 342180 86290 342208 99350
rect 342456 98666 342484 102068
rect 343560 99414 343588 102068
rect 344678 102054 344968 102082
rect 345690 102054 346348 102082
rect 343548 99408 343600 99414
rect 343548 99350 343600 99356
rect 342444 98660 342496 98666
rect 342444 98602 342496 98608
rect 342168 86284 342220 86290
rect 342168 86226 342220 86232
rect 342260 64184 342312 64190
rect 342260 64126 342312 64132
rect 342272 3482 342300 64126
rect 343640 18624 343692 18630
rect 343640 18566 343692 18572
rect 343652 3482 343680 18566
rect 344940 10334 344968 102054
rect 345664 99408 345716 99414
rect 345664 99350 345716 99356
rect 345676 40798 345704 99350
rect 345664 40792 345716 40798
rect 345664 40734 345716 40740
rect 345020 40724 345072 40730
rect 345020 40666 345072 40672
rect 344928 10328 344980 10334
rect 344928 10270 344980 10276
rect 345032 3482 345060 40666
rect 346320 18630 346348 102054
rect 346780 99414 346808 102068
rect 347884 99414 347912 102068
rect 348988 99498 349016 102068
rect 350106 102054 350488 102082
rect 351210 102054 351868 102082
rect 348988 99470 349108 99498
rect 346768 99408 346820 99414
rect 346768 99350 346820 99356
rect 347688 99408 347740 99414
rect 347688 99350 347740 99356
rect 347872 99408 347924 99414
rect 347872 99350 347924 99356
rect 348976 99408 349028 99414
rect 348976 99350 349028 99356
rect 346400 69692 346452 69698
rect 346400 69634 346452 69640
rect 346308 18624 346360 18630
rect 346308 18566 346360 18572
rect 346412 3482 346440 69634
rect 347700 61402 347728 99350
rect 347688 61396 347740 61402
rect 347688 61338 347740 61344
rect 348988 42158 349016 99350
rect 348976 42152 349028 42158
rect 348976 42094 349028 42100
rect 347780 28280 347832 28286
rect 347780 28222 347832 28228
rect 347792 3534 347820 28222
rect 349080 24138 349108 99470
rect 349160 65544 349212 65550
rect 349160 65486 349212 65492
rect 349068 24132 349120 24138
rect 349068 24074 349120 24080
rect 347872 4820 347924 4826
rect 347872 4762 347924 4768
rect 347780 3528 347832 3534
rect 339604 3454 340736 3482
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 343652 3454 344324 3482
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 347780 3470 347832 3476
rect 340708 480 340736 3454
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 3454
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 4762
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 349172 3482 349200 65486
rect 350460 54602 350488 102054
rect 351840 87650 351868 102054
rect 352208 99414 352236 102068
rect 353312 100094 353340 102068
rect 354430 102054 354628 102082
rect 355534 102054 356008 102082
rect 353300 100088 353352 100094
rect 353300 100030 353352 100036
rect 352196 99408 352248 99414
rect 352196 99350 352248 99356
rect 353208 99408 353260 99414
rect 353208 99350 353260 99356
rect 351828 87644 351880 87650
rect 351828 87586 351880 87592
rect 350448 54596 350500 54602
rect 350448 54538 350500 54544
rect 351920 49020 351972 49026
rect 351920 48962 351972 48968
rect 350540 39364 350592 39370
rect 350540 39306 350592 39312
rect 350552 12442 350580 39306
rect 351932 12442 351960 48962
rect 350540 12436 350592 12442
rect 350540 12378 350592 12384
rect 351368 12436 351420 12442
rect 351368 12378 351420 12384
rect 351920 12436 351972 12442
rect 351920 12378 351972 12384
rect 352564 12436 352616 12442
rect 352564 12378 352616 12384
rect 349080 480 349108 3470
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 12378
rect 352576 480 352604 12378
rect 353220 4894 353248 99350
rect 354600 91798 354628 102054
rect 354588 91792 354640 91798
rect 354588 91734 354640 91740
rect 353392 66904 353444 66910
rect 353392 66846 353444 66852
rect 353404 58018 353432 66846
rect 353312 57990 353432 58018
rect 353312 57934 353340 57990
rect 353300 57928 353352 57934
rect 353300 57870 353352 57876
rect 353300 48340 353352 48346
rect 353300 48282 353352 48288
rect 353312 38842 353340 48282
rect 353312 38814 353432 38842
rect 353404 38706 353432 38814
rect 353312 38678 353432 38706
rect 353312 38622 353340 38678
rect 353300 38616 353352 38622
rect 353300 38558 353352 38564
rect 353392 38616 353444 38622
rect 353392 38558 353444 38564
rect 353404 29050 353432 38558
rect 353312 29022 353432 29050
rect 353312 27606 353340 29022
rect 353300 27600 353352 27606
rect 353300 27542 353352 27548
rect 353852 27600 353904 27606
rect 353852 27542 353904 27548
rect 353864 12322 353892 27542
rect 355980 19990 356008 102054
rect 356624 99414 356652 102068
rect 357728 99414 357756 102068
rect 356612 99408 356664 99414
rect 356612 99350 356664 99356
rect 357348 99408 357400 99414
rect 357348 99350 357400 99356
rect 357716 99408 357768 99414
rect 357716 99350 357768 99356
rect 358636 99408 358688 99414
rect 358636 99350 358688 99356
rect 356060 76560 356112 76566
rect 356060 76502 356112 76508
rect 354680 19984 354732 19990
rect 354680 19926 354732 19932
rect 355968 19984 356020 19990
rect 355968 19926 356020 19932
rect 354692 12510 354720 19926
rect 354680 12504 354732 12510
rect 354680 12446 354732 12452
rect 353772 12294 353892 12322
rect 354956 12368 355008 12374
rect 354956 12310 355008 12316
rect 353772 9654 353800 12294
rect 354968 9654 354996 12310
rect 353760 9648 353812 9654
rect 353760 9590 353812 9596
rect 354956 9648 355008 9654
rect 354956 9590 355008 9596
rect 353760 9512 353812 9518
rect 353760 9454 353812 9460
rect 354956 9512 355008 9518
rect 354956 9454 355008 9460
rect 353208 4888 353260 4894
rect 353208 4830 353260 4836
rect 353772 480 353800 9454
rect 354968 480 354996 9454
rect 356072 7614 356100 76502
rect 357360 49026 357388 99350
rect 358648 76566 358676 99350
rect 358636 76560 358688 76566
rect 358636 76502 358688 76508
rect 357348 49020 357400 49026
rect 357348 48962 357400 48968
rect 356152 42084 356204 42090
rect 356152 42026 356204 42032
rect 356060 7608 356112 7614
rect 356060 7550 356112 7556
rect 356164 480 356192 42026
rect 358740 7682 358768 102068
rect 359858 102054 360148 102082
rect 360962 102054 361528 102082
rect 360120 53106 360148 102054
rect 361500 77994 361528 102054
rect 362052 99414 362080 102068
rect 362224 100088 362276 100094
rect 362224 100030 362276 100036
rect 362040 99408 362092 99414
rect 362040 99350 362092 99356
rect 360200 77988 360252 77994
rect 360200 77930 360252 77936
rect 361488 77988 361540 77994
rect 361488 77930 361540 77936
rect 358820 53100 358872 53106
rect 358820 53042 358872 53048
rect 360108 53100 360160 53106
rect 360108 53042 360160 53048
rect 358832 12442 358860 53042
rect 358820 12436 358872 12442
rect 358820 12378 358872 12384
rect 359740 12436 359792 12442
rect 359740 12378 359792 12384
rect 358728 7676 358780 7682
rect 358728 7618 358780 7624
rect 357348 7608 357400 7614
rect 357348 7550 357400 7556
rect 357360 480 357388 7550
rect 358544 7540 358596 7546
rect 358544 7482 358596 7488
rect 358556 480 358584 7482
rect 359752 480 359780 12378
rect 360212 3482 360240 77930
rect 362236 11762 362264 100030
rect 363156 99414 363184 102068
rect 362868 99408 362920 99414
rect 362868 99350 362920 99356
rect 363144 99408 363196 99414
rect 363144 99350 363196 99356
rect 364156 99408 364208 99414
rect 364156 99350 364208 99356
rect 362880 25566 362908 99350
rect 364168 90370 364196 99350
rect 364156 90364 364208 90370
rect 364156 90306 364208 90312
rect 364260 79354 364288 102068
rect 365286 102054 365668 102082
rect 366390 102054 367048 102082
rect 364340 79416 364392 79422
rect 364340 79358 364392 79364
rect 364248 79348 364300 79354
rect 364248 79290 364300 79296
rect 362960 32428 363012 32434
rect 362960 32370 363012 32376
rect 362868 25560 362920 25566
rect 362868 25502 362920 25508
rect 361580 11756 361632 11762
rect 361580 11698 361632 11704
rect 362224 11756 362276 11762
rect 362224 11698 362276 11704
rect 361592 3482 361620 11698
rect 362972 3482 363000 32370
rect 360212 3454 360976 3482
rect 361592 3454 362172 3482
rect 362972 3454 363368 3482
rect 360948 480 360976 3454
rect 362144 480 362172 3454
rect 363340 480 363368 3454
rect 364352 3346 364380 79358
rect 365640 39370 365668 102054
rect 367020 57254 367048 102054
rect 367480 99414 367508 102068
rect 368584 99414 368612 102068
rect 367468 99408 367520 99414
rect 367468 99350 367520 99356
rect 368388 99408 368440 99414
rect 368388 99350 368440 99356
rect 368572 99408 368624 99414
rect 368572 99350 368624 99356
rect 368400 93158 368428 99350
rect 368388 93152 368440 93158
rect 368388 93094 368440 93100
rect 369688 60042 369716 102068
rect 369768 99408 369820 99414
rect 369768 99350 369820 99356
rect 369676 60036 369728 60042
rect 369676 59978 369728 59984
rect 367100 57316 367152 57322
rect 367100 57258 367152 57264
rect 367008 57248 367060 57254
rect 367008 57190 367060 57196
rect 365720 43444 365772 43450
rect 365720 43386 365772 43392
rect 365628 39364 365680 39370
rect 365628 39306 365680 39312
rect 365732 3602 365760 43386
rect 365812 8968 365864 8974
rect 365812 8910 365864 8916
rect 365720 3596 365772 3602
rect 365720 3538 365772 3544
rect 365824 3482 365852 8910
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 365732 3454 365852 3482
rect 364352 3318 364564 3346
rect 364536 480 364564 3318
rect 365732 480 365760 3454
rect 366928 480 366956 3538
rect 367112 3346 367140 57258
rect 368480 10396 368532 10402
rect 368480 10338 368532 10344
rect 368492 3346 368520 10338
rect 369780 8974 369808 99350
rect 370792 95946 370820 102068
rect 371818 102054 372568 102082
rect 370780 95940 370832 95946
rect 370780 95882 370832 95888
rect 371240 72480 371292 72486
rect 371240 72422 371292 72428
rect 371252 66230 371280 72422
rect 371240 66224 371292 66230
rect 371240 66166 371292 66172
rect 371240 56636 371292 56642
rect 371240 56578 371292 56584
rect 369860 55888 369912 55894
rect 369860 55830 369912 55836
rect 369872 19310 369900 55830
rect 371252 46918 371280 56578
rect 371240 46912 371292 46918
rect 371240 46854 371292 46860
rect 371240 37324 371292 37330
rect 371240 37266 371292 37272
rect 371252 27606 371280 37266
rect 371240 27600 371292 27606
rect 371240 27542 371292 27548
rect 372540 26926 372568 102054
rect 372908 99414 372936 102068
rect 374012 99414 374040 102068
rect 375130 102054 375328 102082
rect 376234 102054 376708 102082
rect 372896 99408 372948 99414
rect 372896 99350 372948 99356
rect 373908 99408 373960 99414
rect 373908 99350 373960 99356
rect 374000 99408 374052 99414
rect 374000 99350 374052 99356
rect 375196 99408 375248 99414
rect 375196 99350 375248 99356
rect 373920 55894 373948 99350
rect 375208 80714 375236 99350
rect 375196 80708 375248 80714
rect 375196 80650 375248 80656
rect 374000 73840 374052 73846
rect 374000 73782 374052 73788
rect 373908 55888 373960 55894
rect 373908 55830 373960 55836
rect 372620 29640 372672 29646
rect 372620 29582 372672 29588
rect 372528 26920 372580 26926
rect 372528 26862 372580 26868
rect 369860 19304 369912 19310
rect 369860 19246 369912 19252
rect 371240 18012 371292 18018
rect 371240 17954 371292 17960
rect 371252 12510 371280 17954
rect 372632 12510 372660 29582
rect 371240 12504 371292 12510
rect 371240 12446 371292 12452
rect 372620 12504 372672 12510
rect 372620 12446 372672 12452
rect 371608 12368 371660 12374
rect 371608 12310 371660 12316
rect 372804 12368 372856 12374
rect 372804 12310 372856 12316
rect 370412 9716 370464 9722
rect 370412 9658 370464 9664
rect 369768 8968 369820 8974
rect 369768 8910 369820 8916
rect 367112 3318 368060 3346
rect 368492 3318 369256 3346
rect 368032 480 368060 3318
rect 369228 480 369256 3318
rect 370424 480 370452 9658
rect 371620 480 371648 12310
rect 372816 480 372844 12310
rect 374012 7614 374040 73782
rect 374092 36576 374144 36582
rect 374092 36518 374144 36524
rect 374000 7608 374052 7614
rect 374000 7550 374052 7556
rect 374104 1442 374132 36518
rect 375300 28286 375328 102054
rect 376680 62830 376708 102054
rect 377232 99414 377260 102068
rect 378336 99414 378364 102068
rect 377220 99408 377272 99414
rect 377220 99350 377272 99356
rect 378048 99408 378100 99414
rect 378048 99350 378100 99356
rect 378324 99408 378376 99414
rect 378324 99350 378376 99356
rect 376668 62824 376720 62830
rect 376668 62766 376720 62772
rect 376760 58676 376812 58682
rect 376760 58618 376812 58624
rect 375380 31068 375432 31074
rect 375380 31010 375432 31016
rect 375288 28280 375340 28286
rect 375288 28222 375340 28228
rect 375392 12442 375420 31010
rect 376772 12442 376800 58618
rect 375380 12436 375432 12442
rect 375380 12378 375432 12384
rect 376392 12436 376444 12442
rect 376392 12378 376444 12384
rect 376760 12436 376812 12442
rect 376760 12378 376812 12384
rect 377588 12436 377640 12442
rect 377588 12378 377640 12384
rect 375196 7608 375248 7614
rect 375196 7550 375248 7556
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 7550
rect 376404 480 376432 12378
rect 377600 480 377628 12378
rect 378060 4078 378088 99350
rect 378232 80776 378284 80782
rect 378232 80718 378284 80724
rect 378244 77330 378272 80718
rect 378152 77302 378272 77330
rect 378152 77246 378180 77302
rect 378140 77240 378192 77246
rect 378140 77182 378192 77188
rect 378140 67720 378192 67726
rect 378140 67662 378192 67668
rect 378152 67590 378180 67662
rect 378140 67584 378192 67590
rect 378140 67526 378192 67532
rect 379440 58682 379468 102068
rect 380558 102054 380848 102082
rect 381662 102054 382228 102082
rect 380164 99408 380216 99414
rect 380164 99350 380216 99356
rect 379428 58676 379480 58682
rect 379428 58618 379480 58624
rect 378140 57996 378192 58002
rect 378140 57938 378192 57944
rect 378152 57866 378180 57938
rect 378140 57860 378192 57866
rect 378140 57802 378192 57808
rect 378140 48340 378192 48346
rect 378140 48282 378192 48288
rect 378152 38842 378180 48282
rect 378152 38814 378272 38842
rect 378244 38706 378272 38814
rect 378152 38678 378272 38706
rect 378152 38622 378180 38678
rect 378140 38616 378192 38622
rect 378140 38558 378192 38564
rect 380176 29646 380204 99350
rect 380164 29640 380216 29646
rect 380164 29582 380216 29588
rect 378140 29096 378192 29102
rect 378140 29038 378192 29044
rect 378152 28966 378180 29038
rect 378140 28960 378192 28966
rect 378140 28902 378192 28908
rect 378232 28960 378284 28966
rect 378232 28902 378284 28908
rect 378244 19394 378272 28902
rect 378152 19366 378272 19394
rect 378152 19310 378180 19366
rect 378140 19304 378192 19310
rect 378140 19246 378192 19252
rect 379520 13116 379572 13122
rect 379520 13058 379572 13064
rect 378784 9716 378836 9722
rect 378784 9658 378836 9664
rect 378048 4072 378100 4078
rect 378048 4014 378100 4020
rect 378796 480 378824 9658
rect 379532 3346 379560 13058
rect 380820 3806 380848 102054
rect 380900 97300 380952 97306
rect 380900 97242 380952 97248
rect 380808 3800 380860 3806
rect 380808 3742 380860 3748
rect 380912 3346 380940 97242
rect 382200 14482 382228 102054
rect 382752 99414 382780 102068
rect 383764 99414 383792 102068
rect 382740 99408 382792 99414
rect 382740 99350 382792 99356
rect 383568 99408 383620 99414
rect 383568 99350 383620 99356
rect 383752 99408 383804 99414
rect 383752 99350 383804 99356
rect 382280 75200 382332 75206
rect 382280 75142 382332 75148
rect 382188 14476 382240 14482
rect 382188 14418 382240 14424
rect 382292 3482 382320 75142
rect 383580 64190 383608 99350
rect 383568 64184 383620 64190
rect 383568 64126 383620 64132
rect 383660 35216 383712 35222
rect 383660 35158 383712 35164
rect 382372 14544 382424 14550
rect 382372 14486 382424 14492
rect 382384 3602 382412 14486
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 383568 3596 383620 3602
rect 383568 3538 383620 3544
rect 382292 3454 382412 3482
rect 379532 3318 380020 3346
rect 380912 3318 381216 3346
rect 379992 480 380020 3318
rect 381188 480 381216 3318
rect 382384 480 382412 3454
rect 383580 480 383608 3538
rect 383672 3346 383700 35158
rect 384868 21418 384896 102068
rect 385972 100094 386000 102068
rect 387090 102054 387748 102082
rect 385960 100088 386012 100094
rect 385960 100030 386012 100036
rect 384948 99408 385000 99414
rect 384948 99350 385000 99356
rect 384856 21412 384908 21418
rect 384856 21354 384908 21360
rect 384960 4146 384988 99350
rect 385040 83496 385092 83502
rect 385040 83438 385092 83444
rect 384948 4140 385000 4146
rect 384948 4082 385000 4088
rect 385052 3346 385080 83438
rect 386420 21480 386472 21486
rect 386420 21422 386472 21428
rect 386432 3346 386460 21422
rect 387720 3874 387748 102054
rect 388180 99414 388208 102068
rect 388168 99408 388220 99414
rect 388168 99350 388220 99356
rect 389088 99408 389140 99414
rect 389088 99350 389140 99356
rect 387800 44872 387852 44878
rect 387800 44814 387852 44820
rect 387708 3868 387760 3874
rect 387708 3810 387760 3816
rect 387812 3346 387840 44814
rect 389100 31074 389128 99350
rect 389284 94518 389312 102068
rect 390310 102054 390508 102082
rect 391414 102054 391888 102082
rect 389272 94512 389324 94518
rect 389272 94454 389324 94460
rect 389180 33788 389232 33794
rect 389180 33730 389232 33736
rect 389088 31068 389140 31074
rect 389088 31010 389140 31016
rect 389192 19310 389220 33730
rect 389180 19304 389232 19310
rect 389180 19246 389232 19252
rect 389364 19304 389416 19310
rect 389364 19246 389416 19252
rect 389376 9738 389404 19246
rect 389376 9710 389496 9738
rect 389468 9654 389496 9710
rect 389456 9648 389508 9654
rect 389456 9590 389508 9596
rect 389456 9512 389508 9518
rect 389456 9454 389508 9460
rect 383672 3318 384712 3346
rect 385052 3318 385908 3346
rect 386432 3318 387104 3346
rect 387812 3318 388300 3346
rect 384684 480 384712 3318
rect 385880 480 385908 3318
rect 387076 480 387104 3318
rect 388272 480 388300 3318
rect 389468 480 389496 9454
rect 390480 3942 390508 102054
rect 390560 46232 390612 46238
rect 390560 46174 390612 46180
rect 390572 7614 390600 46174
rect 391860 32434 391888 102054
rect 392504 100706 392532 102068
rect 392492 100700 392544 100706
rect 392492 100642 392544 100648
rect 393228 100700 393280 100706
rect 393228 100642 393280 100648
rect 391940 82136 391992 82142
rect 391940 82078 391992 82084
rect 391848 32428 391900 32434
rect 391848 32370 391900 32376
rect 390652 15904 390704 15910
rect 390652 15846 390704 15852
rect 390560 7608 390612 7614
rect 390560 7550 390612 7556
rect 390468 3936 390520 3942
rect 390468 3878 390520 3884
rect 390664 480 390692 15846
rect 391952 12442 391980 82078
rect 393240 65618 393268 100642
rect 393412 100020 393464 100026
rect 393412 99962 393464 99968
rect 393228 65612 393280 65618
rect 393228 65554 393280 65560
rect 393424 12442 393452 99962
rect 393608 99754 393636 102068
rect 393596 99748 393648 99754
rect 393596 99690 393648 99696
rect 394608 99748 394660 99754
rect 394608 99690 394660 99696
rect 391940 12436 391992 12442
rect 391940 12378 391992 12384
rect 393044 12436 393096 12442
rect 393044 12378 393096 12384
rect 393412 12436 393464 12442
rect 393412 12378 393464 12384
rect 394240 12436 394292 12442
rect 394240 12378 394292 12384
rect 391848 7608 391900 7614
rect 391848 7550 391900 7556
rect 391860 480 391888 7550
rect 393056 480 393084 12378
rect 394252 480 394280 12378
rect 394620 4010 394648 99690
rect 394712 99618 394740 102068
rect 396000 99736 396028 102190
rect 396842 102054 397408 102082
rect 395908 99708 396028 99736
rect 394700 99612 394752 99618
rect 394700 99554 394752 99560
rect 395908 96626 395936 99708
rect 395988 99612 396040 99618
rect 395988 99554 396040 99560
rect 395896 96620 395948 96626
rect 395896 96562 395948 96568
rect 395804 87032 395856 87038
rect 395804 86974 395856 86980
rect 395816 80170 395844 86974
rect 395804 80164 395856 80170
rect 395804 80106 395856 80112
rect 395804 80028 395856 80034
rect 395804 79970 395856 79976
rect 395816 66978 395844 79970
rect 395804 66972 395856 66978
rect 395804 66914 395856 66920
rect 394700 37936 394752 37942
rect 394700 37878 394752 37884
rect 394712 12510 394740 37878
rect 396000 33794 396028 99554
rect 396080 68332 396132 68338
rect 396080 68274 396132 68280
rect 395988 33788 396040 33794
rect 395988 33730 396040 33736
rect 394700 12504 394752 12510
rect 394700 12446 394752 12452
rect 396092 12442 396120 68274
rect 396080 12436 396132 12442
rect 396080 12378 396132 12384
rect 396632 12436 396684 12442
rect 396632 12378 396684 12384
rect 395436 12368 395488 12374
rect 395436 12310 395488 12316
rect 395448 9654 395476 12310
rect 395436 9648 395488 9654
rect 395436 9590 395488 9596
rect 395436 9512 395488 9518
rect 395436 9454 395488 9460
rect 394608 4004 394660 4010
rect 394608 3946 394660 3952
rect 395448 480 395476 9454
rect 396644 480 396672 12378
rect 397380 3738 397408 102054
rect 397932 100706 397960 102068
rect 397920 100700 397972 100706
rect 397920 100642 397972 100648
rect 398748 100700 398800 100706
rect 398748 100642 398800 100648
rect 398760 35222 398788 100642
rect 399036 99414 399064 102068
rect 399024 99408 399076 99414
rect 399024 99350 399076 99356
rect 400036 99408 400088 99414
rect 400036 99350 400088 99356
rect 400048 47598 400076 99350
rect 398840 47592 398892 47598
rect 398840 47534 398892 47540
rect 400036 47592 400088 47598
rect 400036 47534 400088 47540
rect 398748 35216 398800 35222
rect 398748 35158 398800 35164
rect 397552 22772 397604 22778
rect 397552 22714 397604 22720
rect 397564 19394 397592 22714
rect 397472 19366 397592 19394
rect 397472 19310 397500 19366
rect 397460 19304 397512 19310
rect 397460 19246 397512 19252
rect 397828 9716 397880 9722
rect 397828 9658 397880 9664
rect 397368 3732 397420 3738
rect 397368 3674 397420 3680
rect 397840 480 397868 9658
rect 398852 3346 398880 47534
rect 400140 3602 400168 102068
rect 401258 102054 401548 102082
rect 402270 102054 402928 102082
rect 400220 71052 400272 71058
rect 400220 70994 400272 71000
rect 400128 3596 400180 3602
rect 400128 3538 400180 3544
rect 398852 3318 399064 3346
rect 399036 480 399064 3318
rect 400232 480 400260 70994
rect 401520 36582 401548 102054
rect 402900 68338 402928 102054
rect 403360 99414 403388 102068
rect 404464 99414 404492 102068
rect 403348 99408 403400 99414
rect 403348 99350 403400 99356
rect 404268 99408 404320 99414
rect 404268 99350 404320 99356
rect 404452 99408 404504 99414
rect 404452 99350 404504 99356
rect 402980 84856 403032 84862
rect 402980 84798 403032 84804
rect 402888 68332 402940 68338
rect 402888 68274 402940 68280
rect 401600 50380 401652 50386
rect 401600 50322 401652 50328
rect 401508 36576 401560 36582
rect 401508 36518 401560 36524
rect 401324 6180 401376 6186
rect 401324 6122 401376 6128
rect 401336 480 401364 6122
rect 401612 3346 401640 50322
rect 402992 3482 403020 84798
rect 404280 3670 404308 99350
rect 405568 69698 405596 102068
rect 406686 102054 407068 102082
rect 407790 102054 408448 102082
rect 405648 99408 405700 99414
rect 405648 99350 405700 99356
rect 405556 69692 405608 69698
rect 405556 69634 405608 69640
rect 405660 37942 405688 99350
rect 405740 51740 405792 51746
rect 405740 51682 405792 51688
rect 405648 37936 405700 37942
rect 405648 37878 405700 37884
rect 404360 17264 404412 17270
rect 404360 17206 404412 17212
rect 404268 3664 404320 3670
rect 404268 3606 404320 3612
rect 404372 3482 404400 17206
rect 405752 3482 405780 51682
rect 402992 3454 403756 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 407040 3466 407068 102054
rect 407120 86284 407172 86290
rect 407120 86226 407172 86232
rect 407132 3482 407160 86226
rect 408420 40730 408448 102054
rect 408788 100706 408816 102068
rect 408776 100700 408828 100706
rect 408776 100642 408828 100648
rect 409788 100700 409840 100706
rect 409788 100642 409840 100648
rect 408500 98660 408552 98666
rect 408500 98602 408552 98608
rect 408408 40724 408460 40730
rect 408408 40666 408460 40672
rect 401612 3318 402560 3346
rect 402532 480 402560 3318
rect 403728 480 403756 3454
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407028 3460 407080 3466
rect 407132 3454 407344 3482
rect 407028 3402 407080 3408
rect 407316 480 407344 3454
rect 408512 480 408540 98602
rect 409800 71058 409828 100642
rect 409892 99822 409920 102068
rect 411180 99906 411208 102190
rect 412114 102054 412588 102082
rect 413218 102054 413968 102082
rect 411904 100088 411956 100094
rect 411904 100030 411956 100036
rect 411088 99878 411208 99906
rect 409880 99816 409932 99822
rect 409880 99758 409932 99764
rect 411088 87038 411116 99878
rect 411168 99816 411220 99822
rect 411168 99758 411220 99764
rect 410984 87032 411036 87038
rect 410984 86974 411036 86980
rect 411076 87032 411128 87038
rect 411076 86974 411128 86980
rect 410996 82142 411024 86974
rect 410984 82136 411036 82142
rect 410984 82078 411036 82084
rect 410984 77376 411036 77382
rect 410904 77324 410984 77330
rect 410904 77318 411036 77324
rect 410904 77302 411024 77318
rect 409788 71052 409840 71058
rect 409788 70994 409840 71000
rect 410904 70446 410932 77302
rect 410892 70440 410944 70446
rect 410892 70382 410944 70388
rect 410984 70304 411036 70310
rect 410984 70246 411036 70252
rect 410996 61470 411024 70246
rect 410708 61464 410760 61470
rect 410708 61406 410760 61412
rect 410984 61464 411036 61470
rect 410984 61406 411036 61412
rect 410720 56574 410748 61406
rect 410708 56568 410760 56574
rect 410708 56510 410760 56516
rect 410984 50992 411036 50998
rect 410984 50934 411036 50940
rect 410996 41585 411024 50934
rect 410982 41576 411038 41585
rect 410982 41511 411038 41520
rect 408592 40792 408644 40798
rect 408592 40734 408644 40740
rect 408604 19310 408632 40734
rect 410890 36000 410946 36009
rect 410890 35935 410946 35944
rect 410904 35902 410932 35935
rect 410892 35896 410944 35902
rect 410892 35838 410944 35844
rect 410984 26308 411036 26314
rect 410984 26250 411036 26256
rect 410996 22166 411024 26250
rect 410984 22160 411036 22166
rect 410984 22102 411036 22108
rect 408592 19304 408644 19310
rect 408592 19246 408644 19252
rect 409696 19304 409748 19310
rect 409696 19246 409748 19252
rect 409708 480 409736 19246
rect 410800 10328 410852 10334
rect 410800 10270 410852 10276
rect 410812 4162 410840 10270
rect 410892 8424 410944 8430
rect 410892 8366 410944 8372
rect 410904 8294 410932 8366
rect 410892 8288 410944 8294
rect 410892 8230 410944 8236
rect 410812 4134 410932 4162
rect 410904 480 410932 4134
rect 411180 3534 411208 99758
rect 411916 18630 411944 100030
rect 412560 42090 412588 102054
rect 413940 61402 413968 102054
rect 414308 100094 414336 102068
rect 414296 100088 414348 100094
rect 414296 100030 414348 100036
rect 412640 61396 412692 61402
rect 412640 61338 412692 61344
rect 413928 61396 413980 61402
rect 413928 61338 413980 61344
rect 412548 42084 412600 42090
rect 412548 42026 412600 42032
rect 411904 18624 411956 18630
rect 411904 18566 411956 18572
rect 412088 18556 412140 18562
rect 412088 18498 412140 18504
rect 411168 3528 411220 3534
rect 411168 3470 411220 3476
rect 412100 480 412128 18498
rect 412652 12442 412680 61338
rect 415320 43450 415348 102068
rect 416438 102054 416728 102082
rect 417542 102054 418108 102082
rect 416700 54534 416728 102054
rect 416780 87644 416832 87650
rect 416780 87586 416832 87592
rect 416688 54528 416740 54534
rect 416688 54470 416740 54476
rect 415308 43444 415360 43450
rect 415308 43386 415360 43392
rect 414020 42152 414072 42158
rect 414020 42094 414072 42100
rect 414032 19310 414060 42094
rect 415400 24132 415452 24138
rect 415400 24074 415452 24080
rect 415412 19310 415440 24074
rect 414020 19304 414072 19310
rect 414020 19246 414072 19252
rect 414480 19304 414532 19310
rect 414480 19246 414532 19252
rect 415400 19304 415452 19310
rect 415400 19246 415452 19252
rect 412640 12436 412692 12442
rect 412640 12378 412692 12384
rect 413284 12436 413336 12442
rect 413284 12378 413336 12384
rect 413296 480 413324 12378
rect 414492 480 414520 19246
rect 415676 9716 415728 9722
rect 415676 9658 415728 9664
rect 415688 480 415716 9658
rect 416792 7614 416820 87586
rect 416872 54596 416924 54602
rect 416872 54538 416924 54544
rect 416780 7608 416832 7614
rect 416780 7550 416832 7556
rect 416884 480 416912 54538
rect 417976 7608 418028 7614
rect 417976 7550 418028 7556
rect 417988 480 418016 7550
rect 418080 4826 418108 102054
rect 418632 100706 418660 102068
rect 418620 100700 418672 100706
rect 418620 100642 418672 100648
rect 419448 100700 419500 100706
rect 419448 100642 419500 100648
rect 419460 89010 419488 100642
rect 419736 99822 419764 102068
rect 419724 99816 419776 99822
rect 419724 99758 419776 99764
rect 420736 99816 420788 99822
rect 420736 99758 420788 99764
rect 419448 89004 419500 89010
rect 419448 88946 419500 88952
rect 420748 72486 420776 99758
rect 420736 72480 420788 72486
rect 420736 72422 420788 72428
rect 419540 11756 419592 11762
rect 419540 11698 419592 11704
rect 419172 4888 419224 4894
rect 419172 4830 419224 4836
rect 418068 4820 418120 4826
rect 418068 4762 418120 4768
rect 419184 480 419212 4830
rect 419552 3482 419580 11698
rect 420840 7614 420868 102068
rect 421866 102054 422248 102082
rect 422970 102054 423628 102082
rect 420920 91792 420972 91798
rect 420920 91734 420972 91740
rect 420828 7608 420880 7614
rect 420828 7550 420880 7556
rect 420932 3482 420960 91734
rect 422220 44878 422248 102054
rect 423600 73846 423628 102054
rect 424060 100706 424088 102068
rect 425164 100706 425192 102068
rect 424048 100700 424100 100706
rect 424048 100642 424100 100648
rect 424968 100700 425020 100706
rect 424968 100642 425020 100648
rect 425152 100700 425204 100706
rect 425152 100642 425204 100648
rect 423588 73840 423640 73846
rect 423588 73782 423640 73788
rect 423680 49020 423732 49026
rect 423680 48962 423732 48968
rect 422208 44872 422260 44878
rect 422208 44814 422260 44820
rect 422300 19984 422352 19990
rect 422300 19926 422352 19932
rect 422312 3482 422340 19926
rect 423692 3482 423720 48962
rect 424980 10334 425008 100642
rect 426452 98954 426480 102326
rect 477342 102190 477540 102218
rect 427294 102054 427768 102082
rect 427084 100700 427136 100706
rect 427084 100642 427136 100648
rect 426360 98926 426480 98954
rect 425060 76560 425112 76566
rect 425060 76502 425112 76508
rect 424968 10328 425020 10334
rect 424968 10270 425020 10276
rect 425072 3482 425100 76502
rect 426360 75206 426388 98926
rect 426348 75200 426400 75206
rect 426348 75142 426400 75148
rect 426440 53100 426492 53106
rect 426440 53042 426492 53048
rect 426348 7676 426400 7682
rect 426348 7618 426400 7624
rect 419552 3454 420408 3482
rect 420932 3454 421604 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 425072 3454 425192 3482
rect 420380 480 420408 3454
rect 421576 480 421604 3454
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425164 480 425192 3454
rect 426360 480 426388 7618
rect 426452 3482 426480 53042
rect 427096 49026 427124 100642
rect 427084 49020 427136 49026
rect 427084 48962 427136 48968
rect 427740 11830 427768 102054
rect 428384 99414 428412 102068
rect 429488 99414 429516 102068
rect 430592 100026 430620 102068
rect 431710 102054 431908 102082
rect 432814 102054 433288 102082
rect 430580 100020 430632 100026
rect 430580 99962 430632 99968
rect 428372 99408 428424 99414
rect 428372 99350 428424 99356
rect 429108 99408 429160 99414
rect 429108 99350 429160 99356
rect 429476 99408 429528 99414
rect 429476 99350 429528 99356
rect 430488 99408 430540 99414
rect 430488 99350 430540 99356
rect 427820 77988 427872 77994
rect 427820 77930 427872 77936
rect 427728 11824 427780 11830
rect 427728 11766 427780 11772
rect 427832 3482 427860 77930
rect 429120 46238 429148 99350
rect 430500 76566 430528 99350
rect 430580 90364 430632 90370
rect 430580 90306 430632 90312
rect 430488 76560 430540 76566
rect 430488 76502 430540 76508
rect 429108 46232 429160 46238
rect 429108 46174 429160 46180
rect 429200 25560 429252 25566
rect 429200 25502 429252 25508
rect 429212 3482 429240 25502
rect 430592 3482 430620 90306
rect 431880 50386 431908 102054
rect 433260 82142 433288 102054
rect 433812 99414 433840 102068
rect 434916 99414 434944 102068
rect 433800 99408 433852 99414
rect 433800 99350 433852 99356
rect 434628 99408 434680 99414
rect 434628 99350 434680 99356
rect 434904 99408 434956 99414
rect 434904 99350 434956 99356
rect 435916 99408 435968 99414
rect 435916 99350 435968 99356
rect 433248 82136 433300 82142
rect 433248 82078 433300 82084
rect 431960 79348 432012 79354
rect 431960 79290 432012 79296
rect 431868 50380 431920 50386
rect 431868 50322 431920 50328
rect 431972 3482 432000 79290
rect 433340 57248 433392 57254
rect 433340 57190 433392 57196
rect 426452 3454 427584 3482
rect 427832 3454 428780 3482
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 431972 3454 432368 3482
rect 427556 480 427584 3454
rect 428752 480 428780 3454
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3454
rect 433352 3398 433380 57190
rect 433432 39364 433484 39370
rect 433432 39306 433484 39312
rect 433444 3482 433472 39306
rect 434640 13122 434668 99350
rect 434720 93152 434772 93158
rect 434720 93094 434772 93100
rect 434628 13116 434680 13122
rect 434628 13058 434680 13064
rect 434732 3482 434760 93094
rect 435928 91798 435956 99350
rect 435916 91792 435968 91798
rect 435916 91734 435968 91740
rect 436020 57254 436048 102068
rect 437138 102054 437428 102082
rect 438242 102054 438808 102082
rect 436008 57248 436060 57254
rect 436008 57190 436060 57196
rect 437400 15910 437428 102054
rect 438124 100088 438176 100094
rect 438124 100030 438176 100036
rect 437480 60036 437532 60042
rect 437480 59978 437532 59984
rect 437388 15904 437440 15910
rect 437388 15846 437440 15852
rect 437020 8968 437072 8974
rect 437020 8910 437072 8916
rect 433444 3454 433564 3482
rect 434732 3454 435864 3482
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433536 480 433564 3454
rect 434628 3392 434680 3398
rect 434628 3334 434680 3340
rect 434640 480 434668 3334
rect 435836 480 435864 3454
rect 437032 480 437060 8910
rect 437492 3482 437520 59978
rect 438136 8974 438164 100030
rect 438780 39370 438808 102054
rect 439332 99414 439360 102068
rect 439320 99408 439372 99414
rect 439320 99350 439372 99356
rect 440148 99408 440200 99414
rect 440148 99350 440200 99356
rect 438860 95940 438912 95946
rect 438860 95882 438912 95888
rect 438768 39364 438820 39370
rect 438768 39306 438820 39312
rect 438124 8968 438176 8974
rect 438124 8910 438176 8916
rect 438872 3482 438900 95882
rect 440160 60042 440188 99350
rect 440344 98666 440372 102068
rect 440332 98660 440384 98666
rect 440332 98602 440384 98608
rect 441448 90370 441476 102068
rect 442566 102054 442948 102082
rect 441436 90364 441488 90370
rect 441436 90306 441488 90312
rect 440148 60036 440200 60042
rect 440148 59978 440200 59984
rect 442920 55894 442948 102054
rect 443656 97306 443684 102068
rect 444760 99414 444788 102068
rect 445864 99414 445892 102068
rect 444748 99408 444800 99414
rect 444748 99350 444800 99356
rect 445668 99408 445720 99414
rect 445668 99350 445720 99356
rect 445852 99408 445904 99414
rect 445852 99350 445904 99356
rect 443644 97300 443696 97306
rect 443644 97242 443696 97248
rect 443000 80708 443052 80714
rect 443000 80650 443052 80656
rect 441620 55888 441672 55894
rect 441620 55830 441672 55836
rect 442908 55888 442960 55894
rect 442908 55830 442960 55836
rect 440240 26920 440292 26926
rect 440240 26862 440292 26868
rect 440252 3482 440280 26862
rect 441632 3482 441660 55830
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 80650
rect 444380 62824 444432 62830
rect 444380 62766 444432 62772
rect 443092 28280 443144 28286
rect 443092 28222 443144 28228
rect 443104 3482 443132 28222
rect 444392 3482 444420 62766
rect 445680 26926 445708 99350
rect 446876 95946 446904 102068
rect 447994 102054 448468 102082
rect 449098 102054 449848 102082
rect 447048 99408 447100 99414
rect 447048 99350 447100 99356
rect 446864 95940 446916 95946
rect 446864 95882 446916 95888
rect 447060 62830 447088 99350
rect 447048 62824 447100 62830
rect 447048 62766 447100 62772
rect 447140 29640 447192 29646
rect 447140 29582 447192 29588
rect 445668 26920 445720 26926
rect 445668 26862 445720 26868
rect 446588 4072 446640 4078
rect 446588 4014 446640 4020
rect 443104 3454 444236 3482
rect 444392 3454 445432 3482
rect 444208 480 444236 3454
rect 445404 480 445432 3454
rect 446600 480 446628 4014
rect 447152 3482 447180 29582
rect 448440 28286 448468 102054
rect 449820 58682 449848 102054
rect 450188 99414 450216 102068
rect 451292 99414 451320 102068
rect 452318 102054 452516 102082
rect 453422 102054 453988 102082
rect 450176 99408 450228 99414
rect 450176 99350 450228 99356
rect 451188 99408 451240 99414
rect 451188 99350 451240 99356
rect 451280 99408 451332 99414
rect 451280 99350 451332 99356
rect 448520 58676 448572 58682
rect 448520 58618 448572 58624
rect 449808 58676 449860 58682
rect 449808 58618 449860 58624
rect 448428 28280 448480 28286
rect 448428 28222 448480 28228
rect 448532 3482 448560 58618
rect 451200 17270 451228 99350
rect 452488 80714 452516 102054
rect 452568 99408 452620 99414
rect 452568 99350 452620 99356
rect 452476 80708 452528 80714
rect 452476 80650 452528 80656
rect 452580 64190 452608 99350
rect 451280 64184 451332 64190
rect 451280 64126 451332 64132
rect 452568 64184 452620 64190
rect 452568 64126 452620 64132
rect 451188 17264 451240 17270
rect 451188 17206 451240 17212
rect 450176 3800 450228 3806
rect 450176 3742 450228 3748
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 3742
rect 451292 3398 451320 64126
rect 453960 22778 453988 102054
rect 454512 99414 454540 102068
rect 455616 99414 455644 102068
rect 454500 99408 454552 99414
rect 454500 99350 454552 99356
rect 455328 99408 455380 99414
rect 455328 99350 455380 99356
rect 455604 99408 455656 99414
rect 455604 99350 455656 99356
rect 456616 99408 456668 99414
rect 456616 99350 456668 99356
rect 455340 51746 455368 99350
rect 456628 79354 456656 99350
rect 456616 79348 456668 79354
rect 456616 79290 456668 79296
rect 455328 51740 455380 51746
rect 455328 51682 455380 51688
rect 453948 22772 454000 22778
rect 453948 22714 454000 22720
rect 454040 21412 454092 21418
rect 454040 21354 454092 21360
rect 451372 14476 451424 14482
rect 451372 14418 451424 14424
rect 451280 3392 451332 3398
rect 451280 3334 451332 3340
rect 451384 1442 451412 14418
rect 453672 4140 453724 4146
rect 453672 4082 453724 4088
rect 452476 3392 452528 3398
rect 452476 3334 452528 3340
rect 451292 1414 451412 1442
rect 451292 480 451320 1414
rect 452488 480 452516 3334
rect 453684 480 453712 4082
rect 454052 3482 454080 21354
rect 456720 18630 456748 102068
rect 457838 102054 458128 102082
rect 458850 102054 459508 102082
rect 458100 53106 458128 102054
rect 459480 77994 459508 102054
rect 459940 100706 459968 102068
rect 461044 100706 461072 102068
rect 462056 102054 462162 102082
rect 463266 102054 463648 102082
rect 464370 102054 465028 102082
rect 459928 100700 459980 100706
rect 459928 100642 459980 100648
rect 460848 100700 460900 100706
rect 460848 100642 460900 100648
rect 461032 100700 461084 100706
rect 461032 100642 461084 100648
rect 459652 94512 459704 94518
rect 459652 94454 459704 94460
rect 459468 77988 459520 77994
rect 459468 77930 459520 77936
rect 458088 53100 458140 53106
rect 458088 53042 458140 53048
rect 458180 31068 458232 31074
rect 458180 31010 458232 31016
rect 455420 18624 455472 18630
rect 455420 18566 455472 18572
rect 456708 18624 456760 18630
rect 456708 18566 456760 18572
rect 455432 3482 455460 18566
rect 457260 3868 457312 3874
rect 457260 3810 457312 3816
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3810
rect 458192 3482 458220 31010
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 94454
rect 460860 14482 460888 100642
rect 462056 96665 462084 102054
rect 462964 100700 463016 100706
rect 462964 100642 463016 100648
rect 462042 96656 462098 96665
rect 462042 96591 462098 96600
rect 462226 96656 462282 96665
rect 462226 96591 462282 96600
rect 462240 89758 462268 96591
rect 462044 89752 462096 89758
rect 462228 89752 462280 89758
rect 462096 89700 462176 89706
rect 462044 89694 462176 89700
rect 462228 89694 462280 89700
rect 462056 89678 462176 89694
rect 462148 80170 462176 89678
rect 462976 86290 463004 100642
rect 462964 86284 463016 86290
rect 462964 86226 463016 86232
rect 462136 80164 462188 80170
rect 462136 80106 462188 80112
rect 462136 80028 462188 80034
rect 462136 79970 462188 79976
rect 462148 70394 462176 79970
rect 462056 70366 462176 70394
rect 462056 65550 462084 70366
rect 462320 65612 462372 65618
rect 462320 65554 462372 65560
rect 462044 65544 462096 65550
rect 462044 65486 462096 65492
rect 460940 32428 460992 32434
rect 460940 32370 460992 32376
rect 460848 14476 460900 14482
rect 460848 14418 460900 14424
rect 460848 3936 460900 3942
rect 460848 3878 460900 3884
rect 460860 480 460888 3878
rect 460952 3482 460980 32370
rect 462332 3482 462360 65554
rect 463620 19990 463648 102054
rect 465000 31074 465028 102054
rect 465368 99754 465396 102068
rect 465356 99748 465408 99754
rect 465356 99690 465408 99696
rect 466368 99748 466420 99754
rect 466368 99690 466420 99696
rect 466380 66910 466408 99690
rect 466472 99414 466500 102068
rect 466460 99408 466512 99414
rect 466460 99350 466512 99356
rect 467576 84862 467604 102068
rect 468694 102054 469168 102082
rect 467748 99408 467800 99414
rect 467748 99350 467800 99356
rect 467564 84856 467616 84862
rect 467564 84798 467616 84804
rect 466460 66972 466512 66978
rect 466460 66914 466512 66920
rect 466368 66904 466420 66910
rect 466368 66846 466420 66852
rect 465080 33788 465132 33794
rect 465080 33730 465132 33736
rect 464988 31068 465040 31074
rect 464988 31010 465040 31016
rect 463608 19984 463660 19990
rect 463608 19926 463660 19932
rect 464436 4004 464488 4010
rect 464436 3946 464488 3952
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3946
rect 465092 3482 465120 33730
rect 466472 3482 466500 66914
rect 467760 21418 467788 99350
rect 467932 35216 467984 35222
rect 467932 35158 467984 35164
rect 467748 21412 467800 21418
rect 467748 21354 467800 21360
rect 467840 3732 467892 3738
rect 467840 3674 467892 3680
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 3210 467880 3674
rect 467944 3398 467972 35158
rect 469140 3806 469168 102054
rect 469784 99414 469812 102068
rect 470888 99414 470916 102068
rect 469772 99408 469824 99414
rect 469772 99350 469824 99356
rect 470508 99408 470560 99414
rect 470508 99350 470560 99356
rect 470876 99408 470928 99414
rect 470876 99350 470928 99356
rect 471796 99408 471848 99414
rect 471796 99350 471848 99356
rect 469220 47592 469272 47598
rect 469220 47534 469272 47540
rect 469128 3800 469180 3806
rect 469128 3742 469180 3748
rect 469232 3482 469260 47534
rect 470520 24138 470548 99350
rect 471808 32434 471836 99350
rect 471796 32428 471848 32434
rect 471796 32370 471848 32376
rect 470508 24132 470560 24138
rect 470508 24074 470560 24080
rect 471900 4146 471928 102068
rect 473018 102054 473308 102082
rect 474122 102054 474688 102082
rect 473280 47598 473308 102054
rect 473360 68332 473412 68338
rect 473360 68274 473412 68280
rect 473268 47592 473320 47598
rect 473268 47534 473320 47540
rect 471980 36576 472032 36582
rect 471980 36518 472032 36524
rect 471888 4140 471940 4146
rect 471888 4082 471940 4088
rect 471520 3596 471572 3602
rect 471520 3538 471572 3544
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 3182 467972 3210
rect 467944 480 467972 3182
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3538
rect 471992 3346 472020 36518
rect 473372 3346 473400 68274
rect 474660 33794 474688 102054
rect 475212 99414 475240 102068
rect 476316 100706 476344 102068
rect 476304 100700 476356 100706
rect 476304 100642 476356 100648
rect 475200 99408 475252 99414
rect 475200 99350 475252 99356
rect 476028 99408 476080 99414
rect 476028 99350 476080 99356
rect 474648 33788 474700 33794
rect 474648 33730 474700 33736
rect 476040 4078 476068 99350
rect 477512 96642 477540 102190
rect 478446 102054 478828 102082
rect 479550 102054 480208 102082
rect 478236 100700 478288 100706
rect 478236 100642 478288 100648
rect 477420 96614 477540 96642
rect 477420 37942 477448 96614
rect 478248 94518 478276 100642
rect 478236 94512 478288 94518
rect 478236 94454 478288 94460
rect 477592 69692 477644 69698
rect 477592 69634 477644 69640
rect 476120 37936 476172 37942
rect 476120 37878 476172 37884
rect 477408 37936 477460 37942
rect 477408 37878 477460 37884
rect 476028 4072 476080 4078
rect 476028 4014 476080 4020
rect 475108 3664 475160 3670
rect 475108 3606 475160 3612
rect 471992 3318 472756 3346
rect 473372 3318 473952 3346
rect 472728 480 472756 3318
rect 473924 480 473952 3318
rect 475120 480 475148 3606
rect 476132 3346 476160 37878
rect 477604 3482 477632 69634
rect 478800 4010 478828 102054
rect 480180 93158 480208 102054
rect 480640 100706 480668 102068
rect 481744 100706 481772 102068
rect 480628 100700 480680 100706
rect 480628 100642 480680 100648
rect 481548 100700 481600 100706
rect 481548 100642 481600 100648
rect 481732 100700 481784 100706
rect 481732 100642 481784 100648
rect 480168 93152 480220 93158
rect 480168 93094 480220 93100
rect 480260 71052 480312 71058
rect 480260 70994 480312 71000
rect 478880 40724 478932 40730
rect 478880 40666 478932 40672
rect 478788 4004 478840 4010
rect 478788 3946 478840 3952
rect 477512 3454 477632 3482
rect 478696 3460 478748 3466
rect 476132 3318 476344 3346
rect 476316 480 476344 3318
rect 477512 480 477540 3454
rect 478696 3402 478748 3408
rect 478708 480 478736 3402
rect 478892 3346 478920 40666
rect 480272 3482 480300 70994
rect 481560 35222 481588 100642
rect 481548 35216 481600 35222
rect 481548 35158 481600 35164
rect 482848 25566 482876 102068
rect 483874 102054 484348 102082
rect 484978 102054 485728 102082
rect 482928 100700 482980 100706
rect 482928 100642 482980 100648
rect 482836 25560 482888 25566
rect 482836 25502 482888 25508
rect 482940 3942 482968 100642
rect 484320 36582 484348 102054
rect 484400 42084 484452 42090
rect 484400 42026 484452 42032
rect 484308 36576 484360 36582
rect 484308 36518 484360 36524
rect 483480 6180 483532 6186
rect 483480 6122 483532 6128
rect 482928 3936 482980 3942
rect 482928 3878 482980 3884
rect 482284 3528 482336 3534
rect 480272 3454 481128 3482
rect 482284 3470 482336 3476
rect 478892 3318 479932 3346
rect 479904 480 479932 3318
rect 481100 480 481128 3454
rect 482296 480 482324 3470
rect 483492 480 483520 6122
rect 484412 3482 484440 42026
rect 485700 3874 485728 102054
rect 486068 99414 486096 102068
rect 487172 99414 487200 102068
rect 488290 102054 488488 102082
rect 489394 102054 489868 102082
rect 486056 99408 486108 99414
rect 486056 99350 486108 99356
rect 487068 99408 487120 99414
rect 487068 99350 487120 99356
rect 487160 99408 487212 99414
rect 487160 99350 487212 99356
rect 488356 99408 488408 99414
rect 488356 99350 488408 99356
rect 485780 61396 485832 61402
rect 485780 61338 485832 61344
rect 485688 3868 485740 3874
rect 485688 3810 485740 3816
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 480 485820 61338
rect 487080 8974 487108 99350
rect 488368 43450 488396 99350
rect 487160 43444 487212 43450
rect 487160 43386 487212 43392
rect 488356 43444 488408 43450
rect 488356 43386 488408 43392
rect 486976 8968 487028 8974
rect 486976 8910 487028 8916
rect 487068 8968 487120 8974
rect 487068 8910 487120 8916
rect 486988 480 487016 8910
rect 487172 3482 487200 43386
rect 488460 3670 488488 102054
rect 488540 54528 488592 54534
rect 488540 54470 488592 54476
rect 488448 3664 488500 3670
rect 488448 3606 488500 3612
rect 488552 3482 488580 54470
rect 489840 6186 489868 102054
rect 490392 99414 490420 102068
rect 491496 99414 491524 102068
rect 492600 100094 492628 102068
rect 493718 102054 494008 102082
rect 494822 102054 495388 102082
rect 492588 100088 492640 100094
rect 492588 100030 492640 100036
rect 490380 99408 490432 99414
rect 490380 99350 490432 99356
rect 491208 99408 491260 99414
rect 491208 99350 491260 99356
rect 491484 99408 491536 99414
rect 491484 99350 491536 99356
rect 492588 99408 492640 99414
rect 492588 99350 492640 99356
rect 491220 83502 491248 99350
rect 491300 89004 491352 89010
rect 491300 88946 491352 88952
rect 491208 83496 491260 83502
rect 491208 83438 491260 83444
rect 489828 6180 489880 6186
rect 489828 6122 489880 6128
rect 490564 4820 490616 4826
rect 490564 4762 490616 4768
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 490576 480 490604 4762
rect 491312 3618 491340 88946
rect 492600 3738 492628 99350
rect 492680 72480 492732 72486
rect 492680 72422 492732 72428
rect 492588 3732 492640 3738
rect 492588 3674 492640 3680
rect 492692 3618 492720 72422
rect 493980 42090 494008 102054
rect 494060 44872 494112 44878
rect 494060 44814 494112 44820
rect 493968 42084 494020 42090
rect 493968 42026 494020 42032
rect 491312 3590 491800 3618
rect 492692 3590 492996 3618
rect 491772 480 491800 3590
rect 492968 480 492996 3590
rect 494072 3534 494100 44814
rect 494152 7608 494204 7614
rect 494152 7550 494204 7556
rect 494060 3528 494112 3534
rect 494060 3470 494112 3476
rect 494164 480 494192 7550
rect 495360 5250 495388 102054
rect 495912 99414 495940 102068
rect 496924 99414 496952 102068
rect 498028 99498 498056 102068
rect 499146 102054 499528 102082
rect 500250 102054 500908 102082
rect 498028 99470 498148 99498
rect 495900 99408 495952 99414
rect 495900 99350 495952 99356
rect 496728 99408 496780 99414
rect 496728 99350 496780 99356
rect 496912 99408 496964 99414
rect 496912 99350 496964 99356
rect 498016 99408 498068 99414
rect 498016 99350 498068 99356
rect 495440 73840 495492 73846
rect 495440 73782 495492 73788
rect 495452 58177 495480 73782
rect 495438 58168 495494 58177
rect 495438 58103 495494 58112
rect 495438 58032 495494 58041
rect 495438 57967 495494 57976
rect 495452 57934 495480 57967
rect 495440 57928 495492 57934
rect 495440 57870 495492 57876
rect 495440 48340 495492 48346
rect 495440 48282 495492 48288
rect 495452 38622 495480 48282
rect 495440 38616 495492 38622
rect 495440 38558 495492 38564
rect 495440 29028 495492 29034
rect 495440 28970 495492 28976
rect 495452 19310 495480 28970
rect 495440 19304 495492 19310
rect 495440 19246 495492 19252
rect 495624 19304 495676 19310
rect 495624 19246 495676 19252
rect 495636 9761 495664 19246
rect 495438 9752 495494 9761
rect 495438 9687 495494 9696
rect 495622 9752 495678 9761
rect 495622 9687 495678 9696
rect 495452 9654 495480 9687
rect 495440 9648 495492 9654
rect 495440 9590 495492 9596
rect 496740 7614 496768 99350
rect 498028 89010 498056 99350
rect 498016 89004 498068 89010
rect 498016 88946 498068 88952
rect 497740 10328 497792 10334
rect 497740 10270 497792 10276
rect 496728 7608 496780 7614
rect 496728 7550 496780 7556
rect 495268 5222 495388 5250
rect 495268 3602 495296 5222
rect 495256 3596 495308 3602
rect 495256 3538 495308 3544
rect 495348 3528 495400 3534
rect 495348 3470 495400 3476
rect 495360 480 495388 3470
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 10270
rect 498120 3466 498148 99470
rect 498200 49020 498252 49026
rect 498200 48962 498252 48968
rect 498108 3460 498160 3466
rect 498108 3402 498160 3408
rect 498212 2854 498240 48962
rect 499500 10334 499528 102054
rect 499580 75200 499632 75206
rect 499580 75142 499632 75148
rect 499592 67590 499620 75142
rect 499580 67584 499632 67590
rect 499580 67526 499632 67532
rect 499580 57996 499632 58002
rect 499580 57938 499632 57944
rect 499488 10328 499540 10334
rect 499488 10270 499540 10276
rect 499592 2854 499620 57938
rect 500880 11762 500908 102054
rect 501340 99414 501368 102068
rect 502984 100020 503036 100026
rect 502984 99962 503036 99968
rect 501328 99408 501380 99414
rect 501328 99350 501380 99356
rect 502248 99408 502300 99414
rect 502248 99350 502300 99356
rect 501236 11824 501288 11830
rect 501236 11766 501288 11772
rect 500868 11756 500920 11762
rect 500868 11698 500920 11704
rect 498200 2848 498252 2854
rect 498200 2790 498252 2796
rect 499580 2848 499632 2854
rect 499580 2790 499632 2796
rect 498936 2780 498988 2786
rect 498936 2722 498988 2728
rect 500132 2780 500184 2786
rect 500132 2722 500184 2728
rect 498948 480 498976 2722
rect 500144 480 500172 2722
rect 501248 480 501276 11766
rect 502260 3738 502288 99350
rect 502340 76560 502392 76566
rect 502340 76502 502392 76508
rect 502248 3732 502300 3738
rect 502248 3674 502300 3680
rect 502352 2106 502380 76502
rect 502432 46232 502484 46238
rect 502432 46174 502484 46180
rect 502340 2100 502392 2106
rect 502340 2042 502392 2048
rect 502444 480 502472 46174
rect 502996 5506 503024 99962
rect 504376 30326 504404 118487
rect 504468 41410 504496 129639
rect 504560 88330 504588 162959
rect 504638 151872 504694 151881
rect 504638 151807 504694 151816
rect 504548 88324 504600 88330
rect 504548 88266 504600 88272
rect 504652 77246 504680 151807
rect 504744 111790 504772 174111
rect 504836 124166 504864 185127
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 505006 140856 505062 140865
rect 505006 140791 505008 140800
rect 505060 140791 505062 140800
rect 527824 140820 527876 140826
rect 505008 140762 505060 140768
rect 527824 140762 527876 140768
rect 504824 124160 504876 124166
rect 504824 124102 504876 124108
rect 504732 111784 504784 111790
rect 504732 111726 504784 111732
rect 514760 98660 514812 98666
rect 514760 98602 514812 98608
rect 509240 91792 509292 91798
rect 509240 91734 509292 91740
rect 506480 82136 506532 82142
rect 506480 82078 506532 82084
rect 504640 77240 504692 77246
rect 504640 77182 504692 77188
rect 505100 50380 505152 50386
rect 505100 50322 505152 50328
rect 504456 41404 504508 41410
rect 504456 41346 504508 41352
rect 504364 30320 504416 30326
rect 504364 30262 504416 30268
rect 502984 5500 503036 5506
rect 502984 5442 503036 5448
rect 504824 5500 504876 5506
rect 504824 5442 504876 5448
rect 503628 2100 503680 2106
rect 503628 2042 503680 2048
rect 503640 480 503668 2042
rect 504836 480 504864 5442
rect 505112 3482 505140 50322
rect 506492 3482 506520 82078
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507872 3482 507900 13058
rect 509252 3482 509280 91734
rect 513380 60036 513432 60042
rect 513380 59978 513432 59984
rect 510620 57248 510672 57254
rect 510620 57190 510672 57196
rect 510632 3482 510660 57190
rect 512000 39364 512052 39370
rect 512000 39306 512052 39312
rect 505112 3454 506060 3482
rect 506492 3454 507256 3482
rect 507872 3454 508452 3482
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 506032 480 506060 3454
rect 507228 480 507256 3454
rect 508424 480 508452 3454
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 3398 512040 39306
rect 512092 15904 512144 15910
rect 512092 15846 512144 15852
rect 512000 3392 512052 3398
rect 512000 3334 512052 3340
rect 512104 1442 512132 15846
rect 513392 3482 513420 59978
rect 514772 3482 514800 98602
rect 518900 97300 518952 97306
rect 518900 97242 518952 97248
rect 516140 90364 516192 90370
rect 516140 90306 516192 90312
rect 516152 3482 516180 90306
rect 517520 55888 517572 55894
rect 517520 55830 517572 55836
rect 517532 3482 517560 55830
rect 518912 3482 518940 97242
rect 521660 95940 521712 95946
rect 521660 95882 521712 95888
rect 520280 62824 520332 62830
rect 520280 62766 520332 62772
rect 520292 4214 520320 62766
rect 520372 26920 520424 26926
rect 520372 26862 520424 26868
rect 520280 4208 520332 4214
rect 520280 4150 520332 4156
rect 520384 3482 520412 26862
rect 521476 4208 521528 4214
rect 521476 4150 521528 4156
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 512012 1414 512132 1442
rect 512012 480 512040 1414
rect 513208 480 513236 3334
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520292 3454 520412 3482
rect 520292 480 520320 3454
rect 521488 480 521516 4150
rect 521672 3482 521700 95882
rect 527836 64870 527864 140762
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 571984 106344 572036 106350
rect 571984 106286 572036 106292
rect 560944 100088 560996 100094
rect 560944 100030 560996 100036
rect 554780 94512 554832 94518
rect 554780 94454 554832 94460
rect 536840 86284 536892 86290
rect 536840 86226 536892 86232
rect 528560 80708 528612 80714
rect 528560 80650 528612 80656
rect 527824 64864 527876 64870
rect 527824 64806 527876 64812
rect 527180 64184 527232 64190
rect 527180 64126 527232 64132
rect 524420 58676 524472 58682
rect 524420 58618 524472 58624
rect 523040 28280 523092 28286
rect 523040 28222 523092 28228
rect 523052 3482 523080 28222
rect 524432 3482 524460 58618
rect 525800 17264 525852 17270
rect 525800 17206 525852 17212
rect 525812 3482 525840 17206
rect 527192 3482 527220 64126
rect 528572 3482 528600 80650
rect 531320 79348 531372 79354
rect 531320 79290 531372 79296
rect 529940 51740 529992 51746
rect 529940 51682 529992 51688
rect 528652 22772 528704 22778
rect 528652 22714 528704 22720
rect 528664 4214 528692 22714
rect 528652 4208 528704 4214
rect 528652 4150 528704 4156
rect 529848 4208 529900 4214
rect 529848 4150 529900 4156
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 525812 3454 526300 3482
rect 527192 3454 527496 3482
rect 528572 3454 528692 3482
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 3454
rect 527468 480 527496 3454
rect 528664 480 528692 3454
rect 529860 480 529888 4150
rect 529952 3482 529980 51682
rect 531332 3482 531360 79290
rect 535460 77988 535512 77994
rect 535460 77930 535512 77936
rect 534080 53100 534132 53106
rect 534080 53042 534132 53048
rect 532700 18624 532752 18630
rect 532700 18566 532752 18572
rect 532712 3482 532740 18566
rect 534092 3482 534120 53042
rect 535472 3482 535500 77930
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536852 3398 536880 86226
rect 545120 84856 545172 84862
rect 545120 84798 545172 84804
rect 542360 66904 542412 66910
rect 542360 66846 542412 66852
rect 538220 65544 538272 65550
rect 538220 65486 538272 65492
rect 536932 14476 536984 14482
rect 536932 14418 536984 14424
rect 536840 3392 536892 3398
rect 536840 3334 536892 3340
rect 536944 480 536972 14418
rect 538232 3482 538260 65486
rect 540980 31068 541032 31074
rect 540980 31010 541032 31016
rect 539600 19984 539652 19990
rect 539600 19926 539652 19932
rect 539612 3482 539640 19926
rect 540992 3482 541020 31010
rect 542372 3482 542400 66846
rect 543740 21412 543792 21418
rect 543740 21354 543792 21360
rect 543752 3482 543780 21354
rect 545132 3482 545160 84798
rect 550640 47592 550692 47598
rect 550640 47534 550692 47540
rect 547880 32428 547932 32434
rect 547880 32370 547932 32376
rect 546592 24132 546644 24138
rect 546592 24074 546644 24080
rect 546500 3800 546552 3806
rect 546500 3742 546552 3748
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 538128 3392 538180 3398
rect 538128 3334 538180 3340
rect 538140 480 538168 3334
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 480 546540 3742
rect 546604 3482 546632 24074
rect 547892 3482 547920 32370
rect 550088 4140 550140 4146
rect 550088 4082 550140 4088
rect 546604 3454 547736 3482
rect 547892 3454 548932 3482
rect 547708 480 547736 3454
rect 548904 480 548932 3454
rect 550100 480 550128 4082
rect 550652 3482 550680 47534
rect 552020 33788 552072 33794
rect 552020 33730 552072 33736
rect 552032 3482 552060 33730
rect 553584 4072 553636 4078
rect 553584 4014 553636 4020
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 4014
rect 554792 480 554820 94454
rect 557540 93152 557592 93158
rect 557540 93094 557592 93100
rect 554872 37936 554924 37942
rect 554872 37878 554924 37884
rect 554884 12442 554912 37878
rect 557552 12442 557580 93094
rect 558920 35216 558972 35222
rect 558920 35158 558972 35164
rect 558932 12442 558960 35158
rect 554872 12436 554924 12442
rect 554872 12378 554924 12384
rect 555976 12436 556028 12442
rect 555976 12378 556028 12384
rect 557540 12436 557592 12442
rect 557540 12378 557592 12384
rect 558368 12436 558420 12442
rect 558368 12378 558420 12384
rect 558920 12436 558972 12442
rect 558920 12378 558972 12384
rect 559564 12436 559616 12442
rect 559564 12378 559616 12384
rect 555988 480 556016 12378
rect 557172 4004 557224 4010
rect 557172 3946 557224 3952
rect 557184 480 557212 3946
rect 558380 480 558408 12378
rect 559576 480 559604 12378
rect 560956 4826 560984 100030
rect 569960 83496 570012 83502
rect 569960 83438 570012 83444
rect 565820 43444 565872 43450
rect 565820 43386 565872 43392
rect 563152 36576 563204 36582
rect 563152 36518 563204 36524
rect 561680 25560 561732 25566
rect 561680 25502 561732 25508
rect 561692 19310 561720 25502
rect 561680 19304 561732 19310
rect 561680 19246 561732 19252
rect 561956 9716 562008 9722
rect 561956 9658 562008 9664
rect 560944 4820 560996 4826
rect 560944 4762 560996 4768
rect 560760 3936 560812 3942
rect 560760 3878 560812 3884
rect 560772 480 560800 3878
rect 561968 480 561996 9658
rect 563164 480 563192 36518
rect 565544 8968 565596 8974
rect 565544 8910 565596 8916
rect 564348 3868 564400 3874
rect 564348 3810 564400 3816
rect 564360 480 564388 3810
rect 565556 480 565584 8910
rect 565832 3482 565860 43386
rect 569040 6180 569092 6186
rect 569040 6122 569092 6128
rect 567200 3664 567252 3670
rect 567200 3606 567252 3612
rect 565832 3454 566780 3482
rect 566752 480 566780 3454
rect 567212 3398 567240 3606
rect 567200 3392 567252 3398
rect 567200 3334 567252 3340
rect 567844 3392 567896 3398
rect 567844 3334 567896 3340
rect 567856 480 567884 3334
rect 569052 480 569080 6122
rect 569972 3482 570000 83438
rect 571996 17950 572024 106286
rect 574744 89004 574796 89010
rect 574744 88946 574796 88952
rect 572720 42084 572772 42090
rect 572720 42026 572772 42032
rect 571984 17944 572036 17950
rect 571984 17886 572036 17892
rect 572628 4820 572680 4826
rect 572628 4762 572680 4768
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 569972 3454 570276 3482
rect 570248 480 570276 3454
rect 571444 480 571472 3538
rect 572640 480 572668 4762
rect 572732 3482 572760 42026
rect 574756 4010 574784 88946
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 581092 11756 581144 11762
rect 581092 11698 581144 11704
rect 579620 10328 579672 10334
rect 579620 10270 579672 10276
rect 576216 7608 576268 7614
rect 576216 7550 576268 7556
rect 574744 4004 574796 4010
rect 574744 3946 574796 3952
rect 575020 3528 575072 3534
rect 572732 3454 573864 3482
rect 575020 3470 575072 3476
rect 573836 480 573864 3454
rect 575032 480 575060 3470
rect 576228 480 576256 7550
rect 577412 4004 577464 4010
rect 577412 3946 577464 3952
rect 577424 480 577452 3946
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 579632 610 579660 10270
rect 581104 626 581132 11698
rect 582196 3732 582248 3738
rect 582196 3674 582248 3680
rect 579620 604 579672 610
rect 579620 546 579672 552
rect 579804 604 579856 610
rect 579804 546 579856 552
rect 581012 598 581132 626
rect 579816 480 579844 546
rect 581012 480 581040 598
rect 582208 480 582236 3674
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3790 682216 3846 682272
rect 3422 667936 3478 667992
rect 3054 653520 3110 653576
rect 3238 624824 3294 624880
rect 3330 595992 3386 596048
rect 3514 610408 3570 610464
rect 3422 567296 3478 567352
rect 3422 553016 3478 553072
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 505006 596264 505062 596320
rect 78678 595856 78734 595912
rect 3514 538600 3570 538656
rect 3422 509904 3478 509960
rect 504638 585112 504694 585168
rect 78678 583888 78734 583944
rect 505006 573996 505008 574016
rect 505008 573996 505060 574016
rect 505060 573996 505062 574016
rect 505006 573960 505062 573996
rect 78678 572056 78734 572112
rect 505006 562980 505008 563000
rect 505008 562980 505060 563000
rect 505060 562980 505062 563000
rect 505006 562944 505062 562980
rect 78678 560088 78734 560144
rect 78678 548256 78734 548312
rect 78678 536288 78734 536344
rect 78678 524456 78734 524512
rect 504178 518508 504180 518528
rect 504180 518508 504232 518528
rect 504232 518508 504234 518528
rect 504178 518472 504234 518508
rect 78678 512488 78734 512544
rect 78678 500656 78734 500712
rect 505006 551792 505062 551848
rect 505006 540640 505062 540696
rect 505006 529624 505062 529680
rect 505006 507320 505062 507376
rect 504362 496304 504418 496360
rect 3514 495488 3570 495544
rect 3422 481072 3478 481128
rect 78678 488688 78734 488744
rect 78678 476856 78734 476912
rect 503718 474000 503774 474056
rect 78678 464888 78734 464944
rect 503810 462984 503866 463040
rect 78678 453056 78734 453112
rect 3422 452376 3478 452432
rect 504178 451832 504234 451888
rect 78678 441088 78734 441144
rect 505006 485152 505062 485208
rect 580170 697992 580226 698048
rect 580262 686296 580318 686352
rect 542358 683168 542414 683224
rect 542726 683168 542782 683224
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 579894 592456 579950 592512
rect 580354 639376 580410 639432
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 580262 545536 580318 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580170 486784 580226 486840
rect 580354 498616 580410 498672
rect 580262 463392 580318 463448
rect 504362 440680 504418 440736
rect 580170 439864 580226 439920
rect 3146 437960 3202 438016
rect 78678 429256 78734 429312
rect 3238 423680 3294 423736
rect 79322 417288 79378 417344
rect 580446 451696 580502 451752
rect 505006 429528 505062 429584
rect 505006 418512 505062 418568
rect 580354 416472 580410 416528
rect 504362 407360 504418 407416
rect 79414 405456 79470 405512
rect 3146 394984 3202 395040
rect 79322 393488 79378 393544
rect 3238 380568 3294 380624
rect 580262 404776 580318 404832
rect 505006 396208 505062 396264
rect 580354 392944 580410 393000
rect 504546 385192 504602 385248
rect 79598 381656 79654 381712
rect 79506 369688 79562 369744
rect 3146 366152 3202 366208
rect 79414 357856 79470 357912
rect 79322 345888 79378 345944
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 3330 308760 3386 308816
rect 505006 374040 505062 374096
rect 580262 369552 580318 369608
rect 505006 362908 505062 362944
rect 505006 362888 505008 362908
rect 505008 362888 505060 362908
rect 505060 362888 505062 362908
rect 580262 357856 580318 357912
rect 504638 351872 504694 351928
rect 580906 346024 580962 346080
rect 505006 340720 505062 340776
rect 79690 333920 79746 333976
rect 79598 322088 79654 322144
rect 79506 310120 79562 310176
rect 79414 298288 79470 298344
rect 3422 294344 3478 294400
rect 79322 286320 79378 286376
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 78678 274488 78734 274544
rect 3146 265648 3202 265704
rect 3422 251232 3478 251288
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 78678 238756 78680 238776
rect 78680 238756 78732 238776
rect 78732 238756 78734 238776
rect 3422 208120 3478 208176
rect 3146 193840 3202 193896
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3514 78920 3570 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 78678 238720 78734 238756
rect 504362 329568 504418 329624
rect 580170 322632 580226 322688
rect 503810 318552 503866 318608
rect 580170 310800 580226 310856
rect 504362 307400 504418 307456
rect 579802 299104 579858 299160
rect 504362 296248 504418 296304
rect 504454 285232 504510 285288
rect 504362 274080 504418 274136
rect 79598 262520 79654 262576
rect 79506 250688 79562 250744
rect 79414 226888 79470 226944
rect 79322 214920 79378 214976
rect 78678 203088 78734 203144
rect 78678 167320 78734 167376
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 504454 262928 504510 262984
rect 504362 240760 504418 240816
rect 579802 252184 579858 252240
rect 504730 251776 504786 251832
rect 504546 229608 504602 229664
rect 504454 207440 504510 207496
rect 504362 196288 504418 196344
rect 79782 191120 79838 191176
rect 79690 179288 79746 179344
rect 79598 155488 79654 155544
rect 79506 143520 79562 143576
rect 78678 131688 78734 131744
rect 79414 119720 79470 119776
rect 79322 107888 79378 107944
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 504638 218456 504694 218512
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 504822 185136 504878 185192
rect 504730 174120 504786 174176
rect 504546 162968 504602 163024
rect 504454 129648 504510 129704
rect 504362 118496 504418 118552
rect 504270 107480 504326 107536
rect 3422 7112 3478 7168
rect 86682 96600 86738 96656
rect 86866 96600 86922 96656
rect 152830 77152 152886 77208
rect 153014 77152 153070 77208
rect 188710 77288 188766 77344
rect 188894 77288 188950 77344
rect 225970 96600 226026 96656
rect 226154 96600 226210 96656
rect 297730 96600 297786 96656
rect 297914 96600 297970 96656
rect 328090 96600 328146 96656
rect 328366 96600 328422 96656
rect 333610 96600 333666 96656
rect 333794 96600 333850 96656
rect 410982 41520 411038 41576
rect 410890 35944 410946 36000
rect 462042 96600 462098 96656
rect 462226 96600 462282 96656
rect 495438 58112 495494 58168
rect 495438 57976 495494 58032
rect 495438 9696 495494 9752
rect 495622 9696 495678 9752
rect 504638 151816 504694 151872
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 505006 140820 505062 140856
rect 505006 140800 505008 140820
rect 505008 140800 505060 140820
rect 505060 140800 505062 140820
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 542353 683226 542419 683229
rect 542721 683226 542787 683229
rect 542353 683224 542787 683226
rect 542353 683168 542358 683224
rect 542414 683168 542726 683224
rect 542782 683168 542787 683224
rect 542353 683166 542787 683168
rect 542353 683163 542419 683166
rect 542721 683163 542787 683166
rect -960 682274 480 682364
rect 3785 682274 3851 682277
rect -960 682272 3851 682274
rect -960 682216 3790 682272
rect 3846 682216 3851 682272
rect -960 682214 3851 682216
rect -960 682124 480 682214
rect 3785 682211 3851 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3233 624882 3299 624885
rect -960 624880 3299 624882
rect -960 624824 3238 624880
rect 3294 624824 3299 624880
rect -960 624822 3299 624824
rect -960 624732 480 624822
rect 3233 624819 3299 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3509 610466 3575 610469
rect -960 610464 3575 610466
rect -960 610408 3514 610464
rect 3570 610408 3575 610464
rect -960 610406 3575 610408
rect -960 610316 480 610406
rect 3509 610403 3575 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 505001 596322 505067 596325
rect 501860 596320 505067 596322
rect 501860 596264 505006 596320
rect 505062 596264 505067 596320
rect 501860 596262 505067 596264
rect 505001 596259 505067 596262
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 78673 595914 78739 595917
rect 78673 595912 82156 595914
rect 78673 595856 78678 595912
rect 78734 595856 82156 595912
rect 78673 595854 82156 595856
rect 78673 595851 78739 595854
rect 579889 592514 579955 592517
rect 583520 592514 584960 592604
rect 579889 592512 584960 592514
rect 579889 592456 579894 592512
rect 579950 592456 584960 592512
rect 579889 592454 584960 592456
rect 579889 592451 579955 592454
rect 583520 592364 584960 592454
rect 504633 585170 504699 585173
rect 501860 585168 504699 585170
rect 501860 585112 504638 585168
rect 504694 585112 504699 585168
rect 501860 585110 504699 585112
rect 504633 585107 504699 585110
rect 78673 583946 78739 583949
rect 78673 583944 82156 583946
rect 78673 583888 78678 583944
rect 78734 583888 82156 583944
rect 78673 583886 82156 583888
rect 78673 583883 78739 583886
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 505001 574018 505067 574021
rect 501860 574016 505067 574018
rect 501860 573960 505006 574016
rect 505062 573960 505067 574016
rect 501860 573958 505067 573960
rect 505001 573955 505067 573958
rect 78673 572114 78739 572117
rect 78673 572112 82156 572114
rect 78673 572056 78678 572112
rect 78734 572056 82156 572112
rect 78673 572054 82156 572056
rect 78673 572051 78739 572054
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 505001 563002 505067 563005
rect 501860 563000 505067 563002
rect 501860 562944 505006 563000
rect 505062 562944 505067 563000
rect 501860 562942 505067 562944
rect 505001 562939 505067 562942
rect 78673 560146 78739 560149
rect 78673 560144 82156 560146
rect 78673 560088 78678 560144
rect 78734 560088 82156 560144
rect 78673 560086 82156 560088
rect 78673 560083 78739 560086
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 505001 551850 505067 551853
rect 501860 551848 505067 551850
rect 501860 551792 505006 551848
rect 505062 551792 505067 551848
rect 501860 551790 505067 551792
rect 505001 551787 505067 551790
rect 78673 548314 78739 548317
rect 78673 548312 82156 548314
rect 78673 548256 78678 548312
rect 78734 548256 82156 548312
rect 78673 548254 82156 548256
rect 78673 548251 78739 548254
rect 580257 545594 580323 545597
rect 583520 545594 584960 545684
rect 580257 545592 584960 545594
rect 580257 545536 580262 545592
rect 580318 545536 584960 545592
rect 580257 545534 584960 545536
rect 580257 545531 580323 545534
rect 583520 545444 584960 545534
rect 505001 540698 505067 540701
rect 501860 540696 505067 540698
rect 501860 540640 505006 540696
rect 505062 540640 505067 540696
rect 501860 540638 505067 540640
rect 505001 540635 505067 540638
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 78673 536346 78739 536349
rect 78673 536344 82156 536346
rect 78673 536288 78678 536344
rect 78734 536288 82156 536344
rect 78673 536286 82156 536288
rect 78673 536283 78739 536286
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 505001 529682 505067 529685
rect 501860 529680 505067 529682
rect 501860 529624 505006 529680
rect 505062 529624 505067 529680
rect 501860 529622 505067 529624
rect 505001 529619 505067 529622
rect 78673 524514 78739 524517
rect 78673 524512 82156 524514
rect 78673 524456 78678 524512
rect 78734 524456 82156 524512
rect 78673 524454 82156 524456
rect 78673 524451 78739 524454
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 504173 518530 504239 518533
rect 501860 518528 504239 518530
rect 501860 518472 504178 518528
rect 504234 518472 504239 518528
rect 501860 518470 504239 518472
rect 504173 518467 504239 518470
rect 78673 512546 78739 512549
rect 78673 512544 82156 512546
rect 78673 512488 78678 512544
rect 78734 512488 82156 512544
rect 78673 512486 82156 512488
rect 78673 512483 78739 512486
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 505001 507378 505067 507381
rect 501860 507376 505067 507378
rect 501860 507320 505006 507376
rect 505062 507320 505067 507376
rect 501860 507318 505067 507320
rect 505001 507315 505067 507318
rect 78673 500714 78739 500717
rect 78673 500712 82156 500714
rect 78673 500656 78678 500712
rect 78734 500656 82156 500712
rect 78673 500654 82156 500656
rect 78673 500651 78739 500654
rect 580349 498674 580415 498677
rect 583520 498674 584960 498764
rect 580349 498672 584960 498674
rect 580349 498616 580354 498672
rect 580410 498616 584960 498672
rect 580349 498614 584960 498616
rect 580349 498611 580415 498614
rect 583520 498524 584960 498614
rect 504357 496362 504423 496365
rect 501860 496360 504423 496362
rect 501860 496304 504362 496360
rect 504418 496304 504423 496360
rect 501860 496302 504423 496304
rect 504357 496299 504423 496302
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 78673 488746 78739 488749
rect 78673 488744 82156 488746
rect 78673 488688 78678 488744
rect 78734 488688 82156 488744
rect 78673 488686 82156 488688
rect 78673 488683 78739 488686
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 505001 485210 505067 485213
rect 501860 485208 505067 485210
rect 501860 485152 505006 485208
rect 505062 485152 505067 485208
rect 501860 485150 505067 485152
rect 505001 485147 505067 485150
rect -960 481130 480 481220
rect 3417 481130 3483 481133
rect -960 481128 3483 481130
rect -960 481072 3422 481128
rect 3478 481072 3483 481128
rect -960 481070 3483 481072
rect -960 480980 480 481070
rect 3417 481067 3483 481070
rect 78673 476914 78739 476917
rect 78673 476912 82156 476914
rect 78673 476856 78678 476912
rect 78734 476856 82156 476912
rect 78673 476854 82156 476856
rect 78673 476851 78739 476854
rect 583520 474996 584960 475236
rect 503713 474058 503779 474061
rect 501860 474056 503779 474058
rect 501860 474000 503718 474056
rect 503774 474000 503779 474056
rect 501860 473998 503779 474000
rect 503713 473995 503779 473998
rect -960 466700 480 466940
rect 78673 464946 78739 464949
rect 78673 464944 82156 464946
rect 78673 464888 78678 464944
rect 78734 464888 82156 464944
rect 78673 464886 82156 464888
rect 78673 464883 78739 464886
rect 580257 463450 580323 463453
rect 583520 463450 584960 463540
rect 580257 463448 584960 463450
rect 580257 463392 580262 463448
rect 580318 463392 584960 463448
rect 580257 463390 584960 463392
rect 580257 463387 580323 463390
rect 583520 463300 584960 463390
rect 503805 463042 503871 463045
rect 501860 463040 503871 463042
rect 501860 462984 503810 463040
rect 503866 462984 503871 463040
rect 501860 462982 503871 462984
rect 503805 462979 503871 462982
rect 78673 453114 78739 453117
rect 78673 453112 82156 453114
rect 78673 453056 78678 453112
rect 78734 453056 82156 453112
rect 78673 453054 82156 453056
rect 78673 453051 78739 453054
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 504173 451890 504239 451893
rect 501860 451888 504239 451890
rect 501860 451832 504178 451888
rect 504234 451832 504239 451888
rect 501860 451830 504239 451832
rect 504173 451827 504239 451830
rect 580441 451754 580507 451757
rect 583520 451754 584960 451844
rect 580441 451752 584960 451754
rect 580441 451696 580446 451752
rect 580502 451696 584960 451752
rect 580441 451694 584960 451696
rect 580441 451691 580507 451694
rect 583520 451604 584960 451694
rect 78673 441146 78739 441149
rect 78673 441144 82156 441146
rect 78673 441088 78678 441144
rect 78734 441088 82156 441144
rect 78673 441086 82156 441088
rect 78673 441083 78739 441086
rect 504357 440738 504423 440741
rect 501860 440736 504423 440738
rect 501860 440680 504362 440736
rect 504418 440680 504423 440736
rect 501860 440678 504423 440680
rect 504357 440675 504423 440678
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 505001 429586 505067 429589
rect 501860 429584 505067 429586
rect 501860 429528 505006 429584
rect 505062 429528 505067 429584
rect 501860 429526 505067 429528
rect 505001 429523 505067 429526
rect 78673 429314 78739 429317
rect 78673 429312 82156 429314
rect 78673 429256 78678 429312
rect 78734 429256 82156 429312
rect 78673 429254 82156 429256
rect 78673 429251 78739 429254
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 505001 418570 505067 418573
rect 501860 418568 505067 418570
rect 501860 418512 505006 418568
rect 505062 418512 505067 418568
rect 501860 418510 505067 418512
rect 505001 418507 505067 418510
rect 79317 417346 79383 417349
rect 79317 417344 82156 417346
rect 79317 417288 79322 417344
rect 79378 417288 82156 417344
rect 79317 417286 82156 417288
rect 79317 417283 79383 417286
rect 580349 416530 580415 416533
rect 583520 416530 584960 416620
rect 580349 416528 584960 416530
rect 580349 416472 580354 416528
rect 580410 416472 584960 416528
rect 580349 416470 584960 416472
rect 580349 416467 580415 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 504357 407418 504423 407421
rect 501860 407416 504423 407418
rect 501860 407360 504362 407416
rect 504418 407360 504423 407416
rect 501860 407358 504423 407360
rect 504357 407355 504423 407358
rect 79409 405514 79475 405517
rect 79409 405512 82156 405514
rect 79409 405456 79414 405512
rect 79470 405456 82156 405512
rect 79409 405454 82156 405456
rect 79409 405451 79475 405454
rect 580257 404834 580323 404837
rect 583520 404834 584960 404924
rect 580257 404832 584960 404834
rect 580257 404776 580262 404832
rect 580318 404776 584960 404832
rect 580257 404774 584960 404776
rect 580257 404771 580323 404774
rect 583520 404684 584960 404774
rect 505001 396266 505067 396269
rect 501860 396264 505067 396266
rect 501860 396208 505006 396264
rect 505062 396208 505067 396264
rect 501860 396206 505067 396208
rect 505001 396203 505067 396206
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 79317 393546 79383 393549
rect 79317 393544 82156 393546
rect 79317 393488 79322 393544
rect 79378 393488 82156 393544
rect 79317 393486 82156 393488
rect 79317 393483 79383 393486
rect 580349 393002 580415 393005
rect 583520 393002 584960 393092
rect 580349 393000 584960 393002
rect 580349 392944 580354 393000
rect 580410 392944 584960 393000
rect 580349 392942 584960 392944
rect 580349 392939 580415 392942
rect 583520 392852 584960 392942
rect 504541 385250 504607 385253
rect 501860 385248 504607 385250
rect 501860 385192 504546 385248
rect 504602 385192 504607 385248
rect 501860 385190 504607 385192
rect 504541 385187 504607 385190
rect 79593 381714 79659 381717
rect 79593 381712 82156 381714
rect 79593 381656 79598 381712
rect 79654 381656 82156 381712
rect 79593 381654 82156 381656
rect 79593 381651 79659 381654
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 505001 374098 505067 374101
rect 501860 374096 505067 374098
rect 501860 374040 505006 374096
rect 505062 374040 505067 374096
rect 501860 374038 505067 374040
rect 505001 374035 505067 374038
rect 79501 369746 79567 369749
rect 79501 369744 82156 369746
rect 79501 369688 79506 369744
rect 79562 369688 82156 369744
rect 79501 369686 82156 369688
rect 79501 369683 79567 369686
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 505001 362946 505067 362949
rect 501860 362944 505067 362946
rect 501860 362888 505006 362944
rect 505062 362888 505067 362944
rect 501860 362886 505067 362888
rect 505001 362883 505067 362886
rect 79409 357914 79475 357917
rect 580257 357914 580323 357917
rect 583520 357914 584960 358004
rect 79409 357912 82156 357914
rect 79409 357856 79414 357912
rect 79470 357856 82156 357912
rect 79409 357854 82156 357856
rect 580257 357912 584960 357914
rect 580257 357856 580262 357912
rect 580318 357856 584960 357912
rect 580257 357854 584960 357856
rect 79409 357851 79475 357854
rect 580257 357851 580323 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 504633 351930 504699 351933
rect 501860 351928 504699 351930
rect 501860 351872 504638 351928
rect 504694 351872 504699 351928
rect 501860 351870 504699 351872
rect 504633 351867 504699 351870
rect 580901 346082 580967 346085
rect 583520 346082 584960 346172
rect 580901 346080 584960 346082
rect 580901 346024 580906 346080
rect 580962 346024 584960 346080
rect 580901 346022 584960 346024
rect 580901 346019 580967 346022
rect 79317 345946 79383 345949
rect 79317 345944 82156 345946
rect 79317 345888 79322 345944
rect 79378 345888 82156 345944
rect 583520 345932 584960 346022
rect 79317 345886 82156 345888
rect 79317 345883 79383 345886
rect 505001 340778 505067 340781
rect 501860 340776 505067 340778
rect 501860 340720 505006 340776
rect 505062 340720 505067 340776
rect 501860 340718 505067 340720
rect 505001 340715 505067 340718
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 583520 334236 584960 334476
rect 79685 333978 79751 333981
rect 79685 333976 82156 333978
rect 79685 333920 79690 333976
rect 79746 333920 82156 333976
rect 79685 333918 82156 333920
rect 79685 333915 79751 333918
rect 504357 329626 504423 329629
rect 501860 329624 504423 329626
rect 501860 329568 504362 329624
rect 504418 329568 504423 329624
rect 501860 329566 504423 329568
rect 504357 329563 504423 329566
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 79593 322146 79659 322149
rect 79593 322144 82156 322146
rect 79593 322088 79598 322144
rect 79654 322088 82156 322144
rect 79593 322086 82156 322088
rect 79593 322083 79659 322086
rect 503805 318610 503871 318613
rect 501860 318608 503871 318610
rect 501860 318552 503810 318608
rect 503866 318552 503871 318608
rect 501860 318550 503871 318552
rect 503805 318547 503871 318550
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 79501 310178 79567 310181
rect 79501 310176 82156 310178
rect 79501 310120 79506 310176
rect 79562 310120 82156 310176
rect 79501 310118 82156 310120
rect 79501 310115 79567 310118
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 504357 307458 504423 307461
rect 501860 307456 504423 307458
rect 501860 307400 504362 307456
rect 504418 307400 504423 307456
rect 501860 307398 504423 307400
rect 504357 307395 504423 307398
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 79409 298346 79475 298349
rect 79409 298344 82156 298346
rect 79409 298288 79414 298344
rect 79470 298288 82156 298344
rect 79409 298286 82156 298288
rect 79409 298283 79475 298286
rect 504357 296306 504423 296309
rect 501860 296304 504423 296306
rect 501860 296248 504362 296304
rect 504418 296248 504423 296304
rect 501860 296246 504423 296248
rect 504357 296243 504423 296246
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 583520 287316 584960 287556
rect 79317 286378 79383 286381
rect 79317 286376 82156 286378
rect 79317 286320 79322 286376
rect 79378 286320 82156 286376
rect 79317 286318 82156 286320
rect 79317 286315 79383 286318
rect 504449 285290 504515 285293
rect 501860 285288 504515 285290
rect 501860 285232 504454 285288
rect 504510 285232 504515 285288
rect 501860 285230 504515 285232
rect 504449 285227 504515 285230
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 78673 274546 78739 274549
rect 78673 274544 82156 274546
rect 78673 274488 78678 274544
rect 78734 274488 82156 274544
rect 78673 274486 82156 274488
rect 78673 274483 78739 274486
rect 504357 274138 504423 274141
rect 501860 274136 504423 274138
rect 501860 274080 504362 274136
rect 504418 274080 504423 274136
rect 501860 274078 504423 274080
rect 504357 274075 504423 274078
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 504449 262986 504515 262989
rect 501860 262984 504515 262986
rect 501860 262928 504454 262984
rect 504510 262928 504515 262984
rect 501860 262926 504515 262928
rect 504449 262923 504515 262926
rect 79593 262578 79659 262581
rect 79593 262576 82156 262578
rect 79593 262520 79598 262576
rect 79654 262520 82156 262576
rect 79593 262518 82156 262520
rect 79593 262515 79659 262518
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect 504725 251834 504791 251837
rect 501860 251832 504791 251834
rect 501860 251776 504730 251832
rect 504786 251776 504791 251832
rect 501860 251774 504791 251776
rect 504725 251771 504791 251774
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 79501 250746 79567 250749
rect 79501 250744 82156 250746
rect 79501 250688 79506 250744
rect 79562 250688 82156 250744
rect 79501 250686 82156 250688
rect 79501 250683 79567 250686
rect 504357 240818 504423 240821
rect 501860 240816 504423 240818
rect 501860 240760 504362 240816
rect 504418 240760 504423 240816
rect 501860 240758 504423 240760
rect 504357 240755 504423 240758
rect 583520 240396 584960 240636
rect 78673 238778 78739 238781
rect 78673 238776 82156 238778
rect 78673 238720 78678 238776
rect 78734 238720 82156 238776
rect 78673 238718 82156 238720
rect 78673 238715 78739 238718
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 504541 229666 504607 229669
rect 501860 229664 504607 229666
rect 501860 229608 504546 229664
rect 504602 229608 504607 229664
rect 501860 229606 504607 229608
rect 504541 229603 504607 229606
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 79409 226946 79475 226949
rect 79409 226944 82156 226946
rect 79409 226888 79414 226944
rect 79470 226888 82156 226944
rect 79409 226886 82156 226888
rect 79409 226883 79475 226886
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 504633 218514 504699 218517
rect 501860 218512 504699 218514
rect 501860 218456 504638 218512
rect 504694 218456 504699 218512
rect 501860 218454 504699 218456
rect 504633 218451 504699 218454
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 79317 214978 79383 214981
rect 79317 214976 82156 214978
rect 79317 214920 79322 214976
rect 79378 214920 82156 214976
rect 79317 214918 82156 214920
rect 79317 214915 79383 214918
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 504449 207498 504515 207501
rect 501860 207496 504515 207498
rect 501860 207440 504454 207496
rect 504510 207440 504515 207496
rect 501860 207438 504515 207440
rect 504449 207435 504515 207438
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 78673 203146 78739 203149
rect 78673 203144 82156 203146
rect 78673 203088 78678 203144
rect 78734 203088 82156 203144
rect 78673 203086 82156 203088
rect 78673 203083 78739 203086
rect 504357 196346 504423 196349
rect 501860 196344 504423 196346
rect 501860 196288 504362 196344
rect 504418 196288 504423 196344
rect 501860 196286 504423 196288
rect 504357 196283 504423 196286
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 79777 191178 79843 191181
rect 79777 191176 82156 191178
rect 79777 191120 79782 191176
rect 79838 191120 82156 191176
rect 79777 191118 82156 191120
rect 79777 191115 79843 191118
rect 504817 185194 504883 185197
rect 501860 185192 504883 185194
rect 501860 185136 504822 185192
rect 504878 185136 504883 185192
rect 501860 185134 504883 185136
rect 504817 185131 504883 185134
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 79685 179346 79751 179349
rect 79685 179344 82156 179346
rect 79685 179288 79690 179344
rect 79746 179288 82156 179344
rect 79685 179286 82156 179288
rect 79685 179283 79751 179286
rect 504725 174178 504791 174181
rect 501860 174176 504791 174178
rect 501860 174120 504730 174176
rect 504786 174120 504791 174176
rect 501860 174118 504791 174120
rect 504725 174115 504791 174118
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 78673 167378 78739 167381
rect 78673 167376 82156 167378
rect 78673 167320 78678 167376
rect 78734 167320 82156 167376
rect 78673 167318 82156 167320
rect 78673 167315 78739 167318
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 504541 163026 504607 163029
rect 501860 163024 504607 163026
rect 501860 162968 504546 163024
rect 504602 162968 504607 163024
rect 501860 162966 504607 162968
rect 504541 162963 504607 162966
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 79593 155546 79659 155549
rect 79593 155544 82156 155546
rect 79593 155488 79598 155544
rect 79654 155488 82156 155544
rect 79593 155486 82156 155488
rect 79593 155483 79659 155486
rect 504633 151874 504699 151877
rect 501860 151872 504699 151874
rect 501860 151816 504638 151872
rect 504694 151816 504699 151872
rect 501860 151814 504699 151816
rect 504633 151811 504699 151814
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 79501 143578 79567 143581
rect 79501 143576 82156 143578
rect 79501 143520 79506 143576
rect 79562 143520 82156 143576
rect 79501 143518 82156 143520
rect 79501 143515 79567 143518
rect 505001 140858 505067 140861
rect 501860 140856 505067 140858
rect 501860 140800 505006 140856
rect 505062 140800 505067 140856
rect 501860 140798 505067 140800
rect 505001 140795 505067 140798
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 78673 131746 78739 131749
rect 78673 131744 82156 131746
rect 78673 131688 78678 131744
rect 78734 131688 82156 131744
rect 78673 131686 82156 131688
rect 78673 131683 78739 131686
rect 504449 129706 504515 129709
rect 501860 129704 504515 129706
rect 501860 129648 504454 129704
rect 504510 129648 504515 129704
rect 501860 129646 504515 129648
rect 504449 129643 504515 129646
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 79409 119778 79475 119781
rect 79409 119776 82156 119778
rect 79409 119720 79414 119776
rect 79470 119720 82156 119776
rect 79409 119718 82156 119720
rect 79409 119715 79475 119718
rect 504357 118554 504423 118557
rect 501860 118552 504423 118554
rect 501860 118496 504362 118552
rect 504418 118496 504423 118552
rect 501860 118494 504423 118496
rect 504357 118491 504423 118494
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect 79317 107946 79383 107949
rect 79317 107944 82156 107946
rect 79317 107888 79322 107944
rect 79378 107888 82156 107944
rect 79317 107886 82156 107888
rect 79317 107883 79383 107886
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 504265 107538 504331 107541
rect 501860 107536 504331 107538
rect 501860 107480 504270 107536
rect 504326 107480 504331 107536
rect 501860 107478 504331 107480
rect 504265 107475 504331 107478
rect 583520 99636 584960 99876
rect 86677 96658 86743 96661
rect 86861 96658 86927 96661
rect 86677 96656 86927 96658
rect 86677 96600 86682 96656
rect 86738 96600 86866 96656
rect 86922 96600 86927 96656
rect 86677 96598 86927 96600
rect 86677 96595 86743 96598
rect 86861 96595 86927 96598
rect 225965 96658 226031 96661
rect 226149 96658 226215 96661
rect 225965 96656 226215 96658
rect 225965 96600 225970 96656
rect 226026 96600 226154 96656
rect 226210 96600 226215 96656
rect 225965 96598 226215 96600
rect 225965 96595 226031 96598
rect 226149 96595 226215 96598
rect 297725 96658 297791 96661
rect 297909 96658 297975 96661
rect 297725 96656 297975 96658
rect 297725 96600 297730 96656
rect 297786 96600 297914 96656
rect 297970 96600 297975 96656
rect 297725 96598 297975 96600
rect 297725 96595 297791 96598
rect 297909 96595 297975 96598
rect 328085 96658 328151 96661
rect 328361 96658 328427 96661
rect 328085 96656 328427 96658
rect 328085 96600 328090 96656
rect 328146 96600 328366 96656
rect 328422 96600 328427 96656
rect 328085 96598 328427 96600
rect 328085 96595 328151 96598
rect 328361 96595 328427 96598
rect 333605 96658 333671 96661
rect 333789 96658 333855 96661
rect 333605 96656 333855 96658
rect 333605 96600 333610 96656
rect 333666 96600 333794 96656
rect 333850 96600 333855 96656
rect 333605 96598 333855 96600
rect 333605 96595 333671 96598
rect 333789 96595 333855 96598
rect 462037 96658 462103 96661
rect 462221 96658 462287 96661
rect 462037 96656 462287 96658
rect 462037 96600 462042 96656
rect 462098 96600 462226 96656
rect 462282 96600 462287 96656
rect 462037 96598 462287 96600
rect 462037 96595 462103 96598
rect 462221 96595 462287 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 188705 77346 188771 77349
rect 188889 77346 188955 77349
rect 188705 77344 188955 77346
rect 188705 77288 188710 77344
rect 188766 77288 188894 77344
rect 188950 77288 188955 77344
rect 188705 77286 188955 77288
rect 188705 77283 188771 77286
rect 188889 77283 188955 77286
rect 152825 77210 152891 77213
rect 153009 77210 153075 77213
rect 152825 77208 153075 77210
rect 152825 77152 152830 77208
rect 152886 77152 153014 77208
rect 153070 77152 153075 77208
rect 152825 77150 153075 77152
rect 152825 77147 152891 77150
rect 153009 77147 153075 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 495433 58170 495499 58173
rect 495433 58168 495634 58170
rect 495433 58112 495438 58168
rect 495494 58112 495634 58168
rect 495433 58110 495634 58112
rect 495433 58107 495499 58110
rect 495433 58034 495499 58037
rect 495574 58034 495634 58110
rect 495433 58032 495634 58034
rect 495433 57976 495438 58032
rect 495494 57976 495634 58032
rect 495433 57974 495634 57976
rect 495433 57971 495499 57974
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 410977 41580 411043 41581
rect 410926 41578 410932 41580
rect 410886 41518 410932 41578
rect 410996 41576 411043 41580
rect 411038 41520 411043 41576
rect 410926 41516 410932 41518
rect 410996 41516 411043 41520
rect 410977 41515 411043 41516
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 410885 36004 410951 36005
rect 410885 36000 410932 36004
rect 410996 36002 411002 36004
rect -960 35866 480 35956
rect 410885 35944 410890 36000
rect 410885 35940 410932 35944
rect 410996 35942 411042 36002
rect 410996 35940 411002 35942
rect 410885 35939 410951 35940
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 495433 9754 495499 9757
rect 495617 9754 495683 9757
rect 495433 9752 495683 9754
rect 495433 9696 495438 9752
rect 495494 9696 495622 9752
rect 495678 9696 495683 9752
rect 495433 9694 495683 9696
rect 495433 9691 495499 9694
rect 495617 9691 495683 9694
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< via3 >>
rect 410932 41576 410996 41580
rect 410932 41520 410982 41576
rect 410982 41520 410996 41576
rect 410932 41516 410996 41520
rect 410932 36000 410996 36004
rect 410932 35944 410946 36000
rect 410946 35944 410996 36000
rect 410932 35940 410996 35944
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 602000 84204 624698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 602000 91404 631898
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 602000 95004 635498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 602000 98604 603098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 602000 102204 606698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 602000 109404 613898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 602000 113004 617498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 602000 116604 621098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 602000 120204 624698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 602000 127404 631898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 602000 131004 635498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 602000 134604 603098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 602000 138204 606698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 602000 145404 613898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 602000 149004 617498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 602000 152604 621098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 602000 156204 624698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 602000 163404 631898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 602000 167004 635498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 602000 170604 603098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 602000 174204 606698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 602000 181404 613898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 602000 185004 617498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 602000 188604 621098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 602000 192204 624698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 602000 199404 631898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 602000 203004 635498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 602000 206604 603098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 602000 210204 606698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 602000 217404 613898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 602000 221004 617498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 602000 224604 621098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 602000 228204 624698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 602000 235404 631898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 602000 239004 635498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 602000 242604 603098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 602000 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 602000 253404 613898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 602000 257004 617498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 602000 260604 621098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 602000 264204 624698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 602000 271404 631898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 602000 275004 635498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 602000 278604 603098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 602000 282204 606698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 602000 289404 613898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 602000 293004 617498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 602000 296604 621098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 602000 300204 624698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 602000 307404 631898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 602000 311004 635498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 602000 314604 603098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 602000 318204 606698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 602000 325404 613898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 602000 329004 617498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 602000 332604 621098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 602000 336204 624698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 602000 343404 631898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 602000 347004 635498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 602000 350604 603098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 602000 354204 606698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 602000 361404 613898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 602000 365004 617498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 602000 368604 621098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 602000 372204 624698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 602000 379404 631898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 602000 383004 635498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 602000 386604 603098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 602000 390204 606698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 602000 397404 613898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 602000 401004 617498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 602000 404604 621098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 602000 408204 624698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 602000 415404 631898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 602000 419004 635498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 602000 422604 603098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 602000 426204 606698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 602000 433404 613898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 602000 437004 617498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 602000 440604 621098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 602000 444204 624698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 602000 451404 631898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 602000 455004 635498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 602000 458604 603098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 602000 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 602000 469404 613898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 602000 473004 617498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 602000 476604 621098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 602000 480204 624698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 602000 487404 631898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 602000 491004 635498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 602000 494604 603098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 602000 498204 606698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 85254 84204 102000
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 92454 91404 102000
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 96054 95004 102000
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 99654 98604 102000
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 67254 102204 102000
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 74454 109404 102000
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 78054 113004 102000
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 81654 116604 102000
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 85254 120204 102000
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 92454 127404 102000
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 96054 131004 102000
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 99654 134604 102000
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 67254 138204 102000
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 74454 145404 102000
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 78054 149004 102000
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 81654 152604 102000
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 85254 156204 102000
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 92454 163404 102000
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 96054 167004 102000
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 99654 170604 102000
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 67254 174204 102000
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 74454 181404 102000
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 78054 185004 102000
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 81654 188604 102000
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 85254 192204 102000
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 92454 199404 102000
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 96054 203004 102000
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 99654 206604 102000
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 67254 210204 102000
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 74454 217404 102000
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 78054 221004 102000
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 81654 224604 102000
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 85254 228204 102000
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 92454 235404 102000
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 96054 239004 102000
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 99654 242604 102000
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 67254 246204 102000
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 74454 253404 102000
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 78054 257004 102000
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 81654 260604 102000
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 85254 264204 102000
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 92454 271404 102000
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 96054 275004 102000
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 99654 278604 102000
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 67254 282204 102000
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 102000
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 78054 293004 102000
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 81654 296604 102000
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 85254 300204 102000
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 92454 307404 102000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 96054 311004 102000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 99654 314604 102000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 67254 318204 102000
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 74454 325404 102000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 78054 329004 102000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 81654 332604 102000
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 85254 336204 102000
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 92454 343404 102000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 96054 347004 102000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 99654 350604 102000
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 67254 354204 102000
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 74454 361404 102000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 78054 365004 102000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 81654 368604 102000
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 85254 372204 102000
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 92454 379404 102000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 96054 383004 102000
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 99654 386604 102000
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 67254 390204 102000
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 74454 397404 102000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 78054 401004 102000
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 81654 404604 102000
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 85254 408204 102000
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 414804 92454 415404 102000
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 410931 41580 410997 41581
rect 410931 41516 410932 41580
rect 410996 41516 410997 41580
rect 410931 41515 410997 41516
rect 410934 36005 410994 41515
rect 410931 36004 410997 36005
rect 410931 35940 410932 36004
rect 410996 35940 410997 36004
rect 410931 35939 410997 35940
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 96054 419004 102000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 99654 422604 102000
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 67254 426204 102000
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 74454 433404 102000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 78054 437004 102000
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 81654 440604 102000
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 85254 444204 102000
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 92454 451404 102000
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 96054 455004 102000
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 99654 458604 102000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 67254 462204 102000
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 74454 469404 102000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 78054 473004 102000
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 81654 476604 102000
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 85254 480204 102000
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 92454 487404 102000
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 96054 491004 102000
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 99654 494604 102000
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 67254 498204 102000
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use Ibtida_top_dffram_cv  mprj
timestamp 1607603059
transform 1 0 82000 0 1 102000
box 0 0 420000 500000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
