magic
tech sky130A
magscale 1 2
timestamp 1607975982
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 412649 683247 412683 692733
rect 283297 666587 283331 683077
rect 299857 666587 299891 683077
rect 413017 666587 413051 683077
rect 429577 666587 429611 683077
rect 542737 666587 542771 683077
rect 559297 666587 559331 683077
rect 72985 647275 73019 656829
rect 73077 616879 73111 626501
rect 283113 601715 283147 608549
rect 299673 601715 299707 608549
rect 412833 601715 412867 608549
rect 429393 601715 429427 608549
rect 542553 601715 542587 608549
rect 559113 601715 559147 608549
rect 72893 589339 72927 598893
rect 283297 589339 283331 598893
rect 299857 589339 299891 598893
rect 413017 589339 413051 598893
rect 429577 589339 429611 598893
rect 542737 589339 542771 598893
rect 559297 589339 559331 598893
rect 8033 579751 8067 589237
rect 137753 579751 137787 589237
rect 154313 579751 154347 589237
rect 218069 579683 218103 589237
rect 234629 579683 234663 589237
rect 347789 579683 347823 589237
rect 364349 579683 364383 589237
rect 477509 579683 477543 589237
rect 494069 579683 494103 589237
rect 72617 569959 72651 579581
rect 137569 569959 137603 579581
rect 218161 563091 218195 569857
rect 234721 563091 234755 569857
rect 347881 563091 347915 569857
rect 364441 563091 364475 569857
rect 477601 563091 477635 569857
rect 494161 563091 494195 569857
rect 72617 550647 72651 553401
rect 137661 550647 137695 560201
rect 283021 550647 283055 560201
rect 412741 550647 412775 560201
rect 429301 550647 429335 560201
rect 542461 550647 542495 560201
rect 559021 550647 559055 560201
rect 8033 540991 8067 550545
rect 72617 531335 72651 534089
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 283113 485775 283147 492609
rect 299673 485775 299707 492609
rect 412833 485775 412867 492609
rect 429393 485775 429427 492609
rect 542553 485775 542587 492609
rect 559113 485775 559147 492609
rect 283113 466395 283147 473297
rect 299673 466395 299707 473297
rect 412833 466395 412867 473297
rect 429393 466395 429427 473297
rect 542553 466395 542587 473297
rect 559113 466395 559147 473297
rect 299581 447083 299615 453917
rect 8125 437427 8159 444329
rect 137845 437427 137879 444329
rect 154405 437427 154439 444329
rect 283113 427771 283147 434673
rect 299673 427771 299707 434673
rect 412833 427771 412867 434673
rect 429393 427771 429427 434673
rect 542553 427771 542587 434673
rect 559113 427771 559147 434673
rect 198013 95251 198047 100045
rect 370881 99331 370915 102085
rect 92213 85595 92247 89709
rect 198013 85595 198047 95081
rect 198565 85595 198599 89709
rect 227453 87023 227487 89709
rect 267013 89675 267047 96577
rect 278605 87023 278639 96577
rect 342085 87023 342119 98549
rect 92213 67643 92247 80733
rect 104633 77367 104667 82093
rect 104541 67643 104575 77197
rect 151553 67643 151587 77197
rect 198013 75939 198047 80189
rect 239873 77367 239907 81821
rect 267105 77299 267139 80121
rect 239781 67643 239815 77197
rect 518909 75939 518943 85493
rect 532709 75939 532743 85493
rect 267105 67643 267139 70397
rect 274557 67643 274591 71145
rect 92121 48331 92155 57885
rect 96261 56627 96295 66181
rect 200129 56627 200163 66181
rect 239873 57987 239907 62917
rect 267105 57987 267139 62713
rect 341901 56627 341935 66181
rect 518909 56627 518943 66181
rect 532709 56627 532743 66181
rect 569969 56627 570003 65501
rect 96261 46971 96295 56457
rect 239689 48331 239723 51085
rect 267105 48331 267139 51085
rect 267749 46971 267783 53125
rect 138029 37315 138063 46869
rect 200129 37315 200163 46869
rect 267013 38675 267047 41497
rect 509249 37315 509283 46869
rect 518909 37315 518943 46869
rect 527189 37315 527223 46869
rect 532709 37315 532743 46869
rect 567853 38675 567887 48229
rect 569969 37315 570003 46869
rect 198105 19363 198139 28917
rect 215033 27659 215067 37213
rect 227361 27659 227395 37213
rect 198749 9707 198783 27421
rect 200129 9707 200163 22797
rect 267105 19363 267139 28917
rect 267749 9707 267783 22661
rect 491309 9707 491343 19261
rect 492689 9707 492723 19261
rect 509249 9707 509283 27557
rect 510629 9707 510663 19261
rect 516149 9707 516183 19261
rect 518909 18003 518943 27557
rect 527189 18003 527223 27557
rect 532709 9707 532743 27557
rect 550649 12359 550683 19261
rect 553409 9707 553443 19261
rect 568037 18003 568071 27557
rect 569969 9707 570003 27557
rect 144837 4879 144871 8653
rect 154589 3927 154623 4845
rect 486525 3451 486559 7293
rect 511951 3485 512043 3519
rect 499589 3315 499623 3417
rect 509157 3315 509191 3485
rect 512009 3451 512043 3485
rect 517897 595 517931 9605
rect 518909 3451 518943 3553
rect 519093 595 519127 9605
rect 528477 3451 528511 3553
rect 545313 595 545347 9605
rect 548901 595 548935 9605
rect 550097 595 550131 9605
rect 559021 3315 559055 3485
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 412649 692733 412683 692767
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 412649 683213 412683 683247
rect 154313 676209 154347 676243
rect 283297 683077 283331 683111
rect 72801 676073 72835 676107
rect 283297 666553 283331 666587
rect 299857 683077 299891 683111
rect 299857 666553 299891 666587
rect 413017 683077 413051 683111
rect 413017 666553 413051 666587
rect 429577 683077 429611 683111
rect 429577 666553 429611 666587
rect 542737 683077 542771 683111
rect 542737 666553 542771 666587
rect 559297 683077 559331 683111
rect 559297 666553 559331 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 73077 626501 73111 626535
rect 73077 616845 73111 616879
rect 283113 608549 283147 608583
rect 283113 601681 283147 601715
rect 299673 608549 299707 608583
rect 299673 601681 299707 601715
rect 412833 608549 412867 608583
rect 412833 601681 412867 601715
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 542553 608549 542587 608583
rect 542553 601681 542587 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 72893 598893 72927 598927
rect 72893 589305 72927 589339
rect 283297 598893 283331 598927
rect 283297 589305 283331 589339
rect 299857 598893 299891 598927
rect 299857 589305 299891 589339
rect 413017 598893 413051 598927
rect 413017 589305 413051 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 542737 598893 542771 598927
rect 542737 589305 542771 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 8033 589237 8067 589271
rect 8033 579717 8067 579751
rect 137753 589237 137787 589271
rect 137753 579717 137787 579751
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 218069 589237 218103 589271
rect 218069 579649 218103 579683
rect 234629 589237 234663 589271
rect 234629 579649 234663 579683
rect 347789 589237 347823 589271
rect 347789 579649 347823 579683
rect 364349 589237 364383 589271
rect 364349 579649 364383 579683
rect 477509 589237 477543 589271
rect 477509 579649 477543 579683
rect 494069 589237 494103 589271
rect 494069 579649 494103 579683
rect 72617 579581 72651 579615
rect 72617 569925 72651 569959
rect 137569 579581 137603 579615
rect 137569 569925 137603 569959
rect 218161 569857 218195 569891
rect 218161 563057 218195 563091
rect 234721 569857 234755 569891
rect 234721 563057 234755 563091
rect 347881 569857 347915 569891
rect 347881 563057 347915 563091
rect 364441 569857 364475 569891
rect 364441 563057 364475 563091
rect 477601 569857 477635 569891
rect 477601 563057 477635 563091
rect 494161 569857 494195 569891
rect 494161 563057 494195 563091
rect 137661 560201 137695 560235
rect 72617 553401 72651 553435
rect 72617 550613 72651 550647
rect 137661 550613 137695 550647
rect 283021 560201 283055 560235
rect 283021 550613 283055 550647
rect 412741 560201 412775 560235
rect 412741 550613 412775 550647
rect 429301 560201 429335 560235
rect 429301 550613 429335 550647
rect 542461 560201 542495 560235
rect 542461 550613 542495 550647
rect 559021 560201 559055 560235
rect 559021 550613 559055 550647
rect 8033 550545 8067 550579
rect 8033 540957 8067 540991
rect 72617 534089 72651 534123
rect 72617 531301 72651 531335
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 154405 502333 154439 502367
rect 283113 492609 283147 492643
rect 283113 485741 283147 485775
rect 299673 492609 299707 492643
rect 299673 485741 299707 485775
rect 412833 492609 412867 492643
rect 412833 485741 412867 485775
rect 429393 492609 429427 492643
rect 429393 485741 429427 485775
rect 542553 492609 542587 492643
rect 542553 485741 542587 485775
rect 559113 492609 559147 492643
rect 559113 485741 559147 485775
rect 283113 473297 283147 473331
rect 283113 466361 283147 466395
rect 299673 473297 299707 473331
rect 299673 466361 299707 466395
rect 412833 473297 412867 473331
rect 412833 466361 412867 466395
rect 429393 473297 429427 473331
rect 429393 466361 429427 466395
rect 542553 473297 542587 473331
rect 542553 466361 542587 466395
rect 559113 473297 559147 473331
rect 559113 466361 559147 466395
rect 299581 453917 299615 453951
rect 299581 447049 299615 447083
rect 8125 444329 8159 444363
rect 8125 437393 8159 437427
rect 137845 444329 137879 444363
rect 137845 437393 137879 437427
rect 154405 444329 154439 444363
rect 154405 437393 154439 437427
rect 283113 434673 283147 434707
rect 283113 427737 283147 427771
rect 299673 434673 299707 434707
rect 299673 427737 299707 427771
rect 412833 434673 412867 434707
rect 412833 427737 412867 427771
rect 429393 434673 429427 434707
rect 429393 427737 429427 427771
rect 542553 434673 542587 434707
rect 542553 427737 542587 427771
rect 559113 434673 559147 434707
rect 559113 427737 559147 427771
rect 370881 102085 370915 102119
rect 198013 100045 198047 100079
rect 370881 99297 370915 99331
rect 342085 98549 342119 98583
rect 198013 95217 198047 95251
rect 267013 96577 267047 96611
rect 198013 95081 198047 95115
rect 92213 89709 92247 89743
rect 92213 85561 92247 85595
rect 198013 85561 198047 85595
rect 198565 89709 198599 89743
rect 227453 89709 227487 89743
rect 267013 89641 267047 89675
rect 278605 96577 278639 96611
rect 227453 86989 227487 87023
rect 278605 86989 278639 87023
rect 342085 86989 342119 87023
rect 198565 85561 198599 85595
rect 518909 85493 518943 85527
rect 104633 82093 104667 82127
rect 92213 80733 92247 80767
rect 239873 81821 239907 81855
rect 104633 77333 104667 77367
rect 198013 80189 198047 80223
rect 92213 67609 92247 67643
rect 104541 77197 104575 77231
rect 104541 67609 104575 67643
rect 151553 77197 151587 77231
rect 239873 77333 239907 77367
rect 267105 80121 267139 80155
rect 267105 77265 267139 77299
rect 198013 75905 198047 75939
rect 239781 77197 239815 77231
rect 151553 67609 151587 67643
rect 518909 75905 518943 75939
rect 532709 85493 532743 85527
rect 532709 75905 532743 75939
rect 274557 71145 274591 71179
rect 239781 67609 239815 67643
rect 267105 70397 267139 70431
rect 267105 67609 267139 67643
rect 274557 67609 274591 67643
rect 96261 66181 96295 66215
rect 92121 57885 92155 57919
rect 96261 56593 96295 56627
rect 200129 66181 200163 66215
rect 341901 66181 341935 66215
rect 239873 62917 239907 62951
rect 239873 57953 239907 57987
rect 267105 62713 267139 62747
rect 267105 57953 267139 57987
rect 200129 56593 200163 56627
rect 341901 56593 341935 56627
rect 518909 66181 518943 66215
rect 518909 56593 518943 56627
rect 532709 66181 532743 66215
rect 532709 56593 532743 56627
rect 569969 65501 570003 65535
rect 569969 56593 570003 56627
rect 92121 48297 92155 48331
rect 96261 56457 96295 56491
rect 267749 53125 267783 53159
rect 239689 51085 239723 51119
rect 239689 48297 239723 48331
rect 267105 51085 267139 51119
rect 267105 48297 267139 48331
rect 96261 46937 96295 46971
rect 267749 46937 267783 46971
rect 567853 48229 567887 48263
rect 138029 46869 138063 46903
rect 138029 37281 138063 37315
rect 200129 46869 200163 46903
rect 509249 46869 509283 46903
rect 267013 41497 267047 41531
rect 267013 38641 267047 38675
rect 200129 37281 200163 37315
rect 509249 37281 509283 37315
rect 518909 46869 518943 46903
rect 518909 37281 518943 37315
rect 527189 46869 527223 46903
rect 527189 37281 527223 37315
rect 532709 46869 532743 46903
rect 567853 38641 567887 38675
rect 569969 46869 570003 46903
rect 532709 37281 532743 37315
rect 569969 37281 570003 37315
rect 215033 37213 215067 37247
rect 198105 28917 198139 28951
rect 215033 27625 215067 27659
rect 227361 37213 227395 37247
rect 227361 27625 227395 27659
rect 267105 28917 267139 28951
rect 198105 19329 198139 19363
rect 198749 27421 198783 27455
rect 198749 9673 198783 9707
rect 200129 22797 200163 22831
rect 509249 27557 509283 27591
rect 267105 19329 267139 19363
rect 267749 22661 267783 22695
rect 200129 9673 200163 9707
rect 267749 9673 267783 9707
rect 491309 19261 491343 19295
rect 491309 9673 491343 9707
rect 492689 19261 492723 19295
rect 492689 9673 492723 9707
rect 518909 27557 518943 27591
rect 509249 9673 509283 9707
rect 510629 19261 510663 19295
rect 510629 9673 510663 9707
rect 516149 19261 516183 19295
rect 518909 17969 518943 18003
rect 527189 27557 527223 27591
rect 527189 17969 527223 18003
rect 532709 27557 532743 27591
rect 516149 9673 516183 9707
rect 568037 27557 568071 27591
rect 550649 19261 550683 19295
rect 550649 12325 550683 12359
rect 553409 19261 553443 19295
rect 532709 9673 532743 9707
rect 568037 17969 568071 18003
rect 569969 27557 570003 27591
rect 553409 9673 553443 9707
rect 569969 9673 570003 9707
rect 517897 9605 517931 9639
rect 144837 8653 144871 8687
rect 486525 7293 486559 7327
rect 144837 4845 144871 4879
rect 154589 4845 154623 4879
rect 154589 3893 154623 3927
rect 509157 3485 509191 3519
rect 511917 3485 511951 3519
rect 486525 3417 486559 3451
rect 499589 3417 499623 3451
rect 499589 3281 499623 3315
rect 512009 3417 512043 3451
rect 509157 3281 509191 3315
rect 519093 9605 519127 9639
rect 518909 3553 518943 3587
rect 518909 3417 518943 3451
rect 517897 561 517931 595
rect 545313 9605 545347 9639
rect 528477 3553 528511 3587
rect 528477 3417 528511 3451
rect 519093 561 519127 595
rect 545313 561 545347 595
rect 548901 9605 548935 9639
rect 548901 561 548935 595
rect 550097 9605 550131 9639
rect 559021 3485 559055 3519
rect 559021 3281 559055 3315
rect 550097 561 550131 595
<< metal1 >>
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 283282 698232 283288 698284
rect 283340 698272 283346 698284
rect 283926 698272 283932 698284
rect 283340 698244 283932 698272
rect 283340 698232 283346 698244
rect 283926 698232 283932 698244
rect 283984 698232 283990 698284
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 201494 697552 201500 697604
rect 201552 697592 201558 697604
rect 202782 697592 202788 697604
rect 201552 697564 202788 697592
rect 201552 697552 201558 697564
rect 202782 697552 202788 697564
rect 202840 697552 202846 697604
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 331214 697552 331220 697604
rect 331272 697592 331278 697604
rect 332502 697592 332508 697604
rect 331272 697564 332508 697592
rect 331272 697552 331278 697564
rect 332502 697552 332508 697564
rect 332560 697552 332566 697604
rect 567838 696940 567844 696992
rect 567896 696980 567902 696992
rect 580166 696980 580172 696992
rect 567896 696952 580172 696980
rect 567896 696940 567902 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 283098 694084 283104 694136
rect 283156 694124 283162 694136
rect 283282 694124 283288 694136
rect 283156 694096 283288 694124
rect 283156 694084 283162 694096
rect 283282 694084 283288 694096
rect 283340 694084 283346 694136
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 218054 692792 218060 692844
rect 218112 692832 218118 692844
rect 219066 692832 219072 692844
rect 218112 692804 219072 692832
rect 218112 692792 218118 692804
rect 219066 692792 219072 692804
rect 219124 692792 219130 692844
rect 234614 692792 234620 692844
rect 234672 692832 234678 692844
rect 235258 692832 235264 692844
rect 234672 692804 235264 692832
rect 234672 692792 234678 692804
rect 235258 692792 235264 692804
rect 235316 692792 235322 692844
rect 347774 692792 347780 692844
rect 347832 692832 347838 692844
rect 348878 692832 348884 692844
rect 347832 692804 348884 692832
rect 347832 692792 347838 692804
rect 348878 692792 348884 692804
rect 348936 692792 348942 692844
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 283098 692724 283104 692776
rect 283156 692764 283162 692776
rect 283282 692764 283288 692776
rect 283156 692736 283288 692764
rect 283156 692724 283162 692736
rect 283282 692724 283288 692736
rect 283340 692724 283346 692776
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 542538 692724 542544 692776
rect 542596 692764 542602 692776
rect 542722 692764 542728 692776
rect 542596 692736 542728 692764
rect 542596 692724 542602 692736
rect 542722 692724 542728 692736
rect 542780 692724 542786 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 299474 684428 299480 684480
rect 299532 684468 299538 684480
rect 300118 684468 300124 684480
rect 299532 684440 300124 684468
rect 299532 684428 299538 684440
rect 300118 684428 300124 684440
rect 300176 684428 300182 684480
rect 429194 684428 429200 684480
rect 429252 684468 429258 684480
rect 429838 684468 429844 684480
rect 429252 684440 429844 684468
rect 429252 684428 429258 684440
rect 429838 684428 429844 684440
rect 429896 684428 429902 684480
rect 558914 684428 558920 684480
rect 558972 684468 558978 684480
rect 559650 684468 559656 684480
rect 558972 684440 559656 684468
rect 558972 684428 558978 684440
rect 559650 684428 559656 684440
rect 559708 684428 559714 684480
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 282914 683068 282920 683120
rect 282972 683108 282978 683120
rect 283285 683111 283343 683117
rect 283285 683108 283297 683111
rect 282972 683080 283297 683108
rect 282972 683068 282978 683080
rect 283285 683077 283297 683080
rect 283331 683077 283343 683111
rect 283285 683071 283343 683077
rect 299474 683068 299480 683120
rect 299532 683108 299538 683120
rect 299845 683111 299903 683117
rect 299845 683108 299857 683111
rect 299532 683080 299857 683108
rect 299532 683068 299538 683080
rect 299845 683077 299857 683080
rect 299891 683077 299903 683111
rect 299845 683071 299903 683077
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 429194 683068 429200 683120
rect 429252 683108 429258 683120
rect 429565 683111 429623 683117
rect 429565 683108 429577 683111
rect 429252 683080 429577 683108
rect 429252 683068 429258 683080
rect 429565 683077 429577 683080
rect 429611 683077 429623 683111
rect 429565 683071 429623 683077
rect 542354 683068 542360 683120
rect 542412 683108 542418 683120
rect 542725 683111 542783 683117
rect 542725 683108 542737 683111
rect 542412 683080 542737 683108
rect 542412 683068 542418 683080
rect 542725 683077 542737 683080
rect 542771 683077 542783 683111
rect 542725 683071 542783 683077
rect 558914 683068 558920 683120
rect 558972 683108 558978 683120
rect 559285 683111 559343 683117
rect 559285 683108 559297 683111
rect 558972 683080 559297 683108
rect 558972 683068 558978 683080
rect 559285 683077 559297 683080
rect 559331 683077 559343 683111
rect 559285 683071 559343 683077
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 8938 681748 8944 681760
rect 3568 681720 8944 681748
rect 3568 681708 3574 681720
rect 8938 681708 8944 681720
rect 8996 681708 9002 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 218054 673480 218060 673532
rect 218112 673520 218118 673532
rect 218238 673520 218244 673532
rect 218112 673492 218244 673520
rect 218112 673480 218118 673492
rect 218238 673480 218244 673492
rect 218296 673480 218302 673532
rect 234614 673480 234620 673532
rect 234672 673520 234678 673532
rect 234798 673520 234804 673532
rect 234672 673492 234804 673520
rect 234672 673480 234678 673492
rect 234798 673480 234804 673492
rect 234856 673480 234862 673532
rect 347774 673480 347780 673532
rect 347832 673520 347838 673532
rect 347958 673520 347964 673532
rect 347832 673492 347964 673520
rect 347832 673480 347838 673492
rect 347958 673480 347964 673492
rect 348016 673480 348022 673532
rect 364334 673480 364340 673532
rect 364392 673520 364398 673532
rect 364518 673520 364524 673532
rect 364392 673492 364524 673520
rect 364392 673480 364398 673492
rect 364518 673480 364524 673492
rect 364576 673480 364582 673532
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 494054 673480 494060 673532
rect 494112 673520 494118 673532
rect 494238 673520 494244 673532
rect 494112 673492 494244 673520
rect 494112 673480 494118 673492
rect 494238 673480 494244 673492
rect 494296 673480 494302 673532
rect 558178 673480 558184 673532
rect 558236 673520 558242 673532
rect 580166 673520 580172 673532
rect 558236 673492 580172 673520
rect 558236 673480 558242 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 283285 666587 283343 666593
rect 283285 666553 283297 666587
rect 283331 666584 283343 666587
rect 283374 666584 283380 666596
rect 283331 666556 283380 666584
rect 283331 666553 283343 666556
rect 283285 666547 283343 666553
rect 283374 666544 283380 666556
rect 283432 666544 283438 666596
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 218054 654100 218060 654152
rect 218112 654140 218118 654152
rect 218238 654140 218244 654152
rect 218112 654112 218244 654140
rect 218112 654100 218118 654112
rect 218238 654100 218244 654112
rect 218296 654100 218302 654152
rect 234614 654100 234620 654152
rect 234672 654140 234678 654152
rect 234798 654140 234804 654152
rect 234672 654112 234804 654140
rect 234672 654100 234678 654112
rect 234798 654100 234804 654112
rect 234856 654100 234862 654152
rect 347774 654100 347780 654152
rect 347832 654140 347838 654152
rect 347958 654140 347964 654152
rect 347832 654112 347964 654140
rect 347832 654100 347838 654112
rect 347958 654100 347964 654112
rect 348016 654100 348022 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 14458 652780 14464 652792
rect 3108 652752 14464 652780
rect 3108 652740 3114 652752
rect 14458 652740 14464 652752
rect 14516 652740 14522 652792
rect 566458 650020 566464 650072
rect 566516 650060 566522 650072
rect 580166 650060 580172 650072
rect 566516 650032 580172 650060
rect 566516 650020 566522 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 283098 647232 283104 647284
rect 283156 647272 283162 647284
rect 283190 647272 283196 647284
rect 283156 647244 283196 647272
rect 283156 647232 283162 647244
rect 283190 647232 283196 647244
rect 283248 647232 283254 647284
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 283098 640364 283104 640416
rect 283156 640404 283162 640416
rect 283190 640404 283196 640416
rect 283156 640376 283196 640404
rect 283156 640364 283162 640376
rect 283190 640364 283196 640376
rect 283248 640364 283254 640416
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 573358 638936 573364 638988
rect 573416 638976 573422 638988
rect 580166 638976 580172 638988
rect 573416 638948 580172 638976
rect 573416 638936 573422 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 72786 637508 72792 637560
rect 72844 637548 72850 637560
rect 72878 637548 72884 637560
rect 72844 637520 72884 637548
rect 72844 637508 72850 637520
rect 72878 637508 72884 637520
rect 72936 637508 72942 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 218054 634788 218060 634840
rect 218112 634828 218118 634840
rect 218238 634828 218244 634840
rect 218112 634800 218244 634828
rect 218112 634788 218118 634800
rect 218238 634788 218244 634800
rect 218296 634788 218302 634840
rect 234614 634788 234620 634840
rect 234672 634828 234678 634840
rect 234798 634828 234804 634840
rect 234672 634800 234804 634828
rect 234672 634788 234678 634800
rect 234798 634788 234804 634800
rect 234856 634788 234862 634840
rect 347774 634788 347780 634840
rect 347832 634828 347838 634840
rect 347958 634828 347964 634840
rect 347832 634800 347964 634828
rect 347832 634788 347838 634800
rect 347958 634788 347964 634800
rect 348016 634788 348022 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 283006 630640 283012 630692
rect 283064 630680 283070 630692
rect 283190 630680 283196 630692
rect 283064 630652 283196 630680
rect 283064 630640 283070 630652
rect 283190 630640 283196 630652
rect 283248 630640 283254 630692
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 556798 626560 556804 626612
rect 556856 626600 556862 626612
rect 580166 626600 580172 626612
rect 556856 626572 580172 626600
rect 556856 626560 556862 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 73062 626532 73068 626544
rect 73023 626504 73068 626532
rect 73062 626492 73068 626504
rect 73120 626492 73126 626544
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 29638 623812 29644 623824
rect 3292 623784 29644 623812
rect 3292 623772 3298 623784
rect 29638 623772 29644 623784
rect 29696 623772 29702 623824
rect 73062 616876 73068 616888
rect 73023 616848 73068 616876
rect 73062 616836 73068 616848
rect 73120 616836 73126 616888
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 218054 615476 218060 615528
rect 218112 615516 218118 615528
rect 218238 615516 218244 615528
rect 218112 615488 218244 615516
rect 218112 615476 218118 615488
rect 218238 615476 218244 615488
rect 218296 615476 218302 615528
rect 234614 615476 234620 615528
rect 234672 615516 234678 615528
rect 234798 615516 234804 615528
rect 234672 615488 234804 615516
rect 234672 615476 234678 615488
rect 234798 615476 234804 615488
rect 234856 615476 234862 615528
rect 347774 615476 347780 615528
rect 347832 615516 347838 615528
rect 347958 615516 347964 615528
rect 347832 615488 347964 615516
rect 347832 615476 347838 615488
rect 347958 615476 347964 615488
rect 348016 615476 348022 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 477494 615476 477500 615528
rect 477552 615516 477558 615528
rect 477678 615516 477684 615528
rect 477552 615488 477684 615516
rect 477552 615476 477558 615488
rect 477678 615476 477684 615488
rect 477736 615476 477742 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 73062 611436 73068 611448
rect 72896 611408 73068 611436
rect 72896 611312 72924 611408
rect 73062 611396 73068 611408
rect 73120 611396 73126 611448
rect 283006 611328 283012 611380
rect 283064 611368 283070 611380
rect 283190 611368 283196 611380
rect 283064 611340 283196 611368
rect 283064 611328 283070 611340
rect 283190 611328 283196 611340
rect 283248 611328 283254 611380
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 72878 611260 72884 611312
rect 72936 611260 72942 611312
rect 283098 608580 283104 608592
rect 283059 608552 283104 608580
rect 283098 608540 283104 608552
rect 283156 608540 283162 608592
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 412818 608580 412824 608592
rect 412779 608552 412824 608580
rect 412818 608540 412824 608552
rect 412876 608540 412882 608592
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 542538 608580 542544 608592
rect 542499 608552 542544 608580
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 565078 603100 565084 603152
rect 565136 603140 565142 603152
rect 580166 603140 580172 603152
rect 565136 603112 580172 603140
rect 565136 603100 565142 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 283101 601715 283159 601721
rect 283101 601681 283113 601715
rect 283147 601712 283159 601715
rect 283282 601712 283288 601724
rect 283147 601684 283288 601712
rect 283147 601681 283159 601684
rect 283101 601675 283159 601681
rect 283282 601672 283288 601684
rect 283340 601672 283346 601724
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 412821 601715 412879 601721
rect 412821 601681 412833 601715
rect 412867 601712 412879 601715
rect 413002 601712 413008 601724
rect 412867 601684 413008 601712
rect 412867 601681 412879 601684
rect 412821 601675 412879 601681
rect 413002 601672 413008 601684
rect 413060 601672 413066 601724
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 542541 601715 542599 601721
rect 542541 601681 542553 601715
rect 542587 601712 542599 601715
rect 542722 601712 542728 601724
rect 542587 601684 542728 601712
rect 542587 601681 542599 601684
rect 542541 601675 542599 601681
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 72970 601536 72976 601588
rect 73028 601576 73034 601588
rect 73154 601576 73160 601588
rect 73028 601548 73160 601576
rect 73028 601536 73034 601548
rect 73154 601536 73160 601548
rect 73212 601536 73218 601588
rect 72881 598927 72939 598933
rect 72881 598893 72893 598927
rect 72927 598924 72939 598927
rect 72970 598924 72976 598936
rect 72927 598896 72976 598924
rect 72927 598893 72939 598896
rect 72881 598887 72939 598893
rect 72970 598884 72976 598896
rect 73028 598884 73034 598936
rect 283282 598924 283288 598936
rect 283243 598896 283288 598924
rect 283282 598884 283288 598896
rect 283340 598884 283346 598936
rect 299842 598924 299848 598936
rect 299803 598896 299848 598924
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 413002 598924 413008 598936
rect 412963 598896 413008 598924
rect 413002 598884 413008 598896
rect 413060 598884 413066 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 542722 598924 542728 598936
rect 542683 598896 542728 598924
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 137738 596164 137744 596216
rect 137796 596204 137802 596216
rect 137922 596204 137928 596216
rect 137796 596176 137928 596204
rect 137796 596164 137802 596176
rect 137922 596164 137928 596176
rect 137980 596164 137986 596216
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 218054 596164 218060 596216
rect 218112 596204 218118 596216
rect 218238 596204 218244 596216
rect 218112 596176 218244 596204
rect 218112 596164 218118 596176
rect 218238 596164 218244 596176
rect 218296 596164 218302 596216
rect 234614 596164 234620 596216
rect 234672 596204 234678 596216
rect 234798 596204 234804 596216
rect 234672 596176 234804 596204
rect 234672 596164 234678 596176
rect 234798 596164 234804 596176
rect 234856 596164 234862 596216
rect 347774 596164 347780 596216
rect 347832 596204 347838 596216
rect 347958 596204 347964 596216
rect 347832 596176 347964 596204
rect 347832 596164 347838 596176
rect 347958 596164 347964 596176
rect 348016 596164 348022 596216
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 477494 596164 477500 596216
rect 477552 596204 477558 596216
rect 477678 596204 477684 596216
rect 477552 596176 477684 596204
rect 477552 596164 477558 596176
rect 477678 596164 477684 596176
rect 477736 596164 477742 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 44818 594844 44824 594856
rect 3384 594816 44824 594844
rect 3384 594804 3390 594816
rect 44818 594804 44824 594816
rect 44876 594804 44882 594856
rect 570598 592016 570604 592068
rect 570656 592056 570662 592068
rect 580166 592056 580172 592068
rect 570656 592028 580172 592056
rect 570656 592016 570662 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 72878 589336 72884 589348
rect 72839 589308 72884 589336
rect 72878 589296 72884 589308
rect 72936 589296 72942 589348
rect 283285 589339 283343 589345
rect 283285 589305 283297 589339
rect 283331 589336 283343 589339
rect 283374 589336 283380 589348
rect 283331 589308 283380 589336
rect 283331 589305 283343 589308
rect 283285 589299 283343 589305
rect 283374 589296 283380 589308
rect 283432 589296 283438 589348
rect 299845 589339 299903 589345
rect 299845 589305 299857 589339
rect 299891 589336 299903 589339
rect 299934 589336 299940 589348
rect 299891 589308 299940 589336
rect 299891 589305 299903 589308
rect 299845 589299 299903 589305
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 413005 589339 413063 589345
rect 413005 589305 413017 589339
rect 413051 589336 413063 589339
rect 413094 589336 413100 589348
rect 413051 589308 413100 589336
rect 413051 589305 413063 589308
rect 413005 589299 413063 589305
rect 413094 589296 413100 589308
rect 413152 589296 413158 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 542725 589339 542783 589345
rect 542725 589305 542737 589339
rect 542771 589336 542783 589339
rect 542814 589336 542820 589348
rect 542771 589308 542820 589336
rect 542771 589305 542783 589308
rect 542725 589299 542783 589305
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 8018 589268 8024 589280
rect 7979 589240 8024 589268
rect 8018 589228 8024 589240
rect 8076 589228 8082 589280
rect 137738 589268 137744 589280
rect 137699 589240 137744 589268
rect 137738 589228 137744 589240
rect 137796 589228 137802 589280
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 218057 589271 218115 589277
rect 218057 589237 218069 589271
rect 218103 589268 218115 589271
rect 218146 589268 218152 589280
rect 218103 589240 218152 589268
rect 218103 589237 218115 589240
rect 218057 589231 218115 589237
rect 218146 589228 218152 589240
rect 218204 589228 218210 589280
rect 234617 589271 234675 589277
rect 234617 589237 234629 589271
rect 234663 589268 234675 589271
rect 234706 589268 234712 589280
rect 234663 589240 234712 589268
rect 234663 589237 234675 589240
rect 234617 589231 234675 589237
rect 234706 589228 234712 589240
rect 234764 589228 234770 589280
rect 347777 589271 347835 589277
rect 347777 589237 347789 589271
rect 347823 589268 347835 589271
rect 347866 589268 347872 589280
rect 347823 589240 347872 589268
rect 347823 589237 347835 589240
rect 347777 589231 347835 589237
rect 347866 589228 347872 589240
rect 347924 589228 347930 589280
rect 364337 589271 364395 589277
rect 364337 589237 364349 589271
rect 364383 589268 364395 589271
rect 364426 589268 364432 589280
rect 364383 589240 364432 589268
rect 364383 589237 364395 589240
rect 364337 589231 364395 589237
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 477497 589271 477555 589277
rect 477497 589237 477509 589271
rect 477543 589268 477555 589271
rect 477586 589268 477592 589280
rect 477543 589240 477592 589268
rect 477543 589237 477555 589240
rect 477497 589231 477555 589237
rect 477586 589228 477592 589240
rect 477644 589228 477650 589280
rect 494057 589271 494115 589277
rect 494057 589237 494069 589271
rect 494103 589268 494115 589271
rect 494146 589268 494152 589280
rect 494103 589240 494152 589268
rect 494103 589237 494115 589240
rect 494057 589231 494115 589237
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 283374 582468 283380 582480
rect 283300 582440 283380 582468
rect 72694 582360 72700 582412
rect 72752 582400 72758 582412
rect 72878 582400 72884 582412
rect 72752 582372 72884 582400
rect 72752 582360 72758 582372
rect 72878 582360 72884 582372
rect 72936 582360 72942 582412
rect 283300 582344 283328 582440
rect 283374 582428 283380 582440
rect 283432 582428 283438 582480
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 413094 582468 413100 582480
rect 413020 582440 413100 582468
rect 413020 582344 413048 582440
rect 413094 582428 413100 582440
rect 413152 582428 413158 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 283282 582292 283288 582344
rect 283340 582292 283346 582344
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 413002 582292 413008 582344
rect 413060 582292 413066 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 8018 579748 8024 579760
rect 7979 579720 8024 579748
rect 8018 579708 8024 579720
rect 8076 579708 8082 579760
rect 137738 579748 137744 579760
rect 137699 579720 137744 579748
rect 137738 579708 137744 579720
rect 137796 579708 137802 579760
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 218054 579680 218060 579692
rect 218015 579652 218060 579680
rect 218054 579640 218060 579652
rect 218112 579640 218118 579692
rect 234614 579680 234620 579692
rect 234575 579652 234620 579680
rect 234614 579640 234620 579652
rect 234672 579640 234678 579692
rect 347774 579640 347780 579692
rect 347832 579680 347838 579692
rect 364334 579680 364340 579692
rect 347832 579652 347877 579680
rect 364295 579652 364340 579680
rect 347832 579640 347838 579652
rect 364334 579640 364340 579652
rect 364392 579640 364398 579692
rect 477494 579680 477500 579692
rect 477455 579652 477500 579680
rect 477494 579640 477500 579652
rect 477552 579640 477558 579692
rect 494054 579680 494060 579692
rect 494015 579652 494060 579680
rect 494054 579640 494060 579652
rect 494112 579640 494118 579692
rect 555418 579640 555424 579692
rect 555476 579680 555482 579692
rect 580166 579680 580172 579692
rect 555476 579652 580172 579680
rect 555476 579640 555482 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 7926 579572 7932 579624
rect 7984 579612 7990 579624
rect 8110 579612 8116 579624
rect 7984 579584 8116 579612
rect 7984 579572 7990 579584
rect 8110 579572 8116 579584
rect 8168 579572 8174 579624
rect 72605 579615 72663 579621
rect 72605 579581 72617 579615
rect 72651 579612 72663 579615
rect 72694 579612 72700 579624
rect 72651 579584 72700 579612
rect 72651 579581 72663 579584
rect 72605 579575 72663 579581
rect 72694 579572 72700 579584
rect 72752 579572 72758 579624
rect 137557 579615 137615 579621
rect 137557 579581 137569 579615
rect 137603 579612 137615 579615
rect 137646 579612 137652 579624
rect 137603 579584 137652 579612
rect 137603 579581 137615 579584
rect 137557 579575 137615 579581
rect 137646 579572 137652 579584
rect 137704 579572 137710 579624
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 72602 569956 72608 569968
rect 72563 569928 72608 569956
rect 72602 569916 72608 569928
rect 72660 569916 72666 569968
rect 137554 569956 137560 569968
rect 137515 569928 137560 569956
rect 137554 569916 137560 569928
rect 137612 569916 137618 569968
rect 218146 569888 218152 569900
rect 218107 569860 218152 569888
rect 218146 569848 218152 569860
rect 218204 569848 218210 569900
rect 234706 569888 234712 569900
rect 234667 569860 234712 569888
rect 234706 569848 234712 569860
rect 234764 569848 234770 569900
rect 347866 569888 347872 569900
rect 347827 569860 347872 569888
rect 347866 569848 347872 569860
rect 347924 569848 347930 569900
rect 364426 569888 364432 569900
rect 364387 569860 364432 569888
rect 364426 569848 364432 569860
rect 364484 569848 364490 569900
rect 477586 569888 477592 569900
rect 477547 569860 477592 569888
rect 477586 569848 477592 569860
rect 477644 569848 477650 569900
rect 494146 569888 494152 569900
rect 494107 569860 494152 569888
rect 494146 569848 494152 569860
rect 494204 569848 494210 569900
rect 4062 567196 4068 567248
rect 4120 567236 4126 567248
rect 13078 567236 13084 567248
rect 4120 567208 13084 567236
rect 4120 567196 4126 567208
rect 13078 567196 13084 567208
rect 13136 567196 13142 567248
rect 283006 563116 283012 563168
rect 283064 563116 283070 563168
rect 412726 563116 412732 563168
rect 412784 563116 412790 563168
rect 429286 563116 429292 563168
rect 429344 563116 429350 563168
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 72602 563048 72608 563100
rect 72660 563048 72666 563100
rect 137554 563048 137560 563100
rect 137612 563048 137618 563100
rect 218149 563091 218207 563097
rect 218149 563057 218161 563091
rect 218195 563088 218207 563091
rect 218330 563088 218336 563100
rect 218195 563060 218336 563088
rect 218195 563057 218207 563060
rect 218149 563051 218207 563057
rect 218330 563048 218336 563060
rect 218388 563048 218394 563100
rect 234709 563091 234767 563097
rect 234709 563057 234721 563091
rect 234755 563088 234767 563091
rect 234890 563088 234896 563100
rect 234755 563060 234896 563088
rect 234755 563057 234767 563060
rect 234709 563051 234767 563057
rect 234890 563048 234896 563060
rect 234948 563048 234954 563100
rect 7926 562912 7932 562964
rect 7984 562952 7990 562964
rect 8110 562952 8116 562964
rect 7984 562924 8116 562952
rect 7984 562912 7990 562924
rect 8110 562912 8116 562924
rect 8168 562912 8174 562964
rect 72620 562952 72648 563048
rect 72694 562952 72700 562964
rect 72620 562924 72700 562952
rect 72694 562912 72700 562924
rect 72752 562912 72758 562964
rect 137572 562952 137600 563048
rect 283024 563032 283052 563116
rect 347869 563091 347927 563097
rect 347869 563057 347881 563091
rect 347915 563088 347927 563091
rect 348050 563088 348056 563100
rect 347915 563060 348056 563088
rect 347915 563057 347927 563060
rect 347869 563051 347927 563057
rect 348050 563048 348056 563060
rect 348108 563048 348114 563100
rect 364429 563091 364487 563097
rect 364429 563057 364441 563091
rect 364475 563088 364487 563091
rect 364610 563088 364616 563100
rect 364475 563060 364616 563088
rect 364475 563057 364487 563060
rect 364429 563051 364487 563057
rect 364610 563048 364616 563060
rect 364668 563048 364674 563100
rect 412744 563032 412772 563116
rect 429304 563032 429332 563116
rect 477589 563091 477647 563097
rect 477589 563057 477601 563091
rect 477635 563088 477647 563091
rect 477770 563088 477776 563100
rect 477635 563060 477776 563088
rect 477635 563057 477647 563060
rect 477589 563051 477647 563057
rect 477770 563048 477776 563060
rect 477828 563048 477834 563100
rect 494149 563091 494207 563097
rect 494149 563057 494161 563091
rect 494195 563088 494207 563091
rect 494330 563088 494336 563100
rect 494195 563060 494336 563088
rect 494195 563057 494207 563060
rect 494149 563051 494207 563057
rect 494330 563048 494336 563060
rect 494388 563048 494394 563100
rect 542464 563032 542492 563116
rect 559024 563032 559052 563116
rect 283006 562980 283012 563032
rect 283064 562980 283070 563032
rect 412726 562980 412732 563032
rect 412784 562980 412790 563032
rect 429286 562980 429292 563032
rect 429344 562980 429350 563032
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 137646 562952 137652 562964
rect 137572 562924 137652 562952
rect 137646 562912 137652 562924
rect 137704 562912 137710 562964
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 137646 560232 137652 560244
rect 137607 560204 137652 560232
rect 137646 560192 137652 560204
rect 137704 560192 137710 560244
rect 283006 560232 283012 560244
rect 282967 560204 283012 560232
rect 283006 560192 283012 560204
rect 283064 560192 283070 560244
rect 412726 560232 412732 560244
rect 412687 560204 412732 560232
rect 412726 560192 412732 560204
rect 412784 560192 412790 560244
rect 429286 560232 429292 560244
rect 429247 560204 429292 560232
rect 429286 560192 429292 560204
rect 429344 560192 429350 560244
rect 542446 560232 542452 560244
rect 542407 560204 542452 560232
rect 542446 560192 542452 560204
rect 542504 560192 542510 560244
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 563698 556180 563704 556232
rect 563756 556220 563762 556232
rect 580166 556220 580172 556232
rect 563756 556192 580172 556220
rect 563756 556180 563762 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 72602 553432 72608 553444
rect 72563 553404 72608 553432
rect 72602 553392 72608 553404
rect 72660 553392 72666 553444
rect 72602 550644 72608 550656
rect 72563 550616 72608 550644
rect 72602 550604 72608 550616
rect 72660 550604 72666 550656
rect 137649 550647 137707 550653
rect 137649 550613 137661 550647
rect 137695 550644 137707 550647
rect 137830 550644 137836 550656
rect 137695 550616 137836 550644
rect 137695 550613 137707 550616
rect 137649 550607 137707 550613
rect 137830 550604 137836 550616
rect 137888 550604 137894 550656
rect 218146 550604 218152 550656
rect 218204 550644 218210 550656
rect 218422 550644 218428 550656
rect 218204 550616 218428 550644
rect 218204 550604 218210 550616
rect 218422 550604 218428 550616
rect 218480 550604 218486 550656
rect 234706 550604 234712 550656
rect 234764 550644 234770 550656
rect 234982 550644 234988 550656
rect 234764 550616 234988 550644
rect 234764 550604 234770 550616
rect 234982 550604 234988 550616
rect 235040 550604 235046 550656
rect 283009 550647 283067 550653
rect 283009 550613 283021 550647
rect 283055 550644 283067 550647
rect 283190 550644 283196 550656
rect 283055 550616 283196 550644
rect 283055 550613 283067 550616
rect 283009 550607 283067 550613
rect 283190 550604 283196 550616
rect 283248 550604 283254 550656
rect 299474 550604 299480 550656
rect 299532 550644 299538 550656
rect 299750 550644 299756 550656
rect 299532 550616 299756 550644
rect 299532 550604 299538 550616
rect 299750 550604 299756 550616
rect 299808 550604 299814 550656
rect 347866 550604 347872 550656
rect 347924 550644 347930 550656
rect 348142 550644 348148 550656
rect 347924 550616 348148 550644
rect 347924 550604 347930 550616
rect 348142 550604 348148 550616
rect 348200 550604 348206 550656
rect 364426 550604 364432 550656
rect 364484 550644 364490 550656
rect 364702 550644 364708 550656
rect 364484 550616 364708 550644
rect 364484 550604 364490 550616
rect 364702 550604 364708 550616
rect 364760 550604 364766 550656
rect 412729 550647 412787 550653
rect 412729 550613 412741 550647
rect 412775 550644 412787 550647
rect 412910 550644 412916 550656
rect 412775 550616 412916 550644
rect 412775 550613 412787 550616
rect 412729 550607 412787 550613
rect 412910 550604 412916 550616
rect 412968 550604 412974 550656
rect 429289 550647 429347 550653
rect 429289 550613 429301 550647
rect 429335 550644 429347 550647
rect 429470 550644 429476 550656
rect 429335 550616 429476 550644
rect 429335 550613 429347 550616
rect 429289 550607 429347 550613
rect 429470 550604 429476 550616
rect 429528 550604 429534 550656
rect 477586 550604 477592 550656
rect 477644 550644 477650 550656
rect 477862 550644 477868 550656
rect 477644 550616 477868 550644
rect 477644 550604 477650 550616
rect 477862 550604 477868 550616
rect 477920 550604 477926 550656
rect 494146 550604 494152 550656
rect 494204 550644 494210 550656
rect 494422 550644 494428 550656
rect 494204 550616 494428 550644
rect 494204 550604 494210 550616
rect 494422 550604 494428 550616
rect 494480 550604 494486 550656
rect 542449 550647 542507 550653
rect 542449 550613 542461 550647
rect 542495 550644 542507 550647
rect 542630 550644 542636 550656
rect 542495 550616 542636 550644
rect 542495 550613 542507 550616
rect 542449 550607 542507 550613
rect 542630 550604 542636 550616
rect 542688 550604 542694 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559190 550644 559196 550656
rect 559055 550616 559196 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559190 550604 559196 550616
rect 559248 550604 559254 550656
rect 8018 550576 8024 550588
rect 7979 550548 8024 550576
rect 8018 550536 8024 550548
rect 8076 550536 8082 550588
rect 552658 545096 552664 545148
rect 552716 545136 552722 545148
rect 580166 545136 580172 545148
rect 552716 545108 580172 545136
rect 552716 545096 552722 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 218422 543844 218428 543856
rect 218348 543816 218428 543844
rect 72602 543736 72608 543788
rect 72660 543736 72666 543788
rect 72620 543640 72648 543736
rect 218348 543720 218376 543816
rect 218422 543804 218428 543816
rect 218480 543804 218486 543856
rect 234982 543844 234988 543856
rect 234908 543816 234988 543844
rect 234908 543720 234936 543816
rect 234982 543804 234988 543816
rect 235040 543804 235046 543856
rect 348142 543844 348148 543856
rect 348068 543816 348148 543844
rect 299474 543736 299480 543788
rect 299532 543736 299538 543788
rect 218330 543668 218336 543720
rect 218388 543668 218394 543720
rect 234890 543668 234896 543720
rect 234948 543668 234954 543720
rect 72694 543640 72700 543652
rect 72620 543612 72700 543640
rect 72694 543600 72700 543612
rect 72752 543600 72758 543652
rect 137646 543600 137652 543652
rect 137704 543640 137710 543652
rect 137830 543640 137836 543652
rect 137704 543612 137836 543640
rect 137704 543600 137710 543612
rect 137830 543600 137836 543612
rect 137888 543600 137894 543652
rect 283006 543600 283012 543652
rect 283064 543640 283070 543652
rect 283190 543640 283196 543652
rect 283064 543612 283196 543640
rect 283064 543600 283070 543612
rect 283190 543600 283196 543612
rect 283248 543600 283254 543652
rect 299492 543640 299520 543736
rect 348068 543720 348096 543816
rect 348142 543804 348148 543816
rect 348200 543804 348206 543856
rect 364702 543844 364708 543856
rect 364628 543816 364708 543844
rect 364628 543720 364656 543816
rect 364702 543804 364708 543816
rect 364760 543804 364766 543856
rect 477862 543844 477868 543856
rect 477788 543816 477868 543844
rect 477788 543720 477816 543816
rect 477862 543804 477868 543816
rect 477920 543804 477926 543856
rect 494422 543844 494428 543856
rect 494348 543816 494428 543844
rect 494348 543720 494376 543816
rect 494422 543804 494428 543816
rect 494480 543804 494486 543856
rect 348050 543668 348056 543720
rect 348108 543668 348114 543720
rect 364610 543668 364616 543720
rect 364668 543668 364674 543720
rect 477770 543668 477776 543720
rect 477828 543668 477834 543720
rect 494330 543668 494336 543720
rect 494388 543668 494394 543720
rect 299566 543640 299572 543652
rect 299492 543612 299572 543640
rect 299566 543600 299572 543612
rect 299624 543600 299630 543652
rect 412726 543600 412732 543652
rect 412784 543640 412790 543652
rect 412910 543640 412916 543652
rect 412784 543612 412916 543640
rect 412784 543600 412790 543612
rect 412910 543600 412916 543612
rect 412968 543600 412974 543652
rect 429286 543600 429292 543652
rect 429344 543640 429350 543652
rect 429470 543640 429476 543652
rect 429344 543612 429476 543640
rect 429344 543600 429350 543612
rect 429470 543600 429476 543612
rect 429528 543600 429534 543652
rect 542446 543600 542452 543652
rect 542504 543640 542510 543652
rect 542630 543640 542636 543652
rect 542504 543612 542636 543640
rect 542504 543600 542510 543612
rect 542630 543600 542636 543612
rect 542688 543600 542694 543652
rect 559006 543600 559012 543652
rect 559064 543640 559070 543652
rect 559190 543640 559196 543652
rect 559064 543612 559196 543640
rect 559064 543600 559070 543612
rect 559190 543600 559196 543612
rect 559248 543600 559254 543652
rect 8021 540991 8079 540997
rect 8021 540957 8033 540991
rect 8067 540988 8079 540991
rect 8202 540988 8208 541000
rect 8067 540960 8208 540988
rect 8067 540957 8079 540960
rect 8021 540951 8079 540957
rect 8202 540948 8208 540960
rect 8260 540948 8266 541000
rect 4062 538228 4068 538280
rect 4120 538268 4126 538280
rect 17218 538268 17224 538280
rect 4120 538240 17224 538268
rect 4120 538228 4126 538240
rect 17218 538228 17224 538240
rect 17276 538228 17282 538280
rect 72602 534120 72608 534132
rect 72563 534092 72608 534120
rect 72602 534080 72608 534092
rect 72660 534080 72666 534132
rect 137646 534012 137652 534064
rect 137704 534052 137710 534064
rect 137830 534052 137836 534064
rect 137704 534024 137836 534052
rect 137704 534012 137710 534024
rect 137830 534012 137836 534024
rect 137888 534012 137894 534064
rect 283006 534012 283012 534064
rect 283064 534052 283070 534064
rect 283190 534052 283196 534064
rect 283064 534024 283196 534052
rect 283064 534012 283070 534024
rect 283190 534012 283196 534024
rect 283248 534012 283254 534064
rect 299566 534012 299572 534064
rect 299624 534052 299630 534064
rect 299750 534052 299756 534064
rect 299624 534024 299756 534052
rect 299624 534012 299630 534024
rect 299750 534012 299756 534024
rect 299808 534012 299814 534064
rect 412726 534012 412732 534064
rect 412784 534052 412790 534064
rect 412910 534052 412916 534064
rect 412784 534024 412916 534052
rect 412784 534012 412790 534024
rect 412910 534012 412916 534024
rect 412968 534012 412974 534064
rect 429286 534012 429292 534064
rect 429344 534052 429350 534064
rect 429470 534052 429476 534064
rect 429344 534024 429476 534052
rect 429344 534012 429350 534024
rect 429470 534012 429476 534024
rect 429528 534012 429534 534064
rect 542446 534012 542452 534064
rect 542504 534052 542510 534064
rect 542630 534052 542636 534064
rect 542504 534024 542636 534052
rect 542504 534012 542510 534024
rect 542630 534012 542636 534024
rect 542688 534012 542694 534064
rect 559006 534012 559012 534064
rect 559064 534052 559070 534064
rect 559190 534052 559196 534064
rect 559064 534024 559196 534052
rect 559064 534012 559070 534024
rect 559190 534012 559196 534024
rect 559248 534012 559254 534064
rect 72602 531332 72608 531344
rect 72563 531304 72608 531332
rect 72602 531292 72608 531304
rect 72660 531292 72666 531344
rect 218146 531292 218152 531344
rect 218204 531332 218210 531344
rect 218422 531332 218428 531344
rect 218204 531304 218428 531332
rect 218204 531292 218210 531304
rect 218422 531292 218428 531304
rect 218480 531292 218486 531344
rect 234706 531292 234712 531344
rect 234764 531332 234770 531344
rect 234982 531332 234988 531344
rect 234764 531304 234988 531332
rect 234764 531292 234770 531304
rect 234982 531292 234988 531304
rect 235040 531292 235046 531344
rect 347866 531292 347872 531344
rect 347924 531332 347930 531344
rect 348142 531332 348148 531344
rect 347924 531304 348148 531332
rect 347924 531292 347930 531304
rect 348142 531292 348148 531304
rect 348200 531292 348206 531344
rect 364426 531292 364432 531344
rect 364484 531332 364490 531344
rect 364702 531332 364708 531344
rect 364484 531304 364708 531332
rect 364484 531292 364490 531304
rect 364702 531292 364708 531304
rect 364760 531292 364766 531344
rect 477586 531292 477592 531344
rect 477644 531332 477650 531344
rect 477862 531332 477868 531344
rect 477644 531304 477868 531332
rect 477644 531292 477650 531304
rect 477862 531292 477868 531304
rect 477920 531292 477926 531344
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 218422 524532 218428 524544
rect 218348 524504 218428 524532
rect 218348 524408 218376 524504
rect 218422 524492 218428 524504
rect 218480 524492 218486 524544
rect 234982 524532 234988 524544
rect 234908 524504 234988 524532
rect 234908 524408 234936 524504
rect 234982 524492 234988 524504
rect 235040 524492 235046 524544
rect 348142 524532 348148 524544
rect 348068 524504 348148 524532
rect 283190 524424 283196 524476
rect 283248 524424 283254 524476
rect 299750 524424 299756 524476
rect 299808 524424 299814 524476
rect 218330 524356 218336 524408
rect 218388 524356 218394 524408
rect 234890 524356 234896 524408
rect 234948 524356 234954 524408
rect 283208 524396 283236 524424
rect 283282 524396 283288 524408
rect 283208 524368 283288 524396
rect 283282 524356 283288 524368
rect 283340 524356 283346 524408
rect 299768 524396 299796 524424
rect 348068 524408 348096 524504
rect 348142 524492 348148 524504
rect 348200 524492 348206 524544
rect 364702 524532 364708 524544
rect 364628 524504 364708 524532
rect 364628 524408 364656 524504
rect 364702 524492 364708 524504
rect 364760 524492 364766 524544
rect 477862 524532 477868 524544
rect 477788 524504 477868 524532
rect 412910 524424 412916 524476
rect 412968 524424 412974 524476
rect 429470 524424 429476 524476
rect 429528 524424 429534 524476
rect 299842 524396 299848 524408
rect 299768 524368 299848 524396
rect 299842 524356 299848 524368
rect 299900 524356 299906 524408
rect 348050 524356 348056 524408
rect 348108 524356 348114 524408
rect 364610 524356 364616 524408
rect 364668 524356 364674 524408
rect 412928 524396 412956 524424
rect 413002 524396 413008 524408
rect 412928 524368 413008 524396
rect 413002 524356 413008 524368
rect 413060 524356 413066 524408
rect 429488 524396 429516 524424
rect 477788 524408 477816 524504
rect 477862 524492 477868 524504
rect 477920 524492 477926 524544
rect 494422 524532 494428 524544
rect 494348 524504 494428 524532
rect 494348 524408 494376 524504
rect 494422 524492 494428 524504
rect 494480 524492 494486 524544
rect 542630 524424 542636 524476
rect 542688 524424 542694 524476
rect 559190 524424 559196 524476
rect 559248 524424 559254 524476
rect 429562 524396 429568 524408
rect 429488 524368 429568 524396
rect 429562 524356 429568 524368
rect 429620 524356 429626 524408
rect 477770 524356 477776 524408
rect 477828 524356 477834 524408
rect 494330 524356 494336 524408
rect 494388 524356 494394 524408
rect 542648 524396 542676 524424
rect 542722 524396 542728 524408
rect 542648 524368 542728 524396
rect 542722 524356 542728 524368
rect 542780 524356 542786 524408
rect 559208 524396 559236 524424
rect 559282 524396 559288 524408
rect 559208 524368 559288 524396
rect 559282 524356 559288 524368
rect 559340 524356 559346 524408
rect 72694 524288 72700 524340
rect 72752 524328 72758 524340
rect 72878 524328 72884 524340
rect 72752 524300 72884 524328
rect 72752 524288 72758 524300
rect 72878 524288 72884 524300
rect 72936 524288 72942 524340
rect 8202 521636 8208 521688
rect 8260 521676 8266 521688
rect 8386 521676 8392 521688
rect 8260 521648 8392 521676
rect 8260 521636 8266 521648
rect 8386 521636 8392 521648
rect 8444 521636 8450 521688
rect 137922 521636 137928 521688
rect 137980 521676 137986 521688
rect 138106 521676 138112 521688
rect 137980 521648 138112 521676
rect 137980 521636 137986 521648
rect 138106 521636 138112 521648
rect 138164 521636 138170 521688
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 218146 511980 218152 512032
rect 218204 512020 218210 512032
rect 218422 512020 218428 512032
rect 218204 511992 218428 512020
rect 218204 511980 218210 511992
rect 218422 511980 218428 511992
rect 218480 511980 218486 512032
rect 234706 511980 234712 512032
rect 234764 512020 234770 512032
rect 234982 512020 234988 512032
rect 234764 511992 234988 512020
rect 234764 511980 234770 511992
rect 234982 511980 234988 511992
rect 235040 511980 235046 512032
rect 283098 511980 283104 512032
rect 283156 512020 283162 512032
rect 283374 512020 283380 512032
rect 283156 511992 283380 512020
rect 283156 511980 283162 511992
rect 283374 511980 283380 511992
rect 283432 511980 283438 512032
rect 299658 511980 299664 512032
rect 299716 512020 299722 512032
rect 299934 512020 299940 512032
rect 299716 511992 299940 512020
rect 299716 511980 299722 511992
rect 299934 511980 299940 511992
rect 299992 511980 299998 512032
rect 347866 511980 347872 512032
rect 347924 512020 347930 512032
rect 348142 512020 348148 512032
rect 347924 511992 348148 512020
rect 347924 511980 347930 511992
rect 348142 511980 348148 511992
rect 348200 511980 348206 512032
rect 364426 511980 364432 512032
rect 364484 512020 364490 512032
rect 364702 512020 364708 512032
rect 364484 511992 364708 512020
rect 364484 511980 364490 511992
rect 364702 511980 364708 511992
rect 364760 511980 364766 512032
rect 412818 511980 412824 512032
rect 412876 512020 412882 512032
rect 413094 512020 413100 512032
rect 412876 511992 413100 512020
rect 412876 511980 412882 511992
rect 413094 511980 413100 511992
rect 413152 511980 413158 512032
rect 429378 511980 429384 512032
rect 429436 512020 429442 512032
rect 429654 512020 429660 512032
rect 429436 511992 429660 512020
rect 429436 511980 429442 511992
rect 429654 511980 429660 511992
rect 429712 511980 429718 512032
rect 477586 511980 477592 512032
rect 477644 512020 477650 512032
rect 477862 512020 477868 512032
rect 477644 511992 477868 512020
rect 477644 511980 477650 511992
rect 477862 511980 477868 511992
rect 477920 511980 477926 512032
rect 494146 511980 494152 512032
rect 494204 512020 494210 512032
rect 494422 512020 494428 512032
rect 494204 511992 494428 512020
rect 494204 511980 494210 511992
rect 494422 511980 494428 511992
rect 494480 511980 494486 512032
rect 542538 511980 542544 512032
rect 542596 512020 542602 512032
rect 542814 512020 542820 512032
rect 542596 511992 542820 512020
rect 542596 511980 542602 511992
rect 542814 511980 542820 511992
rect 542872 511980 542878 512032
rect 559098 511980 559104 512032
rect 559156 512020 559162 512032
rect 559374 512020 559380 512032
rect 559156 511992 559380 512020
rect 559156 511980 559162 511992
rect 559374 511980 559380 511992
rect 559432 511980 559438 512032
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 3878 509260 3884 509312
rect 3936 509300 3942 509312
rect 39298 509300 39304 509312
rect 3936 509272 39304 509300
rect 3936 509260 3942 509272
rect 39298 509260 39304 509272
rect 39356 509260 39362 509312
rect 551278 509260 551284 509312
rect 551336 509300 551342 509312
rect 580166 509300 580172 509312
rect 551336 509272 580172 509300
rect 551336 509260 551342 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 8202 502324 8208 502376
rect 8260 502364 8266 502376
rect 8386 502364 8392 502376
rect 8260 502336 8392 502364
rect 8260 502324 8266 502336
rect 8386 502324 8392 502336
rect 8444 502324 8450 502376
rect 72602 502324 72608 502376
rect 72660 502364 72666 502376
rect 73062 502364 73068 502376
rect 72660 502336 73068 502364
rect 72660 502324 72666 502336
rect 73062 502324 73068 502336
rect 73120 502324 73126 502376
rect 137922 502324 137928 502376
rect 137980 502364 137986 502376
rect 138106 502364 138112 502376
rect 137980 502336 138112 502364
rect 137980 502324 137986 502336
rect 138106 502324 138112 502336
rect 138164 502324 138170 502376
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 218238 502324 218244 502376
rect 218296 502364 218302 502376
rect 218422 502364 218428 502376
rect 218296 502336 218428 502364
rect 218296 502324 218302 502336
rect 218422 502324 218428 502336
rect 218480 502324 218486 502376
rect 234798 502324 234804 502376
rect 234856 502364 234862 502376
rect 234982 502364 234988 502376
rect 234856 502336 234988 502364
rect 234856 502324 234862 502336
rect 234982 502324 234988 502336
rect 235040 502324 235046 502376
rect 283190 502324 283196 502376
rect 283248 502364 283254 502376
rect 283374 502364 283380 502376
rect 283248 502336 283380 502364
rect 283248 502324 283254 502336
rect 283374 502324 283380 502336
rect 283432 502324 283438 502376
rect 299750 502324 299756 502376
rect 299808 502364 299814 502376
rect 299934 502364 299940 502376
rect 299808 502336 299940 502364
rect 299808 502324 299814 502336
rect 299934 502324 299940 502336
rect 299992 502324 299998 502376
rect 347958 502324 347964 502376
rect 348016 502364 348022 502376
rect 348142 502364 348148 502376
rect 348016 502336 348148 502364
rect 348016 502324 348022 502336
rect 348142 502324 348148 502336
rect 348200 502324 348206 502376
rect 364518 502324 364524 502376
rect 364576 502364 364582 502376
rect 364702 502364 364708 502376
rect 364576 502336 364708 502364
rect 364576 502324 364582 502336
rect 364702 502324 364708 502336
rect 364760 502324 364766 502376
rect 412910 502324 412916 502376
rect 412968 502364 412974 502376
rect 413094 502364 413100 502376
rect 412968 502336 413100 502364
rect 412968 502324 412974 502336
rect 413094 502324 413100 502336
rect 413152 502324 413158 502376
rect 429470 502324 429476 502376
rect 429528 502364 429534 502376
rect 429654 502364 429660 502376
rect 429528 502336 429660 502364
rect 429528 502324 429534 502336
rect 429654 502324 429660 502336
rect 429712 502324 429718 502376
rect 477678 502324 477684 502376
rect 477736 502364 477742 502376
rect 477862 502364 477868 502376
rect 477736 502336 477868 502364
rect 477736 502324 477742 502336
rect 477862 502324 477868 502336
rect 477920 502324 477926 502376
rect 494238 502324 494244 502376
rect 494296 502364 494302 502376
rect 494422 502364 494428 502376
rect 494296 502336 494428 502364
rect 494296 502324 494302 502336
rect 494422 502324 494428 502336
rect 494480 502324 494486 502376
rect 542630 502324 542636 502376
rect 542688 502364 542694 502376
rect 542814 502364 542820 502376
rect 542688 502336 542820 502364
rect 542688 502324 542694 502336
rect 542814 502324 542820 502336
rect 542872 502324 542878 502376
rect 559190 502324 559196 502376
rect 559248 502364 559254 502376
rect 559374 502364 559380 502376
rect 559248 502336 559380 502364
rect 559248 502324 559254 502336
rect 559374 502324 559380 502336
rect 559432 502324 559438 502376
rect 569218 498176 569224 498228
rect 569276 498216 569282 498228
rect 580166 498216 580172 498228
rect 569276 498188 580172 498216
rect 569276 498176 569282 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 7926 492600 7932 492652
rect 7984 492640 7990 492652
rect 8110 492640 8116 492652
rect 7984 492612 8116 492640
rect 7984 492600 7990 492612
rect 8110 492600 8116 492612
rect 8168 492600 8174 492652
rect 137646 492600 137652 492652
rect 137704 492640 137710 492652
rect 137830 492640 137836 492652
rect 137704 492612 137836 492640
rect 137704 492600 137710 492612
rect 137830 492600 137836 492612
rect 137888 492600 137894 492652
rect 154206 492600 154212 492652
rect 154264 492640 154270 492652
rect 154390 492640 154396 492652
rect 154264 492612 154396 492640
rect 154264 492600 154270 492612
rect 154390 492600 154396 492612
rect 154448 492600 154454 492652
rect 283098 492640 283104 492652
rect 283059 492612 283104 492640
rect 283098 492600 283104 492612
rect 283156 492600 283162 492652
rect 299658 492640 299664 492652
rect 299619 492612 299664 492640
rect 299658 492600 299664 492612
rect 299716 492600 299722 492652
rect 412818 492640 412824 492652
rect 412779 492612 412824 492640
rect 412818 492600 412824 492612
rect 412876 492600 412882 492652
rect 429378 492640 429384 492652
rect 429339 492612 429384 492640
rect 429378 492600 429384 492612
rect 429436 492600 429442 492652
rect 542538 492640 542544 492652
rect 542499 492612 542544 492640
rect 542538 492600 542544 492612
rect 542596 492600 542602 492652
rect 559098 492640 559104 492652
rect 559059 492612 559104 492640
rect 559098 492600 559104 492612
rect 559156 492600 559162 492652
rect 554038 485800 554044 485852
rect 554096 485840 554102 485852
rect 579890 485840 579896 485852
rect 554096 485812 579896 485840
rect 554096 485800 554102 485812
rect 579890 485800 579896 485812
rect 579948 485800 579954 485852
rect 283098 485772 283104 485784
rect 283059 485744 283104 485772
rect 283098 485732 283104 485744
rect 283156 485732 283162 485784
rect 299658 485772 299664 485784
rect 299619 485744 299664 485772
rect 299658 485732 299664 485744
rect 299716 485732 299722 485784
rect 412818 485772 412824 485784
rect 412779 485744 412824 485772
rect 412818 485732 412824 485744
rect 412876 485732 412882 485784
rect 429378 485772 429384 485784
rect 429339 485744 429384 485772
rect 429378 485732 429384 485744
rect 429436 485732 429442 485784
rect 542538 485772 542544 485784
rect 542499 485744 542544 485772
rect 542538 485732 542544 485744
rect 542596 485732 542602 485784
rect 559098 485772 559104 485784
rect 559059 485744 559104 485772
rect 559098 485732 559104 485744
rect 559156 485732 559162 485784
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 10318 480264 10324 480276
rect 3200 480236 10324 480264
rect 3200 480224 3206 480236
rect 10318 480224 10324 480236
rect 10376 480224 10382 480276
rect 72878 480224 72884 480276
rect 72936 480264 72942 480276
rect 73062 480264 73068 480276
rect 72936 480236 73068 480264
rect 72936 480224 72942 480236
rect 73062 480224 73068 480236
rect 73120 480224 73126 480276
rect 218054 480224 218060 480276
rect 218112 480264 218118 480276
rect 218238 480264 218244 480276
rect 218112 480236 218244 480264
rect 218112 480224 218118 480236
rect 218238 480224 218244 480236
rect 218296 480224 218302 480276
rect 234614 480224 234620 480276
rect 234672 480264 234678 480276
rect 234798 480264 234804 480276
rect 234672 480236 234804 480264
rect 234672 480224 234678 480236
rect 234798 480224 234804 480236
rect 234856 480224 234862 480276
rect 347774 480224 347780 480276
rect 347832 480264 347838 480276
rect 347958 480264 347964 480276
rect 347832 480236 347964 480264
rect 347832 480224 347838 480236
rect 347958 480224 347964 480236
rect 348016 480224 348022 480276
rect 364334 480224 364340 480276
rect 364392 480264 364398 480276
rect 364518 480264 364524 480276
rect 364392 480236 364524 480264
rect 364392 480224 364398 480236
rect 364518 480224 364524 480236
rect 364576 480224 364582 480276
rect 477494 480224 477500 480276
rect 477552 480264 477558 480276
rect 477678 480264 477684 480276
rect 477552 480236 477684 480264
rect 477552 480224 477558 480236
rect 477678 480224 477684 480236
rect 477736 480224 477742 480276
rect 494054 480224 494060 480276
rect 494112 480264 494118 480276
rect 494238 480264 494244 480276
rect 494112 480236 494244 480264
rect 494112 480224 494118 480236
rect 494238 480224 494244 480236
rect 494296 480224 494302 480276
rect 283006 476076 283012 476128
rect 283064 476116 283070 476128
rect 283190 476116 283196 476128
rect 283064 476088 283196 476116
rect 283064 476076 283070 476088
rect 283190 476076 283196 476088
rect 283248 476076 283254 476128
rect 299566 476076 299572 476128
rect 299624 476116 299630 476128
rect 299750 476116 299756 476128
rect 299624 476088 299756 476116
rect 299624 476076 299630 476088
rect 299750 476076 299756 476088
rect 299808 476076 299814 476128
rect 412726 476076 412732 476128
rect 412784 476116 412790 476128
rect 412910 476116 412916 476128
rect 412784 476088 412916 476116
rect 412784 476076 412790 476088
rect 412910 476076 412916 476088
rect 412968 476076 412974 476128
rect 429286 476076 429292 476128
rect 429344 476116 429350 476128
rect 429470 476116 429476 476128
rect 429344 476088 429476 476116
rect 429344 476076 429350 476088
rect 429470 476076 429476 476088
rect 429528 476076 429534 476128
rect 542446 476076 542452 476128
rect 542504 476116 542510 476128
rect 542630 476116 542636 476128
rect 542504 476088 542636 476116
rect 542504 476076 542510 476088
rect 542630 476076 542636 476088
rect 542688 476076 542694 476128
rect 559006 476076 559012 476128
rect 559064 476116 559070 476128
rect 559190 476116 559196 476128
rect 559064 476088 559196 476116
rect 559064 476076 559070 476088
rect 559190 476076 559196 476088
rect 559248 476076 559254 476128
rect 8018 473288 8024 473340
rect 8076 473328 8082 473340
rect 8110 473328 8116 473340
rect 8076 473300 8116 473328
rect 8076 473288 8082 473300
rect 8110 473288 8116 473300
rect 8168 473288 8174 473340
rect 137462 473288 137468 473340
rect 137520 473328 137526 473340
rect 137738 473328 137744 473340
rect 137520 473300 137744 473328
rect 137520 473288 137526 473300
rect 137738 473288 137744 473300
rect 137796 473288 137802 473340
rect 283098 473328 283104 473340
rect 283059 473300 283104 473328
rect 283098 473288 283104 473300
rect 283156 473288 283162 473340
rect 299658 473328 299664 473340
rect 299619 473300 299664 473328
rect 299658 473288 299664 473300
rect 299716 473288 299722 473340
rect 412818 473328 412824 473340
rect 412779 473300 412824 473328
rect 412818 473288 412824 473300
rect 412876 473288 412882 473340
rect 429378 473328 429384 473340
rect 429339 473300 429384 473328
rect 429378 473288 429384 473300
rect 429436 473288 429442 473340
rect 542538 473328 542544 473340
rect 542499 473300 542544 473328
rect 542538 473288 542544 473300
rect 542596 473288 542602 473340
rect 559098 473328 559104 473340
rect 559059 473300 559104 473328
rect 559098 473288 559104 473300
rect 559156 473288 559162 473340
rect 154298 466420 154304 466472
rect 154356 466460 154362 466472
rect 154482 466460 154488 466472
rect 154356 466432 154488 466460
rect 154356 466420 154362 466432
rect 154482 466420 154488 466432
rect 154540 466420 154546 466472
rect 283098 466392 283104 466404
rect 283059 466364 283104 466392
rect 283098 466352 283104 466364
rect 283156 466352 283162 466404
rect 299658 466392 299664 466404
rect 299619 466364 299664 466392
rect 299658 466352 299664 466364
rect 299716 466352 299722 466404
rect 412818 466392 412824 466404
rect 412779 466364 412824 466392
rect 412818 466352 412824 466364
rect 412876 466352 412882 466404
rect 429378 466392 429384 466404
rect 429339 466364 429384 466392
rect 429378 466352 429384 466364
rect 429436 466352 429442 466404
rect 542538 466392 542544 466404
rect 542499 466364 542544 466392
rect 542538 466352 542544 466364
rect 542596 466352 542602 466404
rect 559098 466392 559104 466404
rect 559059 466364 559104 466392
rect 559098 466352 559104 466364
rect 559156 466352 559162 466404
rect 571978 462340 571984 462392
rect 572036 462380 572042 462392
rect 580166 462380 580172 462392
rect 572036 462352 580172 462380
rect 572036 462340 572042 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 72878 460912 72884 460964
rect 72936 460952 72942 460964
rect 73062 460952 73068 460964
rect 72936 460924 73068 460952
rect 72936 460912 72942 460924
rect 73062 460912 73068 460924
rect 73120 460912 73126 460964
rect 218054 460912 218060 460964
rect 218112 460952 218118 460964
rect 218238 460952 218244 460964
rect 218112 460924 218244 460952
rect 218112 460912 218118 460924
rect 218238 460912 218244 460924
rect 218296 460912 218302 460964
rect 234614 460912 234620 460964
rect 234672 460952 234678 460964
rect 234798 460952 234804 460964
rect 234672 460924 234804 460952
rect 234672 460912 234678 460924
rect 234798 460912 234804 460924
rect 234856 460912 234862 460964
rect 347774 460912 347780 460964
rect 347832 460952 347838 460964
rect 347958 460952 347964 460964
rect 347832 460924 347964 460952
rect 347832 460912 347838 460924
rect 347958 460912 347964 460924
rect 348016 460912 348022 460964
rect 364334 460912 364340 460964
rect 364392 460952 364398 460964
rect 364518 460952 364524 460964
rect 364392 460924 364524 460952
rect 364392 460912 364398 460924
rect 364518 460912 364524 460924
rect 364576 460912 364582 460964
rect 477494 460912 477500 460964
rect 477552 460952 477558 460964
rect 477678 460952 477684 460964
rect 477552 460924 477684 460952
rect 477552 460912 477558 460924
rect 477678 460912 477684 460924
rect 477736 460912 477742 460964
rect 494054 460912 494060 460964
rect 494112 460952 494118 460964
rect 494238 460952 494244 460964
rect 494112 460924 494244 460952
rect 494112 460912 494118 460924
rect 494238 460912 494244 460924
rect 494296 460912 494302 460964
rect 299566 453948 299572 453960
rect 299527 453920 299572 453948
rect 299566 453908 299572 453920
rect 299624 453908 299630 453960
rect 3050 451256 3056 451308
rect 3108 451296 3114 451308
rect 6178 451296 6184 451308
rect 3108 451268 6184 451296
rect 3108 451256 3114 451268
rect 6178 451256 6184 451268
rect 6236 451256 6242 451308
rect 8018 447108 8024 447160
rect 8076 447108 8082 447160
rect 137738 447108 137744 447160
rect 137796 447108 137802 447160
rect 154298 447108 154304 447160
rect 154356 447108 154362 447160
rect 282914 447108 282920 447160
rect 282972 447108 282978 447160
rect 412634 447108 412640 447160
rect 412692 447108 412698 447160
rect 429194 447108 429200 447160
rect 429252 447108 429258 447160
rect 542354 447108 542360 447160
rect 542412 447108 542418 447160
rect 558914 447108 558920 447160
rect 558972 447108 558978 447160
rect 8036 447080 8064 447108
rect 8110 447080 8116 447092
rect 8036 447052 8116 447080
rect 8110 447040 8116 447052
rect 8168 447040 8174 447092
rect 137756 447080 137784 447108
rect 137830 447080 137836 447092
rect 137756 447052 137836 447080
rect 137830 447040 137836 447052
rect 137888 447040 137894 447092
rect 154316 447080 154344 447108
rect 154390 447080 154396 447092
rect 154316 447052 154396 447080
rect 154390 447040 154396 447052
rect 154448 447040 154454 447092
rect 282932 447080 282960 447108
rect 283006 447080 283012 447092
rect 282932 447052 283012 447080
rect 283006 447040 283012 447052
rect 283064 447040 283070 447092
rect 299566 447080 299572 447092
rect 299527 447052 299572 447080
rect 299566 447040 299572 447052
rect 299624 447040 299630 447092
rect 412652 447080 412680 447108
rect 412726 447080 412732 447092
rect 412652 447052 412732 447080
rect 412726 447040 412732 447052
rect 412784 447040 412790 447092
rect 429212 447080 429240 447108
rect 429286 447080 429292 447092
rect 429212 447052 429292 447080
rect 429286 447040 429292 447052
rect 429344 447040 429350 447092
rect 542372 447080 542400 447108
rect 542446 447080 542452 447092
rect 542372 447052 542452 447080
rect 542446 447040 542452 447052
rect 542504 447040 542510 447092
rect 558932 447080 558960 447108
rect 559006 447080 559012 447092
rect 558932 447052 559012 447080
rect 559006 447040 559012 447052
rect 559064 447040 559070 447092
rect 8110 444360 8116 444372
rect 8071 444332 8116 444360
rect 8110 444320 8116 444332
rect 8168 444320 8174 444372
rect 137830 444360 137836 444372
rect 137791 444332 137836 444360
rect 137830 444320 137836 444332
rect 137888 444320 137894 444372
rect 154390 444360 154396 444372
rect 154351 444332 154396 444360
rect 154390 444320 154396 444332
rect 154448 444320 154454 444372
rect 218054 441600 218060 441652
rect 218112 441640 218118 441652
rect 218238 441640 218244 441652
rect 218112 441612 218244 441640
rect 218112 441600 218118 441612
rect 218238 441600 218244 441612
rect 218296 441600 218302 441652
rect 234614 441600 234620 441652
rect 234672 441640 234678 441652
rect 234798 441640 234804 441652
rect 234672 441612 234804 441640
rect 234672 441600 234678 441612
rect 234798 441600 234804 441612
rect 234856 441600 234862 441652
rect 347774 441600 347780 441652
rect 347832 441640 347838 441652
rect 347958 441640 347964 441652
rect 347832 441612 347964 441640
rect 347832 441600 347838 441612
rect 347958 441600 347964 441612
rect 348016 441600 348022 441652
rect 364334 441600 364340 441652
rect 364392 441640 364398 441652
rect 364518 441640 364524 441652
rect 364392 441612 364524 441640
rect 364392 441600 364398 441612
rect 364518 441600 364524 441612
rect 364576 441600 364582 441652
rect 477494 441600 477500 441652
rect 477552 441640 477558 441652
rect 477678 441640 477684 441652
rect 477552 441612 477684 441640
rect 477552 441600 477558 441612
rect 477678 441600 477684 441612
rect 477736 441600 477742 441652
rect 494054 441600 494060 441652
rect 494112 441640 494118 441652
rect 494238 441640 494244 441652
rect 494112 441612 494244 441640
rect 494112 441600 494118 441612
rect 494238 441600 494244 441612
rect 494296 441600 494302 441652
rect 560938 438880 560944 438932
rect 560996 438920 561002 438932
rect 580166 438920 580172 438932
rect 560996 438892 580172 438920
rect 560996 438880 561002 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 72786 437452 72792 437504
rect 72844 437492 72850 437504
rect 72970 437492 72976 437504
rect 72844 437464 72976 437492
rect 72844 437452 72850 437464
rect 72970 437452 72976 437464
rect 73028 437452 73034 437504
rect 8110 437424 8116 437436
rect 8071 437396 8116 437424
rect 8110 437384 8116 437396
rect 8168 437384 8174 437436
rect 137830 437424 137836 437436
rect 137791 437396 137836 437424
rect 137830 437384 137836 437396
rect 137888 437384 137894 437436
rect 154390 437424 154396 437436
rect 154351 437396 154396 437424
rect 154390 437384 154396 437396
rect 154448 437384 154454 437436
rect 283098 434704 283104 434716
rect 283059 434676 283104 434704
rect 283098 434664 283104 434676
rect 283156 434664 283162 434716
rect 299658 434704 299664 434716
rect 299619 434676 299664 434704
rect 299658 434664 299664 434676
rect 299716 434664 299722 434716
rect 412818 434704 412824 434716
rect 412779 434676 412824 434704
rect 412818 434664 412824 434676
rect 412876 434664 412882 434716
rect 429378 434704 429384 434716
rect 429339 434676 429384 434704
rect 429378 434664 429384 434676
rect 429436 434664 429442 434716
rect 542538 434704 542544 434716
rect 542499 434676 542544 434704
rect 542538 434664 542544 434676
rect 542596 434664 542602 434716
rect 559098 434704 559104 434716
rect 559059 434676 559104 434704
rect 559098 434664 559104 434676
rect 559156 434664 559162 434716
rect 283098 427768 283104 427780
rect 283059 427740 283104 427768
rect 283098 427728 283104 427740
rect 283156 427728 283162 427780
rect 299658 427768 299664 427780
rect 299619 427740 299664 427768
rect 299658 427728 299664 427740
rect 299716 427728 299722 427780
rect 412818 427768 412824 427780
rect 412779 427740 412824 427768
rect 412818 427728 412824 427740
rect 412876 427728 412882 427780
rect 429378 427768 429384 427780
rect 429339 427740 429384 427768
rect 429378 427728 429384 427740
rect 429436 427728 429442 427780
rect 542538 427768 542544 427780
rect 542499 427740 542544 427768
rect 542538 427728 542544 427740
rect 542596 427728 542602 427780
rect 559098 427768 559104 427780
rect 559059 427740 559104 427768
rect 559098 427728 559104 427740
rect 559156 427728 559162 427780
rect 8018 425076 8024 425128
rect 8076 425116 8082 425128
rect 8202 425116 8208 425128
rect 8076 425088 8208 425116
rect 8076 425076 8082 425088
rect 8202 425076 8208 425088
rect 8260 425076 8266 425128
rect 137738 425076 137744 425128
rect 137796 425116 137802 425128
rect 137922 425116 137928 425128
rect 137796 425088 137928 425116
rect 137796 425076 137802 425088
rect 137922 425076 137928 425088
rect 137980 425076 137986 425128
rect 154298 425076 154304 425128
rect 154356 425116 154362 425128
rect 154482 425116 154488 425128
rect 154356 425088 154488 425116
rect 154356 425076 154362 425088
rect 154482 425076 154488 425088
rect 154540 425076 154546 425128
rect 300026 424872 300032 424924
rect 300084 424912 300090 424924
rect 397454 424912 397460 424924
rect 300084 424884 397460 424912
rect 300084 424872 300090 424884
rect 397454 424872 397460 424884
rect 397512 424872 397518 424924
rect 311802 424804 311808 424856
rect 311860 424844 311866 424856
rect 412910 424844 412916 424856
rect 311860 424816 412916 424844
rect 311860 424804 311866 424816
rect 412910 424804 412916 424816
rect 412968 424804 412974 424856
rect 323578 424736 323584 424788
rect 323636 424776 323642 424788
rect 429470 424776 429476 424788
rect 323636 424748 429476 424776
rect 323636 424736 323642 424748
rect 429470 424736 429476 424748
rect 429528 424736 429534 424788
rect 335446 424668 335452 424720
rect 335504 424708 335510 424720
rect 462314 424708 462320 424720
rect 335504 424680 462320 424708
rect 335504 424668 335510 424680
rect 462314 424668 462320 424680
rect 462372 424668 462378 424720
rect 347222 424600 347228 424652
rect 347280 424640 347286 424652
rect 477678 424640 477684 424652
rect 347280 424612 477684 424640
rect 347280 424600 347286 424612
rect 477678 424600 477684 424612
rect 477736 424600 477742 424652
rect 72786 424532 72792 424584
rect 72844 424572 72850 424584
rect 123202 424572 123208 424584
rect 72844 424544 123208 424572
rect 72844 424532 72850 424544
rect 123202 424532 123208 424544
rect 123260 424532 123266 424584
rect 252922 424532 252928 424584
rect 252980 424572 252986 424584
rect 299750 424572 299756 424584
rect 252980 424544 299756 424572
rect 252980 424532 252986 424544
rect 299750 424532 299756 424544
rect 299808 424532 299814 424584
rect 358998 424532 359004 424584
rect 359056 424572 359062 424584
rect 494238 424572 494244 424584
rect 359056 424544 494244 424572
rect 359056 424532 359062 424544
rect 494238 424532 494244 424544
rect 494296 424532 494302 424584
rect 41322 424464 41328 424516
rect 41380 424504 41386 424516
rect 111426 424504 111432 424516
rect 41380 424476 111432 424504
rect 41380 424464 41386 424476
rect 111426 424464 111432 424476
rect 111484 424464 111490 424516
rect 264698 424464 264704 424516
rect 264756 424504 264762 424516
rect 331214 424504 331220 424516
rect 264756 424476 331220 424504
rect 264756 424464 264762 424476
rect 331214 424464 331220 424476
rect 331272 424464 331278 424516
rect 370774 424464 370780 424516
rect 370832 424504 370838 424516
rect 527174 424504 527180 424516
rect 370832 424476 527180 424504
rect 370832 424464 370838 424476
rect 527174 424464 527180 424476
rect 527232 424464 527238 424516
rect 24762 424396 24768 424448
rect 24820 424436 24826 424448
rect 99650 424436 99656 424448
rect 24820 424408 99656 424436
rect 24820 424396 24826 424408
rect 99650 424396 99656 424408
rect 99708 424396 99714 424448
rect 106182 424396 106188 424448
rect 106240 424436 106246 424448
rect 146754 424436 146760 424448
rect 106240 424408 146760 424436
rect 106240 424396 106246 424408
rect 146754 424396 146760 424408
rect 146812 424396 146818 424448
rect 154298 424396 154304 424448
rect 154356 424436 154362 424448
rect 170398 424436 170404 424448
rect 154356 424408 170404 424436
rect 154356 424396 154362 424408
rect 170398 424396 170404 424408
rect 170456 424396 170462 424448
rect 205726 424396 205732 424448
rect 205784 424436 205790 424448
rect 218238 424436 218244 424448
rect 205784 424408 218244 424436
rect 205784 424396 205790 424408
rect 218238 424396 218244 424408
rect 218296 424396 218302 424448
rect 229278 424396 229284 424448
rect 229336 424436 229342 424448
rect 266354 424436 266360 424448
rect 229336 424408 266360 424436
rect 229336 424396 229342 424408
rect 266354 424396 266360 424408
rect 266412 424396 266418 424448
rect 276474 424396 276480 424448
rect 276532 424436 276538 424448
rect 347958 424436 347964 424448
rect 276532 424408 347964 424436
rect 276532 424396 276538 424408
rect 347958 424396 347964 424408
rect 348016 424396 348022 424448
rect 382550 424396 382556 424448
rect 382608 424436 382614 424448
rect 542630 424436 542636 424448
rect 382608 424408 542636 424436
rect 382608 424396 382614 424408
rect 542630 424396 542636 424408
rect 542688 424396 542694 424448
rect 8018 424328 8024 424380
rect 8076 424368 8082 424380
rect 87874 424368 87880 424380
rect 8076 424340 87880 424368
rect 8076 424328 8082 424340
rect 87874 424328 87880 424340
rect 87932 424328 87938 424380
rect 89622 424328 89628 424380
rect 89680 424368 89686 424380
rect 134978 424368 134984 424380
rect 89680 424340 134984 424368
rect 89680 424328 89686 424340
rect 134978 424328 134984 424340
rect 135036 424328 135042 424380
rect 137738 424328 137744 424380
rect 137796 424368 137802 424380
rect 158530 424368 158536 424380
rect 137796 424340 158536 424368
rect 137796 424328 137802 424340
rect 158530 424328 158536 424340
rect 158588 424328 158594 424380
rect 171042 424328 171048 424380
rect 171100 424368 171106 424380
rect 182174 424368 182180 424380
rect 171100 424340 182180 424368
rect 171100 424328 171106 424340
rect 182174 424328 182180 424340
rect 182232 424328 182238 424380
rect 217502 424328 217508 424380
rect 217560 424368 217566 424380
rect 234798 424368 234804 424380
rect 217560 424340 234804 424368
rect 217560 424328 217566 424340
rect 234798 424328 234804 424340
rect 234856 424328 234862 424380
rect 241054 424328 241060 424380
rect 241112 424368 241118 424380
rect 283190 424368 283196 424380
rect 241112 424340 283196 424368
rect 241112 424328 241118 424340
rect 283190 424328 283196 424340
rect 283248 424328 283254 424380
rect 288250 424328 288256 424380
rect 288308 424368 288314 424380
rect 364518 424368 364524 424380
rect 288308 424340 364524 424368
rect 288308 424328 288314 424340
rect 364518 424328 364524 424340
rect 364576 424328 364582 424380
rect 394326 424328 394332 424380
rect 394384 424368 394390 424380
rect 559190 424368 559196 424380
rect 394384 424340 559196 424368
rect 394384 424328 394390 424340
rect 559190 424328 559196 424340
rect 559248 424328 559254 424380
rect 3326 423648 3332 423700
rect 3384 423688 3390 423700
rect 7558 423688 7564 423700
rect 3384 423660 7564 423688
rect 3384 423648 3390 423660
rect 7558 423648 7564 423660
rect 7616 423648 7622 423700
rect 193950 423648 193956 423700
rect 194008 423688 194014 423700
rect 201494 423688 201500 423700
rect 194008 423660 201500 423688
rect 194008 423648 194014 423660
rect 201494 423648 201500 423660
rect 201552 423648 201558 423700
rect 8938 419432 8944 419484
rect 8996 419472 9002 419484
rect 78674 419472 78680 419484
rect 8996 419444 78680 419472
rect 8996 419432 9002 419444
rect 78674 419432 78680 419444
rect 78732 419432 78738 419484
rect 401594 419432 401600 419484
rect 401652 419472 401658 419484
rect 567838 419472 567844 419484
rect 401652 419444 567844 419472
rect 401652 419432 401658 419444
rect 567838 419432 567844 419444
rect 567896 419432 567902 419484
rect 425698 415420 425704 415472
rect 425756 415460 425762 415472
rect 580166 415460 580172 415472
rect 425756 415432 580172 415460
rect 425756 415420 425762 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 401594 412564 401600 412616
rect 401652 412604 401658 412616
rect 580258 412604 580264 412616
rect 401652 412576 580264 412604
rect 401652 412564 401658 412576
rect 580258 412564 580264 412576
rect 580316 412564 580322 412616
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 78674 411244 78680 411256
rect 3476 411216 78680 411244
rect 3476 411204 3482 411216
rect 78674 411204 78680 411216
rect 78732 411204 78738 411256
rect 401594 405628 401600 405680
rect 401652 405668 401658 405680
rect 558178 405668 558184 405680
rect 401652 405640 558184 405668
rect 401652 405628 401658 405640
rect 558178 405628 558184 405640
rect 558236 405628 558242 405680
rect 14458 404268 14464 404320
rect 14516 404308 14522 404320
rect 78674 404308 78680 404320
rect 14516 404280 78680 404308
rect 14516 404268 14522 404280
rect 78674 404268 78680 404280
rect 78732 404268 78738 404320
rect 401594 398760 401600 398812
rect 401652 398800 401658 398812
rect 566458 398800 566464 398812
rect 401652 398772 566464 398800
rect 401652 398760 401658 398772
rect 566458 398760 566464 398772
rect 566516 398760 566522 398812
rect 29638 395972 29644 396024
rect 29696 396012 29702 396024
rect 78674 396012 78680 396024
rect 29696 395984 78680 396012
rect 29696 395972 29702 395984
rect 78674 395972 78680 395984
rect 78732 395972 78738 396024
rect 3142 394680 3148 394732
rect 3200 394720 3206 394732
rect 21358 394720 21364 394732
rect 3200 394692 21364 394720
rect 3200 394680 3206 394692
rect 21358 394680 21364 394692
rect 21416 394680 21422 394732
rect 407758 391960 407764 392012
rect 407816 392000 407822 392012
rect 580166 392000 580172 392012
rect 407816 391972 580172 392000
rect 407816 391960 407822 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 401594 390464 401600 390516
rect 401652 390504 401658 390516
rect 573358 390504 573364 390516
rect 401652 390476 573364 390504
rect 401652 390464 401658 390476
rect 573358 390464 573364 390476
rect 573416 390464 573422 390516
rect 3510 389104 3516 389156
rect 3568 389144 3574 389156
rect 78674 389144 78680 389156
rect 3568 389116 78680 389144
rect 3568 389104 3574 389116
rect 78674 389104 78680 389116
rect 78732 389104 78738 389156
rect 401594 383596 401600 383648
rect 401652 383636 401658 383648
rect 556798 383636 556804 383648
rect 401652 383608 556804 383636
rect 401652 383596 401658 383608
rect 556798 383596 556804 383608
rect 556856 383596 556862 383648
rect 44818 380808 44824 380860
rect 44876 380848 44882 380860
rect 78674 380848 78680 380860
rect 44876 380820 78680 380848
rect 44876 380808 44882 380820
rect 78674 380808 78680 380820
rect 78732 380808 78738 380860
rect 401594 376660 401600 376712
rect 401652 376700 401658 376712
rect 565078 376700 565084 376712
rect 401652 376672 565084 376700
rect 401652 376660 401658 376672
rect 565078 376660 565084 376672
rect 565136 376660 565142 376712
rect 13078 373940 13084 373992
rect 13136 373980 13142 373992
rect 78674 373980 78680 373992
rect 13136 373952 78680 373980
rect 13136 373940 13142 373952
rect 78674 373940 78680 373952
rect 78732 373940 78738 373992
rect 401594 369792 401600 369844
rect 401652 369832 401658 369844
rect 570598 369832 570604 369844
rect 401652 369804 570604 369832
rect 401652 369792 401658 369804
rect 570598 369792 570604 369804
rect 570656 369792 570662 369844
rect 576118 368500 576124 368552
rect 576176 368540 576182 368552
rect 580166 368540 580172 368552
rect 576176 368512 580172 368540
rect 576176 368500 576182 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3602 365644 3608 365696
rect 3660 365684 3666 365696
rect 78674 365684 78680 365696
rect 3660 365656 78680 365684
rect 3660 365644 3666 365656
rect 78674 365644 78680 365656
rect 78732 365644 78738 365696
rect 401594 362856 401600 362908
rect 401652 362896 401658 362908
rect 555418 362896 555424 362908
rect 401652 362868 555424 362896
rect 401652 362856 401658 362868
rect 555418 362856 555424 362868
rect 555476 362856 555482 362908
rect 17218 358708 17224 358760
rect 17276 358748 17282 358760
rect 78674 358748 78680 358760
rect 17276 358720 78680 358748
rect 17276 358708 17282 358720
rect 78674 358708 78680 358720
rect 78732 358708 78738 358760
rect 404998 357416 405004 357468
rect 405056 357456 405062 357468
rect 579890 357456 579896 357468
rect 405056 357428 579896 357456
rect 405056 357416 405062 357428
rect 579890 357416 579896 357428
rect 579948 357416 579954 357468
rect 401594 355988 401600 356040
rect 401652 356028 401658 356040
rect 563698 356028 563704 356040
rect 401652 356000 563704 356028
rect 401652 355988 401658 356000
rect 563698 355988 563704 356000
rect 563756 355988 563762 356040
rect 39298 350480 39304 350532
rect 39356 350520 39362 350532
rect 78674 350520 78680 350532
rect 39356 350492 78680 350520
rect 39356 350480 39362 350492
rect 78674 350480 78680 350492
rect 78732 350480 78738 350532
rect 401594 347692 401600 347744
rect 401652 347732 401658 347744
rect 552658 347732 552664 347744
rect 401652 347704 552664 347732
rect 401652 347692 401658 347704
rect 552658 347692 552664 347704
rect 552716 347692 552722 347744
rect 403618 345040 403624 345092
rect 403676 345080 403682 345092
rect 580166 345080 580172 345092
rect 403676 345052 580172 345080
rect 403676 345040 403682 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3694 343544 3700 343596
rect 3752 343584 3758 343596
rect 78674 343584 78680 343596
rect 3752 343556 78680 343584
rect 3752 343544 3758 343556
rect 78674 343544 78680 343556
rect 78732 343544 78738 343596
rect 401594 340824 401600 340876
rect 401652 340864 401658 340876
rect 578878 340864 578884 340876
rect 401652 340836 578884 340864
rect 401652 340824 401658 340836
rect 578878 340824 578884 340836
rect 578936 340824 578942 340876
rect 3050 336744 3056 336796
rect 3108 336784 3114 336796
rect 37918 336784 37924 336796
rect 3108 336756 37924 336784
rect 3108 336744 3114 336756
rect 37918 336744 37924 336756
rect 37976 336744 37982 336796
rect 10318 335248 10324 335300
rect 10376 335288 10382 335300
rect 78674 335288 78680 335300
rect 10376 335260 78680 335288
rect 10376 335248 10382 335260
rect 78674 335248 78680 335260
rect 78732 335248 78738 335300
rect 401594 333888 401600 333940
rect 401652 333928 401658 333940
rect 551278 333928 551284 333940
rect 401652 333900 551284 333928
rect 401652 333888 401658 333900
rect 551278 333888 551284 333900
rect 551336 333888 551342 333940
rect 6178 327020 6184 327072
rect 6236 327060 6242 327072
rect 78674 327060 78680 327072
rect 6236 327032 78680 327060
rect 6236 327020 6242 327032
rect 78674 327020 78680 327032
rect 78732 327020 78738 327072
rect 401594 327020 401600 327072
rect 401652 327060 401658 327072
rect 569218 327060 569224 327072
rect 401652 327032 569224 327060
rect 401652 327020 401658 327032
rect 569218 327020 569224 327032
rect 569276 327020 569282 327072
rect 3786 320084 3792 320136
rect 3844 320124 3850 320136
rect 78674 320124 78680 320136
rect 3844 320096 78680 320124
rect 3844 320084 3850 320096
rect 78674 320084 78680 320096
rect 78732 320084 78738 320136
rect 401594 320084 401600 320136
rect 401652 320124 401658 320136
rect 554038 320124 554044 320136
rect 401652 320096 554044 320124
rect 401652 320084 401658 320096
rect 554038 320084 554044 320096
rect 554096 320084 554102 320136
rect 401594 313216 401600 313268
rect 401652 313256 401658 313268
rect 571978 313256 571984 313268
rect 401652 313228 571984 313256
rect 401652 313216 401658 313228
rect 571978 313216 571984 313228
rect 572036 313216 572042 313268
rect 7558 311788 7564 311840
rect 7616 311828 7622 311840
rect 78674 311828 78680 311840
rect 7616 311800 78680 311828
rect 7616 311788 7622 311800
rect 78674 311788 78680 311800
rect 78732 311788 78738 311840
rect 409138 310496 409144 310548
rect 409196 310536 409202 310548
rect 579614 310536 579620 310548
rect 409196 310508 579620 310536
rect 409196 310496 409202 310508
rect 579614 310496 579620 310508
rect 579672 310496 579678 310548
rect 402238 305600 402244 305652
rect 402296 305640 402302 305652
rect 578878 305640 578884 305652
rect 402296 305612 578884 305640
rect 402296 305600 402302 305612
rect 578878 305600 578884 305612
rect 578936 305600 578942 305652
rect 21358 304920 21364 304972
rect 21416 304960 21422 304972
rect 78674 304960 78680 304972
rect 21416 304932 78680 304960
rect 21416 304920 21422 304932
rect 78674 304920 78680 304932
rect 78732 304920 78738 304972
rect 401594 304920 401600 304972
rect 401652 304960 401658 304972
rect 580350 304960 580356 304972
rect 401652 304932 580356 304960
rect 401652 304920 401658 304932
rect 580350 304920 580356 304932
rect 580408 304920 580414 304972
rect 401594 298052 401600 298104
rect 401652 298092 401658 298104
rect 560938 298092 560944 298104
rect 401652 298064 560944 298092
rect 401652 298052 401658 298064
rect 560938 298052 560944 298064
rect 560996 298052 561002 298104
rect 3418 296624 3424 296676
rect 3476 296664 3482 296676
rect 78674 296664 78680 296676
rect 3476 296636 78680 296664
rect 3476 296624 3482 296636
rect 78674 296624 78680 296636
rect 78732 296624 78738 296676
rect 401594 291116 401600 291168
rect 401652 291156 401658 291168
rect 425698 291156 425704 291168
rect 401652 291128 425704 291156
rect 401652 291116 401658 291128
rect 425698 291116 425704 291128
rect 425756 291116 425762 291168
rect 3510 289756 3516 289808
rect 3568 289796 3574 289808
rect 78674 289796 78680 289808
rect 3568 289768 78680 289796
rect 3568 289756 3574 289768
rect 78674 289756 78680 289768
rect 78732 289756 78738 289808
rect 401594 284248 401600 284300
rect 401652 284288 401658 284300
rect 580258 284288 580264 284300
rect 401652 284260 580264 284288
rect 401652 284248 401658 284260
rect 580258 284248 580264 284260
rect 580316 284248 580322 284300
rect 37918 281460 37924 281512
rect 37976 281500 37982 281512
rect 78674 281500 78680 281512
rect 37976 281472 78680 281500
rect 37976 281460 37982 281472
rect 78674 281460 78680 281472
rect 78732 281460 78738 281512
rect 401594 277312 401600 277364
rect 401652 277352 401658 277364
rect 407758 277352 407764 277364
rect 401652 277324 407764 277352
rect 401652 277312 401658 277324
rect 407758 277312 407764 277324
rect 407816 277312 407822 277364
rect 425698 274660 425704 274712
rect 425756 274700 425762 274712
rect 580166 274700 580172 274712
rect 425756 274672 580172 274700
rect 425756 274660 425762 274672
rect 580166 274660 580172 274672
rect 580224 274660 580230 274712
rect 3602 274592 3608 274644
rect 3660 274632 3666 274644
rect 78674 274632 78680 274644
rect 3660 274604 78680 274632
rect 3660 274592 3666 274604
rect 78674 274592 78680 274604
rect 78732 274592 78738 274644
rect 401594 270444 401600 270496
rect 401652 270484 401658 270496
rect 576118 270484 576124 270496
rect 401652 270456 576124 270484
rect 401652 270444 401658 270456
rect 576118 270444 576124 270456
rect 576176 270444 576182 270496
rect 3694 266296 3700 266348
rect 3752 266336 3758 266348
rect 78674 266336 78680 266348
rect 3752 266308 78680 266336
rect 3752 266296 3758 266308
rect 78674 266296 78680 266308
rect 78732 266296 78738 266348
rect 407758 263576 407764 263628
rect 407816 263616 407822 263628
rect 579798 263616 579804 263628
rect 407816 263588 579804 263616
rect 407816 263576 407822 263588
rect 579798 263576 579804 263588
rect 579856 263576 579862 263628
rect 401594 262148 401600 262200
rect 401652 262188 401658 262200
rect 404998 262188 405004 262200
rect 401652 262160 405004 262188
rect 401652 262148 401658 262160
rect 404998 262148 405004 262160
rect 405056 262148 405062 262200
rect 3418 259360 3424 259412
rect 3476 259400 3482 259412
rect 78674 259400 78680 259412
rect 3476 259372 78680 259400
rect 3476 259360 3482 259372
rect 78674 259360 78680 259372
rect 78732 259360 78738 259412
rect 401594 255076 401600 255128
rect 401652 255116 401658 255128
rect 403618 255116 403624 255128
rect 401652 255088 403624 255116
rect 401652 255076 401658 255088
rect 403618 255076 403624 255088
rect 403676 255076 403682 255128
rect 403618 251200 403624 251252
rect 403676 251240 403682 251252
rect 580166 251240 580172 251252
rect 403676 251212 580172 251240
rect 403676 251200 403682 251212
rect 580166 251200 580172 251212
rect 580224 251200 580230 251252
rect 3510 251132 3516 251184
rect 3568 251172 3574 251184
rect 78674 251172 78680 251184
rect 3568 251144 78680 251172
rect 3568 251132 3574 251144
rect 78674 251132 78680 251144
rect 78732 251132 78738 251184
rect 3602 244196 3608 244248
rect 3660 244236 3666 244248
rect 78674 244236 78680 244248
rect 3660 244208 78680 244236
rect 3660 244196 3666 244208
rect 78674 244196 78680 244208
rect 78732 244196 78738 244248
rect 401594 241408 401600 241460
rect 401652 241448 401658 241460
rect 409138 241448 409144 241460
rect 401652 241420 409144 241448
rect 401652 241408 401658 241420
rect 409138 241408 409144 241420
rect 409196 241408 409202 241460
rect 3418 235900 3424 235952
rect 3476 235940 3482 235952
rect 78674 235940 78680 235952
rect 3476 235912 78680 235940
rect 3476 235900 3482 235912
rect 78674 235900 78680 235912
rect 78732 235900 78738 235952
rect 401594 234540 401600 234592
rect 401652 234580 401658 234592
rect 578878 234580 578884 234592
rect 401652 234552 578884 234580
rect 401652 234540 401658 234552
rect 578878 234540 578884 234552
rect 578936 234540 578942 234592
rect 3510 229032 3516 229084
rect 3568 229072 3574 229084
rect 78674 229072 78680 229084
rect 3568 229044 78680 229072
rect 3568 229032 3574 229044
rect 78674 229032 78680 229044
rect 78732 229032 78738 229084
rect 404998 227740 405004 227792
rect 405056 227780 405062 227792
rect 580166 227780 580172 227792
rect 405056 227752 580172 227780
rect 405056 227740 405062 227752
rect 580166 227740 580172 227752
rect 580224 227740 580230 227792
rect 401594 227672 401600 227724
rect 401652 227712 401658 227724
rect 425698 227712 425704 227724
rect 401652 227684 425704 227712
rect 401652 227672 401658 227684
rect 425698 227672 425704 227684
rect 425756 227672 425762 227724
rect 2958 220736 2964 220788
rect 3016 220776 3022 220788
rect 78674 220776 78680 220788
rect 3016 220748 78680 220776
rect 3016 220736 3022 220748
rect 78674 220736 78680 220748
rect 78732 220736 78738 220788
rect 401594 220736 401600 220788
rect 401652 220776 401658 220788
rect 407758 220776 407764 220788
rect 401652 220748 407764 220776
rect 401652 220736 401658 220748
rect 407758 220736 407764 220748
rect 407816 220736 407822 220788
rect 401594 212372 401600 212424
rect 401652 212412 401658 212424
rect 403618 212412 403624 212424
rect 401652 212384 403624 212412
rect 401652 212372 401658 212384
rect 403618 212372 403624 212384
rect 403676 212372 403682 212424
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 79318 208332 79324 208344
rect 3476 208304 79324 208332
rect 3476 208292 3482 208304
rect 79318 208292 79324 208304
rect 79376 208292 79382 208344
rect 401594 205572 401600 205624
rect 401652 205612 401658 205624
rect 404998 205612 405004 205624
rect 401652 205584 405004 205612
rect 401652 205572 401658 205584
rect 404998 205572 405004 205584
rect 405056 205572 405062 205624
rect 401594 198636 401600 198688
rect 401652 198676 401658 198688
rect 580258 198676 580264 198688
rect 401652 198648 580264 198676
rect 401652 198636 401658 198648
rect 580258 198636 580264 198648
rect 580316 198636 580322 198688
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 79318 194528 79324 194540
rect 3200 194500 79324 194528
rect 3200 194488 3206 194500
rect 79318 194488 79324 194500
rect 79376 194488 79382 194540
rect 401594 191768 401600 191820
rect 401652 191808 401658 191820
rect 580350 191808 580356 191820
rect 401652 191780 580356 191808
rect 401652 191768 401658 191780
rect 580350 191768 580356 191780
rect 580408 191768 580414 191820
rect 401594 182112 401600 182164
rect 401652 182152 401658 182164
rect 580166 182152 580172 182164
rect 401652 182124 580172 182152
rect 401652 182112 401658 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 79410 180792 79416 180804
rect 3292 180764 79416 180792
rect 3292 180752 3298 180764
rect 79410 180752 79416 180764
rect 79468 180752 79474 180804
rect 402238 171028 402244 171080
rect 402296 171068 402302 171080
rect 580166 171068 580172 171080
rect 402296 171040 580172 171068
rect 402296 171028 402302 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 21358 165588 21364 165640
rect 21416 165628 21422 165640
rect 78674 165628 78680 165640
rect 21416 165600 78680 165628
rect 21416 165588 21422 165600
rect 78674 165588 78680 165600
rect 78732 165588 78738 165640
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 79318 165560 79324 165572
rect 3568 165532 79324 165560
rect 3568 165520 3574 165532
rect 79318 165520 79324 165532
rect 79376 165520 79382 165572
rect 402238 158652 402244 158704
rect 402296 158692 402302 158704
rect 579798 158692 579804 158704
rect 402296 158664 579804 158692
rect 402296 158652 402302 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 79502 151756 79508 151768
rect 3200 151728 79508 151756
rect 3200 151716 3206 151728
rect 79502 151716 79508 151728
rect 79560 151716 79566 151768
rect 8938 143556 8944 143608
rect 8996 143596 9002 143608
rect 78674 143596 78680 143608
rect 8996 143568 78680 143596
rect 8996 143556 9002 143568
rect 78674 143556 78680 143568
rect 78732 143556 78738 143608
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 79410 136592 79416 136604
rect 3292 136564 79416 136592
rect 3292 136552 3298 136564
rect 79410 136552 79416 136564
rect 79468 136552 79474 136604
rect 402330 135192 402336 135244
rect 402388 135232 402394 135244
rect 580166 135232 580172 135244
rect 402388 135204 580172 135232
rect 402388 135192 402394 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 401594 125604 401600 125656
rect 401652 125644 401658 125656
rect 578878 125644 578884 125656
rect 401652 125616 578884 125644
rect 401652 125604 401658 125616
rect 578878 125604 578884 125616
rect 578936 125604 578942 125656
rect 402238 124108 402244 124160
rect 402296 124148 402302 124160
rect 580166 124148 580172 124160
rect 402296 124120 580172 124148
rect 402296 124108 402302 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 21358 122788 21364 122800
rect 3476 122760 21364 122788
rect 3476 122748 3482 122760
rect 21358 122748 21364 122760
rect 21416 122748 21422 122800
rect 21358 120096 21364 120148
rect 21416 120136 21422 120148
rect 78674 120136 78680 120148
rect 21416 120108 78680 120136
rect 21416 120096 21422 120108
rect 78674 120096 78680 120108
rect 78732 120096 78738 120148
rect 402606 111732 402612 111784
rect 402664 111772 402670 111784
rect 579798 111772 579804 111784
rect 402664 111744 579804 111772
rect 402664 111732 402670 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 79318 108984 79324 108996
rect 3292 108956 79324 108984
rect 3292 108944 3298 108956
rect 79318 108944 79324 108956
rect 79376 108944 79382 108996
rect 401594 104864 401600 104916
rect 401652 104904 401658 104916
rect 555418 104904 555424 104916
rect 401652 104876 555424 104904
rect 401652 104864 401658 104876
rect 555418 104864 555424 104876
rect 555476 104864 555482 104916
rect 370866 102116 370872 102128
rect 370827 102088 370872 102116
rect 370866 102076 370872 102088
rect 370924 102076 370930 102128
rect 89714 100648 89720 100700
rect 89772 100688 89778 100700
rect 90910 100688 90916 100700
rect 89772 100660 90916 100688
rect 89772 100648 89778 100660
rect 90910 100648 90916 100660
rect 90968 100648 90974 100700
rect 97166 100648 97172 100700
rect 97224 100688 97230 100700
rect 97902 100688 97908 100700
rect 97224 100660 97908 100688
rect 97224 100648 97230 100660
rect 97902 100648 97908 100660
rect 97960 100648 97966 100700
rect 97994 100648 98000 100700
rect 98052 100688 98058 100700
rect 99282 100688 99288 100700
rect 98052 100660 99288 100688
rect 98052 100648 98058 100660
rect 99282 100648 99288 100660
rect 99340 100648 99346 100700
rect 99650 100648 99656 100700
rect 99708 100688 99714 100700
rect 100570 100688 100576 100700
rect 99708 100660 100576 100688
rect 99708 100648 99714 100660
rect 100570 100648 100576 100660
rect 100628 100648 100634 100700
rect 102134 100648 102140 100700
rect 102192 100688 102198 100700
rect 103330 100688 103336 100700
rect 102192 100660 103336 100688
rect 102192 100648 102198 100660
rect 103330 100648 103336 100660
rect 103388 100648 103394 100700
rect 105354 100648 105360 100700
rect 105412 100688 105418 100700
rect 106182 100688 106188 100700
rect 105412 100660 106188 100688
rect 105412 100648 105418 100660
rect 106182 100648 106188 100660
rect 106240 100648 106246 100700
rect 107838 100648 107844 100700
rect 107896 100688 107902 100700
rect 108942 100688 108948 100700
rect 107896 100660 108948 100688
rect 107896 100648 107902 100660
rect 108942 100648 108948 100660
rect 109000 100648 109006 100700
rect 153194 100648 153200 100700
rect 153252 100688 153258 100700
rect 154482 100688 154488 100700
rect 153252 100660 154488 100688
rect 153252 100648 153258 100660
rect 154482 100648 154488 100660
rect 154540 100648 154546 100700
rect 154850 100648 154856 100700
rect 154908 100688 154914 100700
rect 155770 100688 155776 100700
rect 154908 100660 155776 100688
rect 154908 100648 154914 100660
rect 155770 100648 155776 100660
rect 155828 100648 155834 100700
rect 201862 100648 201868 100700
rect 201920 100688 201926 100700
rect 202782 100688 202788 100700
rect 201920 100660 202788 100688
rect 201920 100648 201926 100660
rect 202782 100648 202788 100660
rect 202840 100648 202846 100700
rect 204346 100648 204352 100700
rect 204404 100688 204410 100700
rect 205450 100688 205456 100700
rect 204404 100660 205456 100688
rect 204404 100648 204410 100660
rect 205450 100648 205456 100660
rect 205508 100648 205514 100700
rect 234890 100648 234896 100700
rect 234948 100688 234954 100700
rect 236638 100688 236644 100700
rect 234948 100660 236644 100688
rect 234948 100648 234954 100660
rect 236638 100648 236644 100660
rect 236696 100648 236702 100700
rect 237374 100648 237380 100700
rect 237432 100688 237438 100700
rect 238662 100688 238668 100700
rect 237432 100660 238668 100688
rect 237432 100648 237438 100660
rect 238662 100648 238668 100660
rect 238720 100648 238726 100700
rect 243078 100648 243084 100700
rect 243136 100688 243142 100700
rect 244090 100688 244096 100700
rect 243136 100660 244096 100688
rect 243136 100648 243142 100660
rect 244090 100648 244096 100660
rect 244148 100648 244154 100700
rect 263778 100648 263784 100700
rect 263836 100688 263842 100700
rect 264790 100688 264796 100700
rect 263836 100660 264796 100688
rect 263836 100648 263842 100660
rect 264790 100648 264796 100660
rect 264848 100648 264854 100700
rect 267826 100648 267832 100700
rect 267884 100688 267890 100700
rect 269022 100688 269028 100700
rect 267884 100660 269028 100688
rect 267884 100648 267890 100660
rect 269022 100648 269028 100660
rect 269080 100648 269086 100700
rect 271966 100648 271972 100700
rect 272024 100688 272030 100700
rect 273162 100688 273168 100700
rect 272024 100660 273168 100688
rect 272024 100648 272030 100660
rect 273162 100648 273168 100660
rect 273220 100648 273226 100700
rect 276106 100648 276112 100700
rect 276164 100688 276170 100700
rect 277302 100688 277308 100700
rect 276164 100660 277308 100688
rect 276164 100648 276170 100660
rect 277302 100648 277308 100660
rect 277360 100648 277366 100700
rect 345382 100648 345388 100700
rect 345440 100688 345446 100700
rect 346302 100688 346308 100700
rect 345440 100660 346308 100688
rect 345440 100648 345446 100660
rect 346302 100648 346308 100660
rect 346360 100648 346366 100700
rect 347866 100648 347872 100700
rect 347924 100688 347930 100700
rect 348970 100688 348976 100700
rect 347924 100660 348976 100688
rect 347924 100648 347930 100660
rect 348970 100648 348976 100660
rect 349028 100648 349034 100700
rect 349522 100648 349528 100700
rect 349580 100688 349586 100700
rect 350350 100688 350356 100700
rect 349580 100660 350356 100688
rect 349580 100648 349586 100660
rect 350350 100648 350356 100660
rect 350408 100648 350414 100700
rect 370130 100648 370136 100700
rect 370188 100688 370194 100700
rect 371142 100688 371148 100700
rect 370188 100660 371148 100688
rect 370188 100648 370194 100660
rect 371142 100648 371148 100660
rect 371200 100648 371206 100700
rect 374270 100648 374276 100700
rect 374328 100688 374334 100700
rect 375190 100688 375196 100700
rect 374328 100660 375196 100688
rect 374328 100648 374334 100660
rect 375190 100648 375196 100660
rect 375248 100648 375254 100700
rect 375926 100648 375932 100700
rect 375984 100688 375990 100700
rect 376662 100688 376668 100700
rect 375984 100660 376668 100688
rect 375984 100648 375990 100660
rect 376662 100648 376668 100660
rect 376720 100648 376726 100700
rect 93854 100580 93860 100632
rect 93912 100620 93918 100632
rect 97258 100620 97264 100632
rect 93912 100592 97264 100620
rect 93912 100580 93918 100592
rect 97258 100580 97264 100592
rect 97316 100580 97322 100632
rect 265342 100376 265348 100428
rect 265400 100416 265406 100428
rect 266170 100416 266176 100428
rect 265400 100388 266176 100416
rect 265400 100376 265406 100388
rect 266170 100376 266176 100388
rect 266228 100376 266234 100428
rect 262122 100172 262128 100224
rect 262180 100212 262186 100224
rect 291838 100212 291844 100224
rect 262180 100184 291844 100212
rect 262180 100172 262186 100184
rect 291838 100172 291844 100184
rect 291896 100172 291902 100224
rect 293402 100172 293408 100224
rect 293460 100212 293466 100224
rect 309778 100212 309784 100224
rect 293460 100184 309784 100212
rect 293460 100172 293466 100184
rect 309778 100172 309784 100184
rect 309836 100172 309842 100224
rect 379146 100172 379152 100224
rect 379204 100212 379210 100224
rect 403618 100212 403624 100224
rect 379204 100184 403624 100212
rect 379204 100172 379210 100184
rect 403618 100172 403624 100184
rect 403676 100172 403682 100224
rect 152366 100104 152372 100156
rect 152424 100144 152430 100156
rect 153102 100144 153108 100156
rect 152424 100116 153108 100144
rect 152424 100104 152430 100116
rect 153102 100104 153108 100116
rect 153160 100104 153166 100156
rect 165614 100104 165620 100156
rect 165672 100144 165678 100156
rect 174538 100144 174544 100156
rect 165672 100116 174544 100144
rect 165672 100104 165678 100116
rect 174538 100104 174544 100116
rect 174596 100104 174602 100156
rect 180426 100104 180432 100156
rect 180484 100144 180490 100156
rect 203518 100144 203524 100156
rect 180484 100116 203524 100144
rect 180484 100104 180490 100116
rect 203518 100104 203524 100116
rect 203576 100104 203582 100156
rect 217594 100104 217600 100156
rect 217652 100144 217658 100156
rect 224218 100144 224224 100156
rect 217652 100116 224224 100144
rect 217652 100104 217658 100116
rect 224218 100104 224224 100116
rect 224276 100104 224282 100156
rect 240686 100104 240692 100156
rect 240744 100144 240750 100156
rect 241422 100144 241428 100156
rect 240744 100116 241428 100144
rect 240744 100104 240750 100116
rect 241422 100104 241428 100116
rect 241480 100104 241486 100156
rect 246298 100144 246304 100156
rect 244200 100116 246304 100144
rect 108666 100036 108672 100088
rect 108724 100076 108730 100088
rect 135898 100076 135904 100088
rect 108724 100048 135904 100076
rect 108724 100036 108730 100048
rect 135898 100036 135904 100048
rect 135956 100036 135962 100088
rect 172238 100036 172244 100088
rect 172296 100076 172302 100088
rect 198001 100079 198059 100085
rect 198001 100076 198013 100079
rect 172296 100048 198013 100076
rect 172296 100036 172302 100048
rect 198001 100045 198013 100048
rect 198047 100045 198059 100079
rect 198001 100039 198059 100045
rect 221642 100036 221648 100088
rect 221700 100076 221706 100088
rect 231118 100076 231124 100088
rect 221700 100048 231124 100076
rect 221700 100036 221706 100048
rect 231118 100036 231124 100048
rect 231176 100036 231182 100088
rect 238202 100036 238208 100088
rect 238260 100076 238266 100088
rect 244200 100076 244228 100116
rect 246298 100104 246304 100116
rect 246356 100104 246362 100156
rect 255498 100104 255504 100156
rect 255556 100144 255562 100156
rect 261478 100144 261484 100156
rect 255556 100116 261484 100144
rect 255556 100104 255562 100116
rect 261478 100104 261484 100116
rect 261536 100104 261542 100156
rect 280246 100104 280252 100156
rect 280304 100144 280310 100156
rect 281350 100144 281356 100156
rect 280304 100116 281356 100144
rect 280304 100104 280310 100116
rect 281350 100104 281356 100116
rect 281408 100104 281414 100156
rect 289262 100104 289268 100156
rect 289320 100144 289326 100156
rect 322198 100144 322204 100156
rect 289320 100116 322204 100144
rect 289320 100104 289326 100116
rect 322198 100104 322204 100116
rect 322256 100104 322262 100156
rect 335446 100104 335452 100156
rect 335504 100144 335510 100156
rect 355318 100144 355324 100156
rect 335504 100116 355324 100144
rect 335504 100104 335510 100116
rect 355318 100104 355324 100116
rect 355376 100104 355382 100156
rect 372614 100104 372620 100156
rect 372672 100144 372678 100156
rect 373810 100144 373816 100156
rect 372672 100116 373816 100144
rect 372672 100104 372678 100116
rect 373810 100104 373816 100116
rect 373868 100104 373874 100156
rect 392394 100104 392400 100156
rect 392452 100144 392458 100156
rect 446398 100144 446404 100156
rect 392452 100116 446404 100144
rect 392452 100104 392458 100116
rect 446398 100104 446404 100116
rect 446456 100104 446462 100156
rect 238260 100048 244228 100076
rect 238260 100036 238266 100048
rect 261294 100036 261300 100088
rect 261352 100076 261358 100088
rect 294598 100076 294604 100088
rect 261352 100048 294604 100076
rect 261352 100036 261358 100048
rect 294598 100036 294604 100048
rect 294656 100036 294662 100088
rect 331398 100036 331404 100088
rect 331456 100076 331462 100088
rect 420178 100076 420184 100088
rect 331456 100048 420184 100076
rect 331456 100036 331462 100048
rect 420178 100036 420184 100048
rect 420236 100036 420242 100088
rect 85574 99968 85580 100020
rect 85632 100008 85638 100020
rect 106918 100008 106924 100020
rect 85632 99980 106924 100008
rect 85632 99968 85638 99980
rect 106918 99968 106924 99980
rect 106976 99968 106982 100020
rect 133414 99968 133420 100020
rect 133472 100008 133478 100020
rect 178678 100008 178684 100020
rect 133472 99980 178684 100008
rect 133472 99968 133478 99980
rect 178678 99968 178684 99980
rect 178736 99968 178742 100020
rect 197722 99968 197728 100020
rect 197780 100008 197786 100020
rect 266998 100008 267004 100020
rect 197780 99980 267004 100008
rect 197780 99968 197786 99980
rect 266998 99968 267004 99980
rect 267056 99968 267062 100020
rect 271138 99968 271144 100020
rect 271196 100008 271202 100020
rect 272518 100008 272524 100020
rect 271196 99980 272524 100008
rect 271196 99968 271202 99980
rect 272518 99968 272524 99980
rect 272576 99968 272582 100020
rect 273622 99968 273628 100020
rect 273680 100008 273686 100020
rect 283558 100008 283564 100020
rect 273680 99980 283564 100008
rect 273680 99968 273686 99980
rect 283558 99968 283564 99980
rect 283616 99968 283622 100020
rect 292574 99968 292580 100020
rect 292632 100008 292638 100020
rect 300118 100008 300124 100020
rect 292632 99980 300124 100008
rect 292632 99968 292638 99980
rect 300118 99968 300124 99980
rect 300176 99968 300182 100020
rect 309870 99968 309876 100020
rect 309928 100008 309934 100020
rect 344278 100008 344284 100020
rect 309928 99980 344284 100008
rect 309928 99968 309934 99980
rect 344278 99968 344284 99980
rect 344336 99968 344342 100020
rect 384114 99968 384120 100020
rect 384172 100008 384178 100020
rect 493318 100008 493324 100020
rect 384172 99980 493324 100008
rect 384172 99968 384178 99980
rect 493318 99968 493324 99980
rect 493376 99968 493382 100020
rect 269482 99900 269488 99952
rect 269540 99940 269546 99952
rect 270310 99940 270316 99952
rect 269540 99912 270316 99940
rect 269540 99900 269546 99912
rect 270310 99900 270316 99912
rect 270368 99900 270374 99952
rect 376754 99832 376760 99884
rect 376812 99872 376818 99884
rect 377950 99872 377956 99884
rect 376812 99844 377956 99872
rect 376812 99832 376818 99844
rect 377950 99832 377956 99844
rect 378008 99832 378014 99884
rect 95510 99696 95516 99748
rect 95568 99736 95574 99748
rect 96522 99736 96528 99748
rect 95568 99708 96528 99736
rect 95568 99696 95574 99708
rect 96522 99696 96528 99708
rect 96580 99696 96586 99748
rect 149146 99696 149152 99748
rect 149204 99736 149210 99748
rect 150342 99736 150348 99748
rect 149204 99708 150348 99736
rect 149204 99696 149210 99708
rect 150342 99696 150348 99708
rect 150400 99696 150406 99748
rect 150710 99696 150716 99748
rect 150768 99736 150774 99748
rect 151722 99736 151728 99748
rect 150768 99708 151728 99736
rect 150768 99696 150774 99708
rect 151722 99696 151728 99708
rect 151780 99696 151786 99748
rect 200206 99696 200212 99748
rect 200264 99736 200270 99748
rect 201402 99736 201408 99748
rect 200264 99708 201408 99736
rect 200264 99696 200270 99708
rect 201402 99696 201408 99708
rect 201460 99696 201466 99748
rect 239030 99696 239036 99748
rect 239088 99736 239094 99748
rect 240042 99736 240048 99748
rect 239088 99708 240048 99736
rect 239088 99696 239094 99708
rect 240042 99696 240048 99708
rect 240100 99696 240106 99748
rect 281902 99696 281908 99748
rect 281960 99736 281966 99748
rect 282822 99736 282828 99748
rect 281960 99708 282828 99736
rect 281960 99696 281966 99708
rect 282822 99696 282828 99708
rect 282880 99696 282886 99748
rect 103790 99560 103796 99612
rect 103848 99600 103854 99612
rect 104802 99600 104808 99612
rect 103848 99572 104808 99600
rect 103848 99560 103854 99572
rect 104802 99560 104808 99572
rect 104860 99560 104866 99612
rect 306650 99492 306656 99544
rect 306708 99532 306714 99544
rect 313918 99532 313924 99544
rect 306708 99504 313924 99532
rect 306708 99492 306714 99504
rect 313918 99492 313924 99504
rect 313976 99492 313982 99544
rect 87230 99424 87236 99476
rect 87288 99464 87294 99476
rect 88978 99464 88984 99476
rect 87288 99436 88984 99464
rect 87288 99424 87294 99436
rect 88978 99424 88984 99436
rect 89036 99424 89042 99476
rect 130930 99424 130936 99476
rect 130988 99464 130994 99476
rect 131758 99464 131764 99476
rect 130988 99436 131764 99464
rect 130988 99424 130994 99436
rect 131758 99424 131764 99436
rect 131816 99424 131822 99476
rect 164786 99424 164792 99476
rect 164844 99464 164850 99476
rect 169018 99464 169024 99476
rect 164844 99436 169024 99464
rect 164844 99424 164850 99436
rect 169018 99424 169024 99436
rect 169076 99424 169082 99476
rect 183738 99424 183744 99476
rect 183796 99464 183802 99476
rect 186958 99464 186964 99476
rect 183796 99436 186964 99464
rect 183796 99424 183802 99436
rect 186958 99424 186964 99436
rect 187016 99424 187022 99476
rect 202690 99424 202696 99476
rect 202748 99464 202754 99476
rect 207658 99464 207664 99476
rect 202748 99436 207664 99464
rect 202748 99424 202754 99436
rect 207658 99424 207664 99436
rect 207716 99424 207722 99476
rect 241514 99424 241520 99476
rect 241572 99464 241578 99476
rect 250438 99464 250444 99476
rect 241572 99436 250444 99464
rect 241572 99424 241578 99436
rect 250438 99424 250444 99436
rect 250496 99424 250502 99476
rect 302510 99424 302516 99476
rect 302568 99464 302574 99476
rect 304258 99464 304264 99476
rect 302568 99436 304264 99464
rect 302568 99424 302574 99436
rect 304258 99424 304264 99436
rect 304316 99424 304322 99476
rect 311526 99424 311532 99476
rect 311584 99464 311590 99476
rect 318058 99464 318064 99476
rect 311584 99436 318064 99464
rect 311584 99424 311590 99436
rect 318058 99424 318064 99436
rect 318116 99424 318122 99476
rect 361022 99424 361028 99476
rect 361080 99464 361086 99476
rect 363598 99464 363604 99476
rect 361080 99436 363604 99464
rect 361080 99424 361086 99436
rect 363598 99424 363604 99436
rect 363656 99424 363662 99476
rect 364334 99424 364340 99476
rect 364392 99464 364398 99476
rect 367738 99464 367744 99476
rect 364392 99436 367744 99464
rect 364392 99424 364398 99436
rect 367738 99424 367744 99436
rect 367796 99424 367802 99476
rect 378318 99424 378324 99476
rect 378376 99464 378382 99476
rect 381538 99464 381544 99476
rect 378376 99436 381544 99464
rect 378376 99424 378382 99436
rect 381538 99424 381544 99436
rect 381596 99424 381602 99476
rect 383286 99424 383292 99476
rect 383344 99464 383350 99476
rect 385678 99464 385684 99476
rect 383344 99436 385684 99464
rect 383344 99424 383350 99436
rect 385678 99424 385684 99436
rect 385736 99424 385742 99476
rect 88886 99356 88892 99408
rect 88944 99396 88950 99408
rect 89622 99396 89628 99408
rect 88944 99368 89628 99396
rect 88944 99356 88950 99368
rect 89622 99356 89628 99368
rect 89680 99356 89686 99408
rect 109494 99356 109500 99408
rect 109552 99396 109558 99408
rect 111058 99396 111064 99408
rect 109552 99368 111064 99396
rect 109552 99356 109558 99368
rect 111058 99356 111064 99368
rect 111116 99356 111122 99408
rect 111978 99356 111984 99408
rect 112036 99396 112042 99408
rect 115198 99396 115204 99408
rect 112036 99368 115204 99396
rect 112036 99356 112042 99368
rect 115198 99356 115204 99368
rect 115256 99356 115262 99408
rect 116118 99356 116124 99408
rect 116176 99396 116182 99408
rect 117222 99396 117228 99408
rect 116176 99368 117228 99396
rect 116176 99356 116182 99368
rect 117222 99356 117228 99368
rect 117280 99356 117286 99408
rect 117774 99356 117780 99408
rect 117832 99396 117838 99408
rect 118510 99396 118516 99408
rect 117832 99368 118516 99396
rect 117832 99356 117838 99368
rect 118510 99356 118516 99368
rect 118568 99356 118574 99408
rect 120258 99356 120264 99408
rect 120316 99396 120322 99408
rect 121270 99396 121276 99408
rect 120316 99368 121276 99396
rect 120316 99356 120322 99368
rect 121270 99356 121276 99368
rect 121328 99356 121334 99408
rect 121914 99356 121920 99408
rect 121972 99396 121978 99408
rect 122742 99396 122748 99408
rect 121972 99368 122748 99396
rect 121972 99356 121978 99368
rect 122742 99356 122748 99368
rect 122800 99356 122806 99408
rect 124398 99356 124404 99408
rect 124456 99396 124462 99408
rect 125502 99396 125508 99408
rect 124456 99368 125508 99396
rect 124456 99356 124462 99368
rect 125502 99356 125508 99368
rect 125560 99356 125566 99408
rect 126054 99356 126060 99408
rect 126112 99396 126118 99408
rect 126882 99396 126888 99408
rect 126112 99368 126888 99396
rect 126112 99356 126118 99368
rect 126882 99356 126888 99368
rect 126940 99356 126946 99408
rect 128446 99356 128452 99408
rect 128504 99396 128510 99408
rect 129642 99396 129648 99408
rect 128504 99368 129648 99396
rect 128504 99356 128510 99368
rect 129642 99356 129648 99368
rect 129700 99356 129706 99408
rect 130102 99356 130108 99408
rect 130160 99396 130166 99408
rect 131022 99396 131028 99408
rect 130160 99368 131028 99396
rect 130160 99356 130166 99368
rect 131022 99356 131028 99368
rect 131080 99356 131086 99408
rect 132586 99356 132592 99408
rect 132644 99396 132650 99408
rect 133782 99396 133788 99408
rect 132644 99368 133788 99396
rect 132644 99356 132650 99368
rect 133782 99356 133788 99368
rect 133840 99356 133846 99408
rect 134242 99356 134248 99408
rect 134300 99396 134306 99408
rect 135162 99396 135168 99408
rect 134300 99368 135168 99396
rect 134300 99356 134306 99368
rect 135162 99356 135168 99368
rect 135220 99356 135226 99408
rect 136726 99356 136732 99408
rect 136784 99396 136790 99408
rect 137922 99396 137928 99408
rect 136784 99368 137928 99396
rect 136784 99356 136790 99368
rect 137922 99356 137928 99368
rect 137980 99356 137986 99408
rect 138382 99356 138388 99408
rect 138440 99396 138446 99408
rect 139302 99396 139308 99408
rect 138440 99368 139308 99396
rect 138440 99356 138446 99368
rect 139302 99356 139308 99368
rect 139360 99356 139366 99408
rect 140866 99356 140872 99408
rect 140924 99396 140930 99408
rect 142062 99396 142068 99408
rect 140924 99368 142068 99396
rect 140924 99356 140930 99368
rect 142062 99356 142068 99368
rect 142120 99356 142126 99408
rect 142522 99356 142528 99408
rect 142580 99396 142586 99408
rect 143350 99396 143356 99408
rect 142580 99368 143356 99396
rect 142580 99356 142586 99368
rect 143350 99356 143356 99368
rect 143408 99356 143414 99408
rect 145006 99356 145012 99408
rect 145064 99396 145070 99408
rect 146110 99396 146116 99408
rect 145064 99368 146116 99396
rect 145064 99356 145070 99368
rect 146110 99356 146116 99368
rect 146168 99356 146174 99408
rect 146662 99356 146668 99408
rect 146720 99396 146726 99408
rect 147582 99396 147588 99408
rect 146720 99368 147588 99396
rect 146720 99356 146726 99368
rect 147582 99356 147588 99368
rect 147640 99356 147646 99408
rect 157334 99356 157340 99408
rect 157392 99396 157398 99408
rect 158530 99396 158536 99408
rect 157392 99368 158536 99396
rect 157392 99356 157398 99368
rect 158530 99356 158536 99368
rect 158588 99356 158594 99408
rect 158990 99356 158996 99408
rect 159048 99396 159054 99408
rect 159910 99396 159916 99408
rect 159048 99368 159916 99396
rect 159048 99356 159054 99368
rect 159910 99356 159916 99368
rect 159968 99356 159974 99408
rect 160646 99356 160652 99408
rect 160704 99396 160710 99408
rect 161382 99396 161388 99408
rect 160704 99368 161388 99396
rect 160704 99356 160710 99368
rect 161382 99356 161388 99368
rect 161440 99356 161446 99408
rect 161474 99356 161480 99408
rect 161532 99396 161538 99408
rect 162670 99396 162676 99408
rect 161532 99368 162676 99396
rect 161532 99356 161538 99368
rect 162670 99356 162676 99368
rect 162728 99356 162734 99408
rect 163958 99356 163964 99408
rect 164016 99396 164022 99408
rect 164878 99396 164884 99408
rect 164016 99368 164884 99396
rect 164016 99356 164022 99368
rect 164878 99356 164884 99368
rect 164936 99356 164942 99408
rect 167270 99356 167276 99408
rect 167328 99396 167334 99408
rect 168190 99396 168196 99408
rect 167328 99368 168196 99396
rect 167328 99356 167334 99368
rect 168190 99356 168196 99368
rect 168248 99356 168254 99408
rect 168926 99356 168932 99408
rect 168984 99396 168990 99408
rect 169662 99396 169668 99408
rect 168984 99368 169668 99396
rect 168984 99356 168990 99368
rect 169662 99356 169668 99368
rect 169720 99356 169726 99408
rect 169754 99356 169760 99408
rect 169812 99396 169818 99408
rect 170950 99396 170956 99408
rect 169812 99368 170956 99396
rect 169812 99356 169818 99368
rect 170950 99356 170956 99368
rect 171008 99356 171014 99408
rect 171410 99356 171416 99408
rect 171468 99396 171474 99408
rect 172422 99396 172428 99408
rect 171468 99368 172428 99396
rect 171468 99356 171474 99368
rect 172422 99356 172428 99368
rect 172480 99356 172486 99408
rect 173066 99356 173072 99408
rect 173124 99396 173130 99408
rect 173802 99396 173808 99408
rect 173124 99368 173808 99396
rect 173124 99356 173130 99368
rect 173802 99356 173808 99368
rect 173860 99356 173866 99408
rect 175458 99356 175464 99408
rect 175516 99396 175522 99408
rect 176562 99396 176568 99408
rect 175516 99368 176568 99396
rect 175516 99356 175522 99368
rect 176562 99356 176568 99368
rect 176620 99356 176626 99408
rect 179598 99356 179604 99408
rect 179656 99396 179662 99408
rect 180702 99396 180708 99408
rect 179656 99368 180708 99396
rect 179656 99356 179662 99368
rect 180702 99356 180708 99368
rect 180760 99356 180766 99408
rect 181254 99356 181260 99408
rect 181312 99396 181318 99408
rect 182818 99396 182824 99408
rect 181312 99368 182824 99396
rect 181312 99356 181318 99368
rect 182818 99356 182824 99368
rect 182876 99356 182882 99408
rect 185394 99356 185400 99408
rect 185452 99396 185458 99408
rect 186222 99396 186228 99408
rect 185452 99368 186228 99396
rect 185452 99356 185458 99368
rect 186222 99356 186228 99368
rect 186280 99356 186286 99408
rect 187878 99356 187884 99408
rect 187936 99396 187942 99408
rect 188982 99396 188988 99408
rect 187936 99368 188988 99396
rect 187936 99356 187942 99368
rect 188982 99356 188988 99368
rect 189040 99356 189046 99408
rect 189534 99356 189540 99408
rect 189592 99396 189598 99408
rect 191098 99396 191104 99408
rect 189592 99368 191104 99396
rect 189592 99356 189598 99368
rect 191098 99356 191104 99368
rect 191156 99356 191162 99408
rect 192018 99356 192024 99408
rect 192076 99396 192082 99408
rect 193030 99396 193036 99408
rect 192076 99368 193036 99396
rect 192076 99356 192082 99368
rect 193030 99356 193036 99368
rect 193088 99356 193094 99408
rect 206002 99356 206008 99408
rect 206060 99396 206066 99408
rect 206830 99396 206836 99408
rect 206060 99368 206836 99396
rect 206060 99356 206066 99368
rect 206830 99356 206836 99368
rect 206888 99356 206894 99408
rect 208486 99356 208492 99408
rect 208544 99396 208550 99408
rect 209590 99396 209596 99408
rect 208544 99368 209596 99396
rect 208544 99356 208550 99368
rect 209590 99356 209596 99368
rect 209648 99356 209654 99408
rect 210142 99356 210148 99408
rect 210200 99396 210206 99408
rect 210970 99396 210976 99408
rect 210200 99368 210976 99396
rect 210200 99356 210206 99368
rect 210970 99356 210976 99368
rect 211028 99356 211034 99408
rect 212626 99356 212632 99408
rect 212684 99396 212690 99408
rect 213822 99396 213828 99408
rect 212684 99368 213828 99396
rect 212684 99356 212690 99368
rect 213822 99356 213828 99368
rect 213880 99356 213886 99408
rect 214282 99356 214288 99408
rect 214340 99396 214346 99408
rect 215938 99396 215944 99408
rect 214340 99368 215944 99396
rect 214340 99356 214346 99368
rect 215938 99356 215944 99368
rect 215996 99356 216002 99408
rect 216766 99356 216772 99408
rect 216824 99396 216830 99408
rect 217962 99396 217968 99408
rect 216824 99368 217968 99396
rect 216824 99356 216830 99368
rect 217962 99356 217968 99368
rect 218020 99356 218026 99408
rect 218422 99356 218428 99408
rect 218480 99396 218486 99408
rect 219250 99396 219256 99408
rect 218480 99368 219256 99396
rect 218480 99356 218486 99368
rect 219250 99356 219256 99368
rect 219308 99356 219314 99408
rect 220814 99356 220820 99408
rect 220872 99396 220878 99408
rect 222102 99396 222108 99408
rect 220872 99368 222108 99396
rect 220872 99356 220878 99368
rect 222102 99356 222108 99368
rect 222160 99356 222166 99408
rect 222470 99356 222476 99408
rect 222528 99396 222534 99408
rect 223390 99396 223396 99408
rect 222528 99368 223396 99396
rect 222528 99356 222534 99368
rect 223390 99356 223396 99368
rect 223448 99356 223454 99408
rect 224126 99356 224132 99408
rect 224184 99396 224190 99408
rect 224862 99396 224868 99408
rect 224184 99368 224868 99396
rect 224184 99356 224190 99368
rect 224862 99356 224868 99368
rect 224920 99356 224926 99408
rect 224954 99356 224960 99408
rect 225012 99396 225018 99408
rect 226242 99396 226248 99408
rect 225012 99368 226248 99396
rect 225012 99356 225018 99368
rect 226242 99356 226248 99368
rect 226300 99356 226306 99408
rect 226610 99356 226616 99408
rect 226668 99396 226674 99408
rect 227622 99396 227628 99408
rect 226668 99368 227628 99396
rect 226668 99356 226674 99368
rect 227622 99356 227628 99368
rect 227680 99356 227686 99408
rect 229094 99356 229100 99408
rect 229152 99396 229158 99408
rect 230290 99396 230296 99408
rect 229152 99368 230296 99396
rect 229152 99356 229158 99368
rect 230290 99356 230296 99368
rect 230348 99356 230354 99408
rect 232406 99356 232412 99408
rect 232464 99396 232470 99408
rect 233142 99396 233148 99408
rect 232464 99368 233148 99396
rect 232464 99356 232470 99368
rect 233142 99356 233148 99368
rect 233200 99356 233206 99408
rect 233234 99356 233240 99408
rect 233292 99396 233298 99408
rect 234430 99396 234436 99408
rect 233292 99368 234436 99396
rect 233292 99356 233298 99368
rect 234430 99356 234436 99368
rect 234488 99356 234494 99408
rect 244734 99356 244740 99408
rect 244792 99396 244798 99408
rect 245562 99396 245568 99408
rect 244792 99368 245568 99396
rect 244792 99356 244798 99368
rect 245562 99356 245568 99368
rect 245620 99356 245626 99408
rect 247218 99356 247224 99408
rect 247276 99396 247282 99408
rect 248230 99396 248236 99408
rect 247276 99368 248236 99396
rect 247276 99356 247282 99368
rect 248230 99356 248236 99368
rect 248288 99356 248294 99408
rect 251358 99356 251364 99408
rect 251416 99396 251422 99408
rect 252462 99396 252468 99408
rect 251416 99368 252468 99396
rect 251416 99356 251422 99368
rect 252462 99356 252468 99368
rect 252520 99356 252526 99408
rect 253014 99356 253020 99408
rect 253072 99396 253078 99408
rect 254578 99396 254584 99408
rect 253072 99368 254584 99396
rect 253072 99356 253078 99368
rect 254578 99356 254584 99368
rect 254636 99356 254642 99408
rect 259638 99356 259644 99408
rect 259696 99396 259702 99408
rect 260742 99396 260748 99408
rect 259696 99368 260748 99396
rect 259696 99356 259702 99368
rect 260742 99356 260748 99368
rect 260800 99356 260806 99408
rect 284386 99356 284392 99408
rect 284444 99396 284450 99408
rect 285582 99396 285588 99408
rect 284444 99368 285588 99396
rect 284444 99356 284450 99368
rect 285582 99356 285588 99368
rect 285640 99356 285646 99408
rect 286042 99356 286048 99408
rect 286100 99396 286106 99408
rect 286870 99396 286876 99408
rect 286100 99368 286876 99396
rect 286100 99356 286106 99368
rect 286870 99356 286876 99368
rect 286928 99356 286934 99408
rect 287606 99356 287612 99408
rect 287664 99396 287670 99408
rect 288342 99396 288348 99408
rect 287664 99368 288348 99396
rect 287664 99356 287670 99368
rect 288342 99356 288348 99368
rect 288400 99356 288406 99408
rect 288434 99356 288440 99408
rect 288492 99396 288498 99408
rect 289722 99396 289728 99408
rect 288492 99368 289728 99396
rect 288492 99356 288498 99368
rect 289722 99356 289728 99368
rect 289780 99356 289786 99408
rect 290090 99356 290096 99408
rect 290148 99396 290154 99408
rect 291010 99396 291016 99408
rect 290148 99368 291016 99396
rect 290148 99356 290154 99368
rect 291010 99356 291016 99368
rect 291068 99356 291074 99408
rect 294230 99356 294236 99408
rect 294288 99396 294294 99408
rect 295242 99396 295248 99408
rect 294288 99368 295248 99396
rect 294288 99356 294294 99368
rect 295242 99356 295248 99368
rect 295300 99356 295306 99408
rect 295886 99356 295892 99408
rect 295944 99396 295950 99408
rect 296622 99396 296628 99408
rect 295944 99368 296628 99396
rect 295944 99356 295950 99368
rect 296622 99356 296628 99368
rect 296680 99356 296686 99408
rect 296714 99356 296720 99408
rect 296772 99396 296778 99408
rect 297910 99396 297916 99408
rect 296772 99368 297916 99396
rect 296772 99356 296778 99368
rect 297910 99356 297916 99368
rect 297968 99356 297974 99408
rect 298370 99356 298376 99408
rect 298428 99396 298434 99408
rect 299290 99396 299296 99408
rect 298428 99368 299296 99396
rect 298428 99356 298434 99368
rect 299290 99356 299296 99368
rect 299348 99356 299354 99408
rect 300854 99356 300860 99408
rect 300912 99396 300918 99408
rect 302050 99396 302056 99408
rect 300912 99368 302056 99396
rect 300912 99356 300918 99368
rect 302050 99356 302056 99368
rect 302108 99356 302114 99408
rect 304166 99356 304172 99408
rect 304224 99396 304230 99408
rect 304902 99396 304908 99408
rect 304224 99368 304908 99396
rect 304224 99356 304230 99368
rect 304902 99356 304908 99368
rect 304960 99356 304966 99408
rect 309134 99356 309140 99408
rect 309192 99396 309198 99408
rect 310422 99396 310428 99408
rect 309192 99368 310428 99396
rect 309192 99356 309198 99368
rect 310422 99356 310428 99368
rect 310480 99356 310486 99408
rect 310698 99356 310704 99408
rect 310756 99396 310762 99408
rect 311802 99396 311808 99408
rect 310756 99368 311808 99396
rect 310756 99356 310762 99368
rect 311802 99356 311808 99368
rect 311860 99356 311866 99408
rect 314838 99356 314844 99408
rect 314896 99396 314902 99408
rect 315850 99396 315856 99408
rect 314896 99368 315856 99396
rect 314896 99356 314902 99368
rect 315850 99356 315856 99368
rect 315908 99356 315914 99408
rect 316494 99356 316500 99408
rect 316552 99396 316558 99408
rect 317230 99396 317236 99408
rect 316552 99368 317236 99396
rect 316552 99356 316558 99368
rect 317230 99356 317236 99368
rect 317288 99356 317294 99408
rect 318978 99356 318984 99408
rect 319036 99396 319042 99408
rect 319990 99396 319996 99408
rect 319036 99368 319996 99396
rect 319036 99356 319042 99368
rect 319990 99356 319996 99368
rect 320048 99356 320054 99408
rect 320634 99356 320640 99408
rect 320692 99396 320698 99408
rect 321462 99396 321468 99408
rect 320692 99368 321468 99396
rect 320692 99356 320698 99368
rect 321462 99356 321468 99368
rect 321520 99356 321526 99408
rect 323118 99356 323124 99408
rect 323176 99396 323182 99408
rect 324222 99396 324228 99408
rect 323176 99368 324228 99396
rect 323176 99356 323182 99368
rect 324222 99356 324228 99368
rect 324280 99356 324286 99408
rect 324774 99356 324780 99408
rect 324832 99396 324838 99408
rect 326338 99396 326344 99408
rect 324832 99368 326344 99396
rect 324832 99356 324838 99368
rect 326338 99356 326344 99368
rect 326396 99356 326402 99408
rect 327258 99356 327264 99408
rect 327316 99396 327322 99408
rect 328270 99396 328276 99408
rect 327316 99368 328276 99396
rect 327316 99356 327322 99368
rect 328270 99356 328276 99368
rect 328328 99356 328334 99408
rect 328914 99356 328920 99408
rect 328972 99396 328978 99408
rect 331858 99396 331864 99408
rect 328972 99368 331864 99396
rect 328972 99356 328978 99368
rect 331858 99356 331864 99368
rect 331916 99356 331922 99408
rect 332962 99356 332968 99408
rect 333020 99396 333026 99408
rect 333790 99396 333796 99408
rect 333020 99368 333796 99396
rect 333020 99356 333026 99368
rect 333790 99356 333796 99368
rect 333848 99356 333854 99408
rect 337102 99356 337108 99408
rect 337160 99396 337166 99408
rect 337930 99396 337936 99408
rect 337160 99368 337936 99396
rect 337160 99356 337166 99368
rect 337930 99356 337936 99368
rect 337988 99356 337994 99408
rect 339586 99356 339592 99408
rect 339644 99396 339650 99408
rect 340782 99396 340788 99408
rect 339644 99368 340788 99396
rect 339644 99356 339650 99368
rect 340782 99356 340788 99368
rect 340840 99356 340846 99408
rect 352006 99356 352012 99408
rect 352064 99396 352070 99408
rect 353110 99396 353116 99408
rect 352064 99368 353116 99396
rect 352064 99356 352070 99368
rect 353110 99356 353116 99368
rect 353168 99356 353174 99408
rect 353662 99356 353668 99408
rect 353720 99396 353726 99408
rect 354490 99396 354496 99408
rect 353720 99368 354496 99396
rect 353720 99356 353726 99368
rect 354490 99356 354496 99368
rect 354548 99356 354554 99408
rect 356054 99356 356060 99408
rect 356112 99396 356118 99408
rect 357250 99396 357256 99408
rect 356112 99368 357256 99396
rect 356112 99356 356118 99368
rect 357250 99356 357256 99368
rect 357308 99356 357314 99408
rect 357710 99356 357716 99408
rect 357768 99396 357774 99408
rect 358722 99396 358728 99408
rect 357768 99368 358728 99396
rect 357768 99356 357774 99368
rect 358722 99356 358728 99368
rect 358780 99356 358786 99408
rect 359366 99356 359372 99408
rect 359424 99396 359430 99408
rect 360102 99396 360108 99408
rect 359424 99368 360108 99396
rect 359424 99356 359430 99368
rect 360102 99356 360108 99368
rect 360160 99356 360166 99408
rect 360194 99356 360200 99408
rect 360252 99396 360258 99408
rect 361482 99396 361488 99408
rect 360252 99368 361488 99396
rect 360252 99356 360258 99368
rect 361482 99356 361488 99368
rect 361540 99356 361546 99408
rect 361850 99356 361856 99408
rect 361908 99396 361914 99408
rect 362770 99396 362776 99408
rect 361908 99368 362776 99396
rect 361908 99356 361914 99368
rect 362770 99356 362776 99368
rect 362828 99356 362834 99408
rect 365990 99356 365996 99408
rect 366048 99396 366054 99408
rect 366910 99396 366916 99408
rect 366048 99368 366916 99396
rect 366048 99356 366054 99368
rect 366910 99356 366916 99368
rect 366968 99356 366974 99408
rect 367646 99356 367652 99408
rect 367704 99396 367710 99408
rect 368382 99396 368388 99408
rect 367704 99368 368388 99396
rect 367704 99356 367710 99368
rect 368382 99356 368388 99368
rect 368440 99356 368446 99408
rect 368474 99356 368480 99408
rect 368532 99396 368538 99408
rect 369670 99396 369676 99408
rect 368532 99368 369676 99396
rect 368532 99356 368538 99368
rect 369670 99356 369676 99368
rect 369728 99356 369734 99408
rect 379974 99356 379980 99408
rect 380032 99396 380038 99408
rect 380710 99396 380716 99408
rect 380032 99368 380716 99396
rect 380032 99356 380038 99368
rect 380710 99356 380716 99368
rect 380768 99356 380774 99408
rect 382458 99356 382464 99408
rect 382516 99396 382522 99408
rect 383562 99396 383568 99408
rect 382516 99368 383568 99396
rect 382516 99356 382522 99368
rect 383562 99356 383568 99368
rect 383620 99356 383626 99408
rect 386598 99356 386604 99408
rect 386656 99396 386662 99408
rect 387610 99396 387616 99408
rect 386656 99368 387616 99396
rect 386656 99356 386662 99368
rect 387610 99356 387616 99368
rect 387668 99356 387674 99408
rect 388254 99356 388260 99408
rect 388312 99396 388318 99408
rect 388990 99396 388996 99408
rect 388312 99368 388996 99396
rect 388312 99356 388318 99368
rect 388990 99356 388996 99368
rect 389048 99356 389054 99408
rect 390738 99356 390744 99408
rect 390796 99396 390802 99408
rect 391750 99396 391756 99408
rect 390796 99368 391756 99396
rect 390796 99356 390802 99368
rect 391750 99356 391756 99368
rect 391808 99356 391814 99408
rect 396534 99356 396540 99408
rect 396592 99396 396598 99408
rect 398098 99396 398104 99408
rect 396592 99368 398104 99396
rect 396592 99356 396598 99368
rect 398098 99356 398104 99368
rect 398156 99356 398162 99408
rect 399018 99356 399024 99408
rect 399076 99396 399082 99408
rect 400122 99396 400128 99408
rect 399076 99368 400128 99396
rect 399076 99356 399082 99368
rect 400122 99356 400128 99368
rect 400180 99356 400186 99408
rect 370866 99328 370872 99340
rect 370827 99300 370872 99328
rect 370866 99288 370872 99300
rect 370924 99288 370930 99340
rect 228266 98744 228272 98796
rect 228324 98784 228330 98796
rect 333974 98784 333980 98796
rect 228324 98756 333980 98784
rect 228324 98744 228330 98756
rect 333974 98744 333980 98756
rect 334032 98744 334038 98796
rect 317322 98676 317328 98728
rect 317380 98716 317386 98728
rect 462314 98716 462320 98728
rect 317380 98688 462320 98716
rect 317380 98676 317386 98688
rect 462314 98676 462320 98688
rect 462372 98676 462378 98728
rect 91370 98608 91376 98660
rect 91428 98648 91434 98660
rect 92382 98648 92388 98660
rect 91428 98620 92388 98648
rect 91428 98608 91434 98620
rect 92382 98608 92388 98620
rect 92440 98608 92446 98660
rect 145834 98608 145840 98660
rect 145892 98648 145898 98660
rect 215294 98648 215300 98660
rect 145892 98620 215300 98648
rect 145892 98608 145898 98620
rect 215294 98608 215300 98620
rect 215352 98608 215358 98660
rect 333698 98608 333704 98660
rect 333756 98648 333762 98660
rect 485774 98648 485780 98660
rect 333756 98620 485780 98648
rect 333756 98608 333762 98620
rect 485774 98608 485780 98620
rect 485832 98608 485838 98660
rect 342070 98580 342076 98592
rect 342031 98552 342076 98580
rect 342070 98540 342076 98552
rect 342128 98540 342134 98592
rect 163130 97316 163136 97368
rect 163188 97356 163194 97368
rect 240134 97356 240140 97368
rect 163188 97328 240140 97356
rect 163188 97316 163194 97328
rect 240134 97316 240140 97328
rect 240192 97316 240198 97368
rect 312354 97316 312360 97368
rect 312412 97356 312418 97368
rect 455414 97356 455420 97368
rect 312412 97328 455420 97356
rect 312412 97316 312418 97328
rect 455414 97316 455420 97328
rect 455472 97316 455478 97368
rect 230750 97248 230756 97300
rect 230808 97288 230814 97300
rect 338114 97288 338120 97300
rect 230808 97260 338120 97288
rect 230808 97248 230814 97260
rect 338114 97248 338120 97260
rect 338172 97248 338178 97300
rect 341242 97248 341248 97300
rect 341300 97288 341306 97300
rect 496814 97288 496820 97300
rect 341300 97260 496820 97288
rect 341300 97248 341306 97260
rect 496814 97248 496820 97260
rect 496872 97248 496878 97300
rect 278498 96704 278504 96756
rect 278556 96744 278562 96756
rect 278682 96744 278688 96756
rect 278556 96716 278688 96744
rect 278556 96704 278562 96716
rect 278682 96704 278688 96716
rect 278740 96704 278746 96756
rect 266998 96608 267004 96620
rect 266959 96580 267004 96608
rect 266998 96568 267004 96580
rect 267056 96568 267062 96620
rect 278593 96611 278651 96617
rect 278593 96577 278605 96611
rect 278639 96608 278651 96611
rect 278682 96608 278688 96620
rect 278639 96580 278688 96608
rect 278639 96577 278651 96580
rect 278593 96571 278651 96577
rect 278682 96568 278688 96580
rect 278740 96568 278746 96620
rect 304994 95956 305000 96008
rect 305052 95996 305058 96008
rect 444374 95996 444380 96008
rect 305052 95968 444380 95996
rect 305052 95956 305058 95968
rect 444374 95956 444380 95968
rect 444432 95956 444438 96008
rect 149974 95888 149980 95940
rect 150032 95928 150038 95940
rect 220814 95928 220820 95940
rect 150032 95900 220820 95928
rect 150032 95888 150038 95900
rect 220814 95888 220820 95900
rect 220872 95888 220878 95940
rect 225782 95888 225788 95940
rect 225840 95928 225846 95940
rect 331214 95928 331220 95940
rect 225840 95900 331220 95928
rect 225840 95888 225846 95900
rect 331214 95888 331220 95900
rect 331272 95888 331278 95940
rect 343726 95888 343732 95940
rect 343784 95928 343790 95940
rect 500954 95928 500960 95940
rect 343784 95900 500960 95928
rect 343784 95888 343790 95900
rect 500954 95888 500960 95900
rect 501012 95888 501018 95940
rect 92106 95276 92112 95328
rect 92164 95316 92170 95328
rect 92164 95288 92336 95316
rect 92164 95276 92170 95288
rect 92308 95260 92336 95288
rect 92290 95208 92296 95260
rect 92348 95208 92354 95260
rect 197998 95248 198004 95260
rect 197959 95220 198004 95248
rect 197998 95208 198004 95220
rect 198056 95208 198062 95260
rect 197998 95112 198004 95124
rect 197959 95084 198004 95112
rect 197998 95072 198004 95084
rect 198056 95072 198062 95124
rect 277762 94596 277768 94648
rect 277820 94636 277826 94648
rect 405734 94636 405740 94648
rect 277820 94608 405740 94636
rect 277820 94596 277826 94608
rect 405734 94596 405740 94608
rect 405792 94596 405798 94648
rect 346210 94528 346216 94580
rect 346268 94568 346274 94580
rect 503714 94568 503720 94580
rect 346268 94540 503720 94568
rect 346268 94528 346274 94540
rect 503714 94528 503720 94540
rect 503772 94528 503778 94580
rect 196066 94460 196072 94512
rect 196124 94500 196130 94512
rect 287054 94500 287060 94512
rect 196124 94472 287060 94500
rect 196124 94460 196130 94472
rect 287054 94460 287060 94472
rect 287112 94460 287118 94512
rect 394878 94460 394884 94512
rect 394936 94500 394942 94512
rect 574094 94500 574100 94512
rect 394936 94472 574100 94500
rect 394936 94460 394942 94472
rect 574094 94460 574100 94472
rect 574152 94460 574158 94512
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 79686 93820 79692 93832
rect 3476 93792 79692 93820
rect 3476 93780 3482 93792
rect 79686 93780 79692 93792
rect 79744 93780 79750 93832
rect 295058 93168 295064 93220
rect 295116 93208 295122 93220
rect 430574 93208 430580 93220
rect 295116 93180 430580 93208
rect 295116 93168 295122 93180
rect 430574 93168 430580 93180
rect 430632 93168 430638 93220
rect 147490 93100 147496 93152
rect 147548 93140 147554 93152
rect 218054 93140 218060 93152
rect 147548 93112 218060 93140
rect 147548 93100 147554 93112
rect 218054 93100 218060 93112
rect 218112 93100 218118 93152
rect 219250 93100 219256 93152
rect 219308 93140 219314 93152
rect 320174 93140 320180 93152
rect 219308 93112 320180 93140
rect 219308 93100 219314 93112
rect 320174 93100 320180 93112
rect 320232 93100 320238 93152
rect 354490 93100 354496 93152
rect 354548 93140 354554 93152
rect 514754 93140 514760 93152
rect 354548 93112 514760 93140
rect 354548 93100 354554 93112
rect 514754 93100 514760 93112
rect 514812 93100 514818 93152
rect 153102 91808 153108 91860
rect 153160 91848 153166 91860
rect 224954 91848 224960 91860
rect 153160 91820 224960 91848
rect 153160 91808 153166 91820
rect 224954 91808 224960 91820
rect 225012 91808 225018 91860
rect 291010 91808 291016 91860
rect 291068 91848 291074 91860
rect 423674 91848 423680 91860
rect 291068 91820 423680 91848
rect 291068 91808 291074 91820
rect 423674 91808 423680 91820
rect 423732 91808 423738 91860
rect 216582 91740 216588 91792
rect 216640 91780 216646 91792
rect 316034 91780 316040 91792
rect 216640 91752 316040 91780
rect 216640 91740 216646 91752
rect 316034 91740 316040 91752
rect 316092 91740 316098 91792
rect 357250 91740 357256 91792
rect 357308 91780 357314 91792
rect 518894 91780 518900 91792
rect 357308 91752 518900 91780
rect 357308 91740 357314 91752
rect 518894 91740 518900 91752
rect 518952 91740 518958 91792
rect 155770 90380 155776 90432
rect 155828 90420 155834 90432
rect 227714 90420 227720 90432
rect 155828 90392 227720 90420
rect 155828 90380 155834 90392
rect 227714 90380 227720 90392
rect 227772 90380 227778 90432
rect 285490 90380 285496 90432
rect 285548 90420 285554 90432
rect 416774 90420 416780 90432
rect 285548 90392 416780 90420
rect 285548 90380 285554 90392
rect 416774 90380 416780 90392
rect 416832 90380 416838 90432
rect 213730 90312 213736 90364
rect 213788 90352 213794 90364
rect 313274 90352 313280 90364
rect 213788 90324 313280 90352
rect 213788 90312 213794 90324
rect 313274 90312 313280 90324
rect 313332 90312 313338 90364
rect 358538 90312 358544 90364
rect 358596 90352 358602 90364
rect 521654 90352 521660 90364
rect 358596 90324 521660 90352
rect 358596 90312 358602 90324
rect 521654 90312 521660 90324
rect 521712 90312 521718 90364
rect 92198 89740 92204 89752
rect 92159 89712 92204 89740
rect 92198 89700 92204 89712
rect 92256 89700 92262 89752
rect 151446 89700 151452 89752
rect 151504 89740 151510 89752
rect 151630 89740 151636 89752
rect 151504 89712 151636 89740
rect 151504 89700 151510 89712
rect 151630 89700 151636 89712
rect 151688 89700 151694 89752
rect 198550 89740 198556 89752
rect 198511 89712 198556 89740
rect 198550 89700 198556 89712
rect 198608 89700 198614 89752
rect 227438 89740 227444 89752
rect 227399 89712 227444 89740
rect 227438 89700 227444 89712
rect 227496 89700 227502 89752
rect 274358 89700 274364 89752
rect 274416 89740 274422 89752
rect 274542 89740 274548 89752
rect 274416 89712 274548 89740
rect 274416 89700 274422 89712
rect 274542 89700 274548 89712
rect 274600 89700 274606 89752
rect 266998 89672 267004 89684
rect 266959 89644 267004 89672
rect 266998 89632 267004 89644
rect 267056 89632 267062 89684
rect 282730 89088 282736 89140
rect 282788 89128 282794 89140
rect 412634 89128 412640 89140
rect 282788 89100 412640 89128
rect 282788 89088 282794 89100
rect 412634 89088 412640 89100
rect 412692 89088 412698 89140
rect 158530 89020 158536 89072
rect 158588 89060 158594 89072
rect 231854 89060 231860 89072
rect 158588 89032 231860 89060
rect 158588 89020 158594 89032
rect 231854 89020 231860 89032
rect 231912 89020 231918 89072
rect 299290 89020 299296 89072
rect 299348 89060 299354 89072
rect 434714 89060 434720 89072
rect 299348 89032 434720 89060
rect 299348 89020 299354 89032
rect 434714 89020 434720 89032
rect 434772 89020 434778 89072
rect 210970 88952 210976 89004
rect 211028 88992 211034 89004
rect 307754 88992 307760 89004
rect 211028 88964 307760 88992
rect 211028 88952 211034 88964
rect 307754 88952 307760 88964
rect 307812 88952 307818 89004
rect 364242 88952 364248 89004
rect 364300 88992 364306 89004
rect 528554 88992 528560 89004
rect 364300 88964 528560 88992
rect 364300 88952 364306 88964
rect 528554 88952 528560 88964
rect 528612 88952 528618 89004
rect 402514 88272 402520 88324
rect 402572 88312 402578 88324
rect 580166 88312 580172 88324
rect 402572 88284 580172 88312
rect 402572 88272 402578 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 146110 87660 146116 87712
rect 146168 87700 146174 87712
rect 213914 87700 213920 87712
rect 146168 87672 213920 87700
rect 146168 87660 146174 87672
rect 213914 87660 213920 87672
rect 213972 87660 213978 87712
rect 264790 87660 264796 87712
rect 264848 87700 264854 87712
rect 385034 87700 385040 87712
rect 264848 87672 385040 87700
rect 264848 87660 264854 87672
rect 385034 87660 385040 87672
rect 385092 87660 385098 87712
rect 187602 87592 187608 87644
rect 187660 87632 187666 87644
rect 274634 87632 274640 87644
rect 187660 87604 274640 87632
rect 187660 87592 187666 87604
rect 274634 87592 274640 87604
rect 274692 87592 274698 87644
rect 277210 87592 277216 87644
rect 277268 87632 277274 87644
rect 404354 87632 404360 87644
rect 277268 87604 404360 87632
rect 277268 87592 277274 87604
rect 404354 87592 404360 87604
rect 404412 87592 404418 87644
rect 104618 86980 104624 87032
rect 104676 87020 104682 87032
rect 104710 87020 104716 87032
rect 104676 86992 104716 87020
rect 104676 86980 104682 86992
rect 104710 86980 104716 86992
rect 104768 86980 104774 87032
rect 227438 87020 227444 87032
rect 227399 86992 227444 87020
rect 227438 86980 227444 86992
rect 227496 86980 227502 87032
rect 239858 86980 239864 87032
rect 239916 87020 239922 87032
rect 239950 87020 239956 87032
rect 239916 86992 239956 87020
rect 239916 86980 239922 86992
rect 239950 86980 239956 86992
rect 240008 86980 240014 87032
rect 278590 87020 278596 87032
rect 278551 86992 278596 87020
rect 278590 86980 278596 86992
rect 278648 86980 278654 87032
rect 342070 87020 342076 87032
rect 342031 86992 342076 87020
rect 342070 86980 342076 86992
rect 342128 86980 342134 87032
rect 309778 86368 309784 86420
rect 309836 86408 309842 86420
rect 427814 86408 427820 86420
rect 309836 86380 427820 86408
rect 309836 86368 309842 86380
rect 427814 86368 427820 86380
rect 427872 86368 427878 86420
rect 281350 86300 281356 86352
rect 281408 86340 281414 86352
rect 408494 86340 408500 86352
rect 281408 86312 408500 86340
rect 281408 86300 281414 86312
rect 408494 86300 408500 86312
rect 408552 86300 408558 86352
rect 143350 86232 143356 86284
rect 143408 86272 143414 86284
rect 209774 86272 209780 86284
rect 143408 86244 209780 86272
rect 143408 86232 143414 86244
rect 209774 86232 209780 86244
rect 209832 86232 209838 86284
rect 211062 86232 211068 86284
rect 211120 86272 211126 86284
rect 309134 86272 309140 86284
rect 211120 86244 309140 86272
rect 211120 86232 211126 86244
rect 309134 86232 309140 86244
rect 309192 86232 309198 86284
rect 366910 86232 366916 86284
rect 366968 86272 366974 86284
rect 532694 86272 532700 86284
rect 366968 86244 532700 86272
rect 366968 86232 366974 86244
rect 532694 86232 532700 86244
rect 532752 86232 532758 86284
rect 92198 85592 92204 85604
rect 92159 85564 92204 85592
rect 92198 85552 92204 85564
rect 92256 85552 92262 85604
rect 96338 85552 96344 85604
rect 96396 85592 96402 85604
rect 96430 85592 96436 85604
rect 96396 85564 96436 85592
rect 96396 85552 96402 85564
rect 96430 85552 96436 85564
rect 96488 85552 96494 85604
rect 198001 85595 198059 85601
rect 198001 85561 198013 85595
rect 198047 85592 198059 85595
rect 198090 85592 198096 85604
rect 198047 85564 198096 85592
rect 198047 85561 198059 85564
rect 198001 85555 198059 85561
rect 198090 85552 198096 85564
rect 198148 85552 198154 85604
rect 198550 85592 198556 85604
rect 198511 85564 198556 85592
rect 198550 85552 198556 85564
rect 198608 85552 198614 85604
rect 518894 85524 518900 85536
rect 518855 85496 518900 85524
rect 518894 85484 518900 85496
rect 518952 85484 518958 85536
rect 532694 85524 532700 85536
rect 532655 85496 532700 85524
rect 532694 85484 532700 85496
rect 532752 85484 532758 85536
rect 275922 84940 275928 84992
rect 275980 84980 275986 84992
rect 401594 84980 401600 84992
rect 275980 84952 401600 84980
rect 275980 84940 275986 84952
rect 401594 84940 401600 84952
rect 401652 84940 401658 84992
rect 289722 84872 289728 84924
rect 289780 84912 289786 84924
rect 420914 84912 420920 84924
rect 289780 84884 420920 84912
rect 289780 84872 289786 84884
rect 420914 84872 420920 84884
rect 420972 84872 420978 84924
rect 209590 84804 209596 84856
rect 209648 84844 209654 84856
rect 304994 84844 305000 84856
rect 209648 84816 305000 84844
rect 209648 84804 209654 84816
rect 304994 84804 305000 84816
rect 305052 84804 305058 84856
rect 369670 84804 369676 84856
rect 369728 84844 369734 84856
rect 536834 84844 536840 84856
rect 369728 84816 536840 84844
rect 369728 84804 369734 84816
rect 536834 84804 536840 84816
rect 536892 84804 536898 84856
rect 273070 83512 273076 83564
rect 273128 83552 273134 83564
rect 398834 83552 398840 83564
rect 273128 83524 398840 83552
rect 273128 83512 273134 83524
rect 398834 83512 398840 83524
rect 398892 83512 398898 83564
rect 400030 83512 400036 83564
rect 400088 83552 400094 83564
rect 482278 83552 482284 83564
rect 400088 83524 482284 83552
rect 400088 83512 400094 83524
rect 482278 83512 482284 83524
rect 482336 83512 482342 83564
rect 206830 83444 206836 83496
rect 206888 83484 206894 83496
rect 302234 83484 302240 83496
rect 206888 83456 302240 83484
rect 206888 83444 206894 83456
rect 302234 83444 302240 83456
rect 302292 83444 302298 83496
rect 370682 83444 370688 83496
rect 370740 83484 370746 83496
rect 539594 83484 539600 83496
rect 370740 83456 539600 83484
rect 370740 83444 370746 83456
rect 539594 83444 539600 83456
rect 539652 83444 539658 83496
rect 140682 82152 140688 82204
rect 140740 82192 140746 82204
rect 207014 82192 207020 82204
rect 140740 82164 207020 82192
rect 140740 82152 140746 82164
rect 207014 82152 207020 82164
rect 207072 82152 207078 82204
rect 315850 82152 315856 82204
rect 315908 82192 315914 82204
rect 459646 82192 459652 82204
rect 315908 82164 459652 82192
rect 315908 82152 315914 82164
rect 459646 82152 459652 82164
rect 459704 82152 459710 82204
rect 104618 82124 104624 82136
rect 104579 82096 104624 82124
rect 104618 82084 104624 82096
rect 104676 82084 104682 82136
rect 175182 82084 175188 82136
rect 175240 82124 175246 82136
rect 256694 82124 256700 82136
rect 175240 82096 256700 82124
rect 175240 82084 175246 82096
rect 256694 82084 256700 82096
rect 256752 82084 256758 82136
rect 257890 82084 257896 82136
rect 257948 82124 257954 82136
rect 375374 82124 375380 82136
rect 257948 82096 375380 82124
rect 257948 82084 257954 82096
rect 375374 82084 375380 82096
rect 375432 82084 375438 82136
rect 381538 82084 381544 82136
rect 381596 82124 381602 82136
rect 550634 82124 550640 82136
rect 381596 82096 550640 82124
rect 381596 82084 381602 82096
rect 550634 82084 550640 82096
rect 550692 82084 550698 82136
rect 227070 82016 227076 82068
rect 227128 82056 227134 82068
rect 227438 82056 227444 82068
rect 227128 82028 227444 82056
rect 227128 82016 227134 82028
rect 227438 82016 227444 82028
rect 227496 82016 227502 82068
rect 341702 82016 341708 82068
rect 341760 82056 341766 82068
rect 342070 82056 342076 82068
rect 341760 82028 342076 82056
rect 341760 82016 341766 82028
rect 342070 82016 342076 82028
rect 342128 82016 342134 82068
rect 239858 81852 239864 81864
rect 239819 81824 239864 81852
rect 239858 81812 239864 81824
rect 239916 81812 239922 81864
rect 266170 80792 266176 80844
rect 266228 80832 266234 80844
rect 387794 80832 387800 80844
rect 266228 80804 387800 80832
rect 266228 80792 266234 80804
rect 387794 80792 387800 80804
rect 387852 80792 387858 80844
rect 91922 80724 91928 80776
rect 91980 80764 91986 80776
rect 92201 80767 92259 80773
rect 92201 80764 92213 80767
rect 91980 80736 92213 80764
rect 91980 80724 91986 80736
rect 92201 80733 92213 80736
rect 92247 80733 92259 80767
rect 92201 80727 92259 80733
rect 277302 80724 277308 80776
rect 277360 80764 277366 80776
rect 402974 80764 402980 80776
rect 277360 80736 402980 80764
rect 277360 80724 277366 80736
rect 402974 80724 402980 80736
rect 403032 80724 403038 80776
rect 137830 80656 137836 80708
rect 137888 80696 137894 80708
rect 202874 80696 202880 80708
rect 137888 80668 202880 80696
rect 137888 80656 137894 80668
rect 202874 80656 202880 80668
rect 202932 80656 202938 80708
rect 204162 80656 204168 80708
rect 204220 80696 204226 80708
rect 298094 80696 298100 80708
rect 204220 80668 298100 80696
rect 204220 80656 204226 80668
rect 298094 80656 298100 80668
rect 298152 80656 298158 80708
rect 385678 80656 385684 80708
rect 385736 80696 385742 80708
rect 557534 80696 557540 80708
rect 385736 80668 557540 80696
rect 385736 80656 385742 80668
rect 557534 80656 557540 80668
rect 557592 80656 557598 80708
rect 198001 80223 198059 80229
rect 198001 80189 198013 80223
rect 198047 80220 198059 80223
rect 198090 80220 198096 80232
rect 198047 80192 198096 80220
rect 198047 80189 198059 80192
rect 198001 80183 198059 80189
rect 198090 80180 198096 80192
rect 198148 80180 198154 80232
rect 267090 80152 267096 80164
rect 267051 80124 267096 80152
rect 267090 80112 267096 80124
rect 267148 80112 267154 80164
rect 278590 80044 278596 80096
rect 278648 80044 278654 80096
rect 278608 79948 278636 80044
rect 278682 79948 278688 79960
rect 278608 79920 278688 79948
rect 278682 79908 278688 79920
rect 278740 79908 278746 79960
rect 3510 79432 3516 79484
rect 3568 79472 3574 79484
rect 8938 79472 8944 79484
rect 3568 79444 8944 79472
rect 3568 79432 3574 79444
rect 8938 79432 8944 79444
rect 8996 79432 9002 79484
rect 201310 79364 201316 79416
rect 201368 79404 201374 79416
rect 295334 79404 295340 79416
rect 201368 79376 295340 79404
rect 201368 79364 201374 79376
rect 295334 79364 295340 79376
rect 295392 79364 295398 79416
rect 329742 79364 329748 79416
rect 329800 79404 329806 79416
rect 480254 79404 480260 79416
rect 329800 79376 480260 79404
rect 329800 79364 329806 79376
rect 480254 79364 480260 79376
rect 480312 79364 480318 79416
rect 135070 79296 135076 79348
rect 135128 79336 135134 79348
rect 200114 79336 200120 79348
rect 135128 79308 200120 79336
rect 135128 79296 135134 79308
rect 200114 79296 200120 79308
rect 200172 79296 200178 79348
rect 263502 79296 263508 79348
rect 263560 79336 263566 79348
rect 383654 79336 383660 79348
rect 263560 79308 383660 79336
rect 263560 79296 263566 79308
rect 383654 79296 383660 79308
rect 383712 79296 383718 79348
rect 388990 79296 388996 79348
rect 389048 79336 389054 79348
rect 564434 79336 564440 79348
rect 389048 79308 564440 79336
rect 389048 79296 389054 79308
rect 564434 79296 564440 79308
rect 564492 79296 564498 79348
rect 198550 78004 198556 78056
rect 198608 78044 198614 78056
rect 291194 78044 291200 78056
rect 198608 78016 291200 78044
rect 198608 78004 198614 78016
rect 291194 78004 291200 78016
rect 291252 78004 291258 78056
rect 307662 78004 307668 78056
rect 307720 78044 307726 78056
rect 448514 78044 448520 78056
rect 307720 78016 448520 78044
rect 307720 78004 307726 78016
rect 448514 78004 448520 78016
rect 448572 78004 448578 78056
rect 133782 77936 133788 77988
rect 133840 77976 133846 77988
rect 195974 77976 195980 77988
rect 133840 77948 195980 77976
rect 133840 77936 133846 77948
rect 195974 77936 195980 77948
rect 196032 77936 196038 77988
rect 260650 77936 260656 77988
rect 260708 77976 260714 77988
rect 380894 77976 380900 77988
rect 260708 77948 380900 77976
rect 260708 77936 260714 77948
rect 380894 77936 380900 77948
rect 380952 77936 380958 77988
rect 391750 77936 391756 77988
rect 391808 77976 391814 77988
rect 568574 77976 568580 77988
rect 391808 77948 568580 77976
rect 391808 77936 391814 77948
rect 568574 77936 568580 77948
rect 568632 77936 568638 77988
rect 104618 77364 104624 77376
rect 104579 77336 104624 77364
rect 104618 77324 104624 77336
rect 104676 77324 104682 77376
rect 239858 77364 239864 77376
rect 239819 77336 239864 77364
rect 239858 77324 239864 77336
rect 239916 77324 239922 77376
rect 267090 77296 267096 77308
rect 267051 77268 267096 77296
rect 267090 77256 267096 77268
rect 267148 77256 267154 77308
rect 104526 77228 104532 77240
rect 104487 77200 104532 77228
rect 104526 77188 104532 77200
rect 104584 77188 104590 77240
rect 151538 77228 151544 77240
rect 151499 77200 151544 77228
rect 151538 77188 151544 77200
rect 151596 77188 151602 77240
rect 239766 77228 239772 77240
rect 239727 77200 239772 77228
rect 239766 77188 239772 77200
rect 239824 77188 239830 77240
rect 402422 77188 402428 77240
rect 402480 77228 402486 77240
rect 580166 77228 580172 77240
rect 402480 77200 580172 77228
rect 402480 77188 402486 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 254578 76576 254584 76628
rect 254636 76616 254642 76628
rect 369854 76616 369860 76628
rect 254636 76588 369860 76616
rect 254636 76576 254642 76588
rect 369854 76576 369860 76588
rect 369912 76576 369918 76628
rect 131022 76508 131028 76560
rect 131080 76548 131086 76560
rect 193214 76548 193220 76560
rect 131080 76520 193220 76548
rect 131080 76508 131086 76520
rect 193214 76508 193220 76520
rect 193272 76508 193278 76560
rect 194410 76508 194416 76560
rect 194468 76548 194474 76560
rect 284294 76548 284300 76560
rect 194468 76520 284300 76548
rect 194468 76508 194474 76520
rect 284294 76508 284300 76520
rect 284352 76508 284358 76560
rect 304258 76508 304264 76560
rect 304316 76548 304322 76560
rect 441614 76548 441620 76560
rect 304316 76520 441620 76548
rect 304316 76508 304322 76520
rect 441614 76508 441620 76520
rect 441672 76508 441678 76560
rect 197998 75936 198004 75948
rect 197959 75908 198004 75936
rect 197998 75896 198004 75908
rect 198056 75896 198062 75948
rect 518894 75936 518900 75948
rect 518855 75908 518900 75936
rect 518894 75896 518900 75908
rect 518952 75896 518958 75948
rect 532694 75936 532700 75948
rect 532655 75908 532700 75936
rect 532694 75896 532700 75908
rect 532752 75896 532758 75948
rect 191742 75216 191748 75268
rect 191800 75256 191806 75268
rect 280154 75256 280160 75268
rect 191800 75228 280160 75256
rect 191800 75216 191806 75228
rect 280154 75216 280160 75228
rect 280212 75216 280218 75268
rect 300762 75216 300768 75268
rect 300820 75256 300826 75268
rect 437474 75256 437480 75268
rect 300820 75228 437480 75256
rect 300820 75216 300826 75228
rect 437474 75216 437480 75228
rect 437532 75216 437538 75268
rect 128262 75148 128268 75200
rect 128320 75188 128326 75200
rect 189074 75188 189080 75200
rect 128320 75160 189080 75188
rect 128320 75148 128326 75160
rect 189074 75148 189080 75160
rect 189132 75148 189138 75200
rect 245470 75148 245476 75200
rect 245528 75188 245534 75200
rect 358814 75188 358820 75200
rect 245528 75160 358820 75188
rect 245528 75148 245534 75160
rect 358814 75148 358820 75160
rect 358872 75148 358878 75200
rect 393222 75148 393228 75200
rect 393280 75188 393286 75200
rect 571334 75188 571340 75200
rect 393280 75160 571340 75188
rect 393280 75148 393286 75160
rect 571334 75148 571340 75160
rect 571392 75148 571398 75200
rect 215018 74468 215024 74520
rect 215076 74508 215082 74520
rect 215202 74508 215208 74520
rect 215076 74480 215208 74508
rect 215076 74468 215082 74480
rect 215202 74468 215208 74480
rect 215260 74468 215266 74520
rect 188890 73856 188896 73908
rect 188948 73896 188954 73908
rect 277394 73896 277400 73908
rect 188948 73868 277400 73896
rect 188948 73856 188954 73868
rect 277394 73856 277400 73868
rect 277452 73856 277458 73908
rect 300118 73856 300124 73908
rect 300176 73896 300182 73908
rect 426434 73896 426440 73908
rect 300176 73868 426440 73896
rect 300176 73856 300182 73868
rect 426434 73856 426440 73868
rect 426492 73856 426498 73908
rect 244090 73788 244096 73840
rect 244148 73828 244154 73840
rect 356054 73828 356060 73840
rect 244148 73800 356060 73828
rect 244148 73788 244154 73800
rect 356054 73788 356060 73800
rect 356112 73788 356118 73840
rect 395982 73788 395988 73840
rect 396040 73828 396046 73840
rect 575474 73828 575480 73840
rect 396040 73800 575480 73828
rect 396040 73788 396046 73800
rect 575474 73788 575480 73800
rect 575532 73788 575538 73840
rect 186130 72496 186136 72548
rect 186188 72536 186194 72548
rect 273254 72536 273260 72548
rect 186188 72508 273260 72536
rect 186188 72496 186194 72508
rect 273254 72496 273260 72508
rect 273312 72496 273318 72548
rect 282822 72496 282828 72548
rect 282880 72536 282886 72548
rect 411254 72536 411260 72548
rect 282880 72508 411260 72536
rect 282880 72496 282886 72508
rect 411254 72496 411260 72508
rect 411312 72496 411318 72548
rect 224862 72428 224868 72480
rect 224920 72468 224926 72480
rect 328454 72468 328460 72480
rect 224920 72440 328460 72468
rect 224920 72428 224926 72440
rect 328454 72428 328460 72440
rect 328512 72428 328518 72480
rect 375190 72428 375196 72480
rect 375248 72468 375254 72480
rect 545114 72468 545120 72480
rect 375248 72440 545120 72468
rect 375248 72428 375254 72440
rect 545114 72428 545120 72440
rect 545172 72428 545178 72480
rect 274542 71176 274548 71188
rect 274503 71148 274548 71176
rect 274542 71136 274548 71148
rect 274600 71136 274606 71188
rect 285582 71136 285588 71188
rect 285640 71176 285646 71188
rect 415394 71176 415400 71188
rect 285640 71148 415400 71176
rect 285640 71136 285646 71148
rect 415394 71136 415400 71148
rect 415452 71136 415458 71188
rect 186958 71068 186964 71120
rect 187016 71108 187022 71120
rect 270494 71108 270500 71120
rect 187016 71080 270500 71108
rect 187016 71068 187022 71080
rect 270494 71068 270500 71080
rect 270552 71068 270558 71120
rect 303522 71068 303528 71120
rect 303580 71108 303586 71120
rect 442994 71108 443000 71120
rect 303580 71080 443000 71108
rect 303580 71068 303586 71080
rect 442994 71068 443000 71080
rect 443052 71068 443058 71120
rect 125410 71000 125416 71052
rect 125468 71040 125474 71052
rect 184934 71040 184940 71052
rect 125468 71012 184940 71040
rect 125468 71000 125474 71012
rect 184934 71000 184940 71012
rect 184992 71000 184998 71052
rect 219342 71000 219348 71052
rect 219400 71040 219406 71052
rect 321554 71040 321560 71052
rect 219400 71012 321560 71040
rect 219400 71000 219406 71012
rect 321554 71000 321560 71012
rect 321612 71000 321618 71052
rect 377950 71000 377956 71052
rect 378008 71040 378014 71052
rect 547874 71040 547880 71052
rect 378008 71012 547880 71040
rect 378008 71000 378014 71012
rect 547874 71000 547880 71012
rect 547932 71000 547938 71052
rect 227346 70496 227352 70508
rect 227272 70468 227352 70496
rect 227272 70372 227300 70468
rect 227346 70456 227352 70468
rect 227404 70456 227410 70508
rect 341978 70496 341984 70508
rect 341904 70468 341984 70496
rect 267090 70428 267096 70440
rect 267051 70400 267096 70428
rect 267090 70388 267096 70400
rect 267148 70388 267154 70440
rect 341904 70372 341932 70468
rect 341978 70456 341984 70468
rect 342036 70456 342042 70508
rect 227254 70320 227260 70372
rect 227312 70320 227318 70372
rect 341886 70320 341892 70372
rect 341944 70320 341950 70372
rect 182818 69776 182824 69828
rect 182876 69816 182882 69828
rect 266354 69816 266360 69828
rect 182876 69788 266360 69816
rect 182876 69776 182882 69788
rect 266354 69776 266360 69788
rect 266412 69776 266418 69828
rect 209682 69708 209688 69760
rect 209740 69748 209746 69760
rect 306374 69748 306380 69760
rect 209740 69720 306380 69748
rect 209740 69708 209746 69720
rect 306374 69708 306380 69720
rect 306432 69708 306438 69760
rect 322198 69708 322204 69760
rect 322256 69748 322262 69760
rect 422294 69748 422300 69760
rect 322256 69720 422300 69748
rect 322256 69708 322262 69720
rect 422294 69708 422300 69720
rect 422352 69708 422358 69760
rect 122650 69640 122656 69692
rect 122708 69680 122714 69692
rect 182174 69680 182180 69692
rect 122708 69652 182180 69680
rect 122708 69640 122714 69652
rect 182174 69640 182180 69652
rect 182232 69640 182238 69692
rect 256602 69640 256608 69692
rect 256660 69680 256666 69692
rect 373994 69680 374000 69692
rect 256660 69652 374000 69680
rect 256660 69640 256666 69652
rect 373994 69640 374000 69652
rect 374052 69640 374058 69692
rect 382182 69640 382188 69692
rect 382240 69680 382246 69692
rect 554774 69680 554780 69692
rect 382240 69652 554780 69680
rect 382240 69640 382246 69652
rect 554774 69640 554780 69652
rect 554832 69640 554838 69692
rect 292482 68416 292488 68468
rect 292540 68456 292546 68468
rect 425054 68456 425060 68468
rect 292540 68428 425060 68456
rect 292540 68416 292546 68428
rect 425054 68416 425060 68428
rect 425112 68416 425118 68468
rect 179322 68348 179328 68400
rect 179380 68388 179386 68400
rect 262214 68388 262220 68400
rect 179380 68360 262220 68388
rect 179380 68348 179386 68360
rect 262214 68348 262220 68360
rect 262272 68348 262278 68400
rect 302050 68348 302056 68400
rect 302108 68388 302114 68400
rect 438854 68388 438860 68400
rect 302108 68360 438860 68388
rect 302108 68348 302114 68360
rect 438854 68348 438860 68360
rect 438912 68348 438918 68400
rect 121270 68280 121276 68332
rect 121328 68320 121334 68332
rect 178034 68320 178040 68332
rect 121328 68292 178040 68320
rect 121328 68280 121334 68292
rect 178034 68280 178040 68292
rect 178092 68280 178098 68332
rect 215938 68280 215944 68332
rect 215996 68320 216002 68332
rect 313366 68320 313372 68332
rect 215996 68292 313372 68320
rect 215996 68280 216002 68292
rect 313366 68280 313372 68292
rect 313424 68280 313430 68332
rect 387610 68280 387616 68332
rect 387668 68320 387674 68332
rect 563054 68320 563060 68332
rect 387668 68292 563060 68320
rect 387668 68280 387674 68292
rect 563054 68280 563060 68292
rect 563112 68280 563118 68332
rect 92201 67643 92259 67649
rect 92201 67609 92213 67643
rect 92247 67640 92259 67643
rect 92290 67640 92296 67652
rect 92247 67612 92296 67640
rect 92247 67609 92259 67612
rect 92201 67603 92259 67609
rect 92290 67600 92296 67612
rect 92348 67600 92354 67652
rect 104529 67643 104587 67649
rect 104529 67609 104541 67643
rect 104575 67640 104587 67643
rect 104618 67640 104624 67652
rect 104575 67612 104624 67640
rect 104575 67609 104587 67612
rect 104529 67603 104587 67609
rect 104618 67600 104624 67612
rect 104676 67600 104682 67652
rect 151541 67643 151599 67649
rect 151541 67609 151553 67643
rect 151587 67640 151599 67643
rect 151630 67640 151636 67652
rect 151587 67612 151636 67640
rect 151587 67609 151599 67612
rect 151541 67603 151599 67609
rect 151630 67600 151636 67612
rect 151688 67600 151694 67652
rect 239769 67643 239827 67649
rect 239769 67609 239781 67643
rect 239815 67640 239827 67643
rect 239858 67640 239864 67652
rect 239815 67612 239864 67640
rect 239815 67609 239827 67612
rect 239769 67603 239827 67609
rect 239858 67600 239864 67612
rect 239916 67600 239922 67652
rect 267090 67640 267096 67652
rect 267051 67612 267096 67640
rect 267090 67600 267096 67612
rect 267148 67600 267154 67652
rect 274542 67640 274548 67652
rect 274503 67612 274548 67640
rect 274542 67600 274548 67612
rect 274600 67600 274606 67652
rect 550634 67600 550640 67652
rect 550692 67640 550698 67652
rect 550910 67640 550916 67652
rect 550692 67612 550916 67640
rect 550692 67600 550698 67612
rect 550910 67600 550916 67612
rect 550968 67600 550974 67652
rect 151446 67464 151452 67516
rect 151504 67504 151510 67516
rect 151630 67504 151636 67516
rect 151504 67476 151636 67504
rect 151504 67464 151510 67476
rect 151630 67464 151636 67476
rect 151688 67464 151694 67516
rect 274358 67464 274364 67516
rect 274416 67504 274422 67516
rect 274542 67504 274548 67516
rect 274416 67476 274548 67504
rect 274416 67464 274422 67476
rect 274542 67464 274548 67476
rect 274600 67464 274606 67516
rect 278590 66988 278596 67040
rect 278648 67028 278654 67040
rect 407114 67028 407120 67040
rect 278648 67000 407120 67028
rect 278648 66988 278654 67000
rect 407114 66988 407120 67000
rect 407172 66988 407178 67040
rect 176470 66920 176476 66972
rect 176528 66960 176534 66972
rect 259454 66960 259460 66972
rect 176528 66932 259460 66960
rect 176528 66920 176534 66932
rect 259454 66920 259460 66932
rect 259512 66920 259518 66972
rect 295242 66920 295248 66972
rect 295300 66960 295306 66972
rect 429194 66960 429200 66972
rect 295300 66932 429200 66960
rect 295300 66920 295306 66932
rect 429194 66920 429200 66932
rect 429252 66920 429258 66972
rect 118510 66852 118516 66904
rect 118568 66892 118574 66904
rect 175274 66892 175280 66904
rect 118568 66864 175280 66892
rect 118568 66852 118574 66864
rect 175274 66852 175280 66864
rect 175332 66852 175338 66904
rect 212442 66852 212448 66904
rect 212500 66892 212506 66904
rect 310514 66892 310520 66904
rect 212500 66864 310520 66892
rect 212500 66852 212506 66864
rect 310514 66852 310520 66864
rect 310572 66852 310578 66904
rect 389082 66852 389088 66904
rect 389140 66892 389146 66904
rect 565814 66892 565820 66904
rect 389140 66864 565820 66892
rect 389140 66852 389146 66864
rect 565814 66852 565820 66864
rect 565872 66852 565878 66904
rect 96249 66215 96307 66221
rect 96249 66181 96261 66215
rect 96295 66212 96307 66215
rect 96338 66212 96344 66224
rect 96295 66184 96344 66212
rect 96295 66181 96307 66184
rect 96249 66175 96307 66181
rect 96338 66172 96344 66184
rect 96396 66172 96402 66224
rect 200114 66212 200120 66224
rect 200075 66184 200120 66212
rect 200114 66172 200120 66184
rect 200172 66172 200178 66224
rect 227254 66172 227260 66224
rect 227312 66212 227318 66224
rect 227438 66212 227444 66224
rect 227312 66184 227444 66212
rect 227312 66172 227318 66184
rect 227438 66172 227444 66184
rect 227496 66172 227502 66224
rect 341886 66212 341892 66224
rect 341847 66184 341892 66212
rect 341886 66172 341892 66184
rect 341944 66172 341950 66224
rect 518894 66212 518900 66224
rect 518855 66184 518900 66212
rect 518894 66172 518900 66184
rect 518952 66172 518958 66224
rect 532694 66212 532700 66224
rect 532655 66184 532700 66212
rect 532694 66172 532700 66184
rect 532752 66172 532758 66224
rect 268930 65628 268936 65680
rect 268988 65668 268994 65680
rect 391934 65668 391940 65680
rect 268988 65640 391940 65668
rect 268988 65628 268994 65640
rect 391934 65628 391940 65640
rect 391992 65628 391998 65680
rect 173710 65560 173716 65612
rect 173768 65600 173774 65612
rect 255314 65600 255320 65612
rect 173768 65572 255320 65600
rect 173768 65560 173774 65572
rect 255314 65560 255320 65572
rect 255372 65560 255378 65612
rect 297910 65560 297916 65612
rect 297968 65600 297974 65612
rect 433334 65600 433340 65612
rect 297968 65572 433340 65600
rect 297968 65560 297974 65572
rect 433334 65560 433340 65572
rect 433392 65560 433398 65612
rect 206922 65492 206928 65544
rect 206980 65532 206986 65544
rect 303614 65532 303620 65544
rect 206980 65504 303620 65532
rect 206980 65492 206986 65504
rect 303614 65492 303620 65504
rect 303672 65492 303678 65544
rect 391842 65492 391848 65544
rect 391900 65532 391906 65544
rect 569957 65535 570015 65541
rect 569957 65532 569969 65535
rect 391900 65504 569969 65532
rect 391900 65492 391906 65504
rect 569957 65501 569969 65504
rect 570003 65501 570015 65535
rect 569957 65495 570015 65501
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 79594 64852 79600 64864
rect 3384 64824 79600 64852
rect 3384 64812 3390 64824
rect 79594 64812 79600 64824
rect 79652 64812 79658 64864
rect 205450 64200 205456 64252
rect 205508 64240 205514 64252
rect 299474 64240 299480 64252
rect 205508 64212 299480 64240
rect 205508 64200 205514 64212
rect 299474 64200 299480 64212
rect 299532 64200 299538 64252
rect 302142 64200 302148 64252
rect 302200 64240 302206 64252
rect 440234 64240 440240 64252
rect 302200 64212 440240 64240
rect 302200 64200 302206 64212
rect 440234 64200 440240 64212
rect 440292 64200 440298 64252
rect 115842 64132 115848 64184
rect 115900 64172 115906 64184
rect 171134 64172 171140 64184
rect 115900 64144 171140 64172
rect 115900 64132 115906 64144
rect 171134 64132 171140 64144
rect 171192 64132 171198 64184
rect 172422 64132 172428 64184
rect 172480 64172 172486 64184
rect 252554 64172 252560 64184
rect 172480 64144 252560 64172
rect 172480 64132 172486 64144
rect 252554 64132 252560 64144
rect 252612 64132 252618 64184
rect 253842 64132 253848 64184
rect 253900 64172 253906 64184
rect 371234 64172 371240 64184
rect 253900 64144 371240 64172
rect 253900 64132 253906 64144
rect 371234 64132 371240 64144
rect 371292 64132 371298 64184
rect 398098 64132 398104 64184
rect 398156 64172 398162 64184
rect 576854 64172 576860 64184
rect 398156 64144 576860 64172
rect 398156 64132 398162 64144
rect 576854 64132 576860 64144
rect 576912 64132 576918 64184
rect 214926 63452 214932 63504
rect 214984 63492 214990 63504
rect 215018 63492 215024 63504
rect 214984 63464 215024 63492
rect 214984 63452 214990 63464
rect 215018 63452 215024 63464
rect 215076 63452 215082 63504
rect 239858 62948 239864 62960
rect 239819 62920 239864 62948
rect 239858 62908 239864 62920
rect 239916 62908 239922 62960
rect 202782 62840 202788 62892
rect 202840 62880 202846 62892
rect 296714 62880 296720 62892
rect 202840 62852 296720 62880
rect 202840 62840 202846 62852
rect 296714 62840 296720 62852
rect 296772 62840 296778 62892
rect 313918 62840 313924 62892
rect 313976 62880 313982 62892
rect 447134 62880 447140 62892
rect 313976 62852 447140 62880
rect 313976 62840 313982 62852
rect 447134 62840 447140 62852
rect 447192 62840 447198 62892
rect 113082 62772 113088 62824
rect 113140 62812 113146 62824
rect 166994 62812 167000 62824
rect 113140 62784 167000 62812
rect 113140 62772 113146 62784
rect 166994 62772 167000 62784
rect 167052 62772 167058 62824
rect 169662 62772 169668 62824
rect 169720 62812 169726 62824
rect 248414 62812 248420 62824
rect 169720 62784 248420 62812
rect 169720 62772 169726 62784
rect 248414 62772 248420 62784
rect 248472 62772 248478 62824
rect 250438 62772 250444 62824
rect 250496 62812 250502 62824
rect 353294 62812 353300 62824
rect 250496 62784 353300 62812
rect 250496 62772 250502 62784
rect 353294 62772 353300 62784
rect 353352 62772 353358 62824
rect 400122 62772 400128 62824
rect 400180 62812 400186 62824
rect 578878 62812 578884 62824
rect 400180 62784 578884 62812
rect 400180 62772 400186 62784
rect 578878 62772 578884 62784
rect 578936 62772 578942 62824
rect 267090 62744 267096 62756
rect 267051 62716 267096 62744
rect 267090 62704 267096 62716
rect 267148 62704 267154 62756
rect 166902 61412 166908 61464
rect 166960 61452 166966 61464
rect 244274 61452 244280 61464
rect 166960 61424 244280 61452
rect 166960 61412 166966 61424
rect 244274 61412 244280 61424
rect 244332 61412 244338 61464
rect 310422 61412 310428 61464
rect 310480 61452 310486 61464
rect 451274 61452 451280 61464
rect 310480 61424 451280 61452
rect 310480 61412 310486 61424
rect 451274 61412 451280 61424
rect 451332 61412 451338 61464
rect 110322 61344 110328 61396
rect 110380 61384 110386 61396
rect 164234 61384 164240 61396
rect 110380 61356 164240 61384
rect 110380 61344 110386 61356
rect 164234 61344 164240 61356
rect 164292 61344 164298 61396
rect 200022 61344 200028 61396
rect 200080 61384 200086 61396
rect 292574 61384 292580 61396
rect 200080 61356 292580 61384
rect 200080 61344 200086 61356
rect 292574 61344 292580 61356
rect 292632 61344 292638 61396
rect 322842 61344 322848 61396
rect 322900 61384 322906 61396
rect 469214 61384 469220 61396
rect 322900 61356 469220 61384
rect 322900 61344 322906 61356
rect 469214 61344 469220 61356
rect 469272 61344 469278 61396
rect 104618 60840 104624 60852
rect 104544 60812 104624 60840
rect 104544 60716 104572 60812
rect 104618 60800 104624 60812
rect 104676 60800 104682 60852
rect 104526 60664 104532 60716
rect 104584 60664 104590 60716
rect 235902 60052 235908 60104
rect 235960 60092 235966 60104
rect 345014 60092 345020 60104
rect 235960 60064 345020 60092
rect 235960 60052 235966 60064
rect 345014 60052 345020 60064
rect 345072 60052 345078 60104
rect 355318 60052 355324 60104
rect 355376 60092 355382 60104
rect 488534 60092 488540 60104
rect 355376 60064 488540 60092
rect 355376 60052 355382 60064
rect 488534 60052 488540 60064
rect 488592 60052 488598 60104
rect 162670 59984 162676 60036
rect 162728 60024 162734 60036
rect 237374 60024 237380 60036
rect 162728 59996 237380 60024
rect 162728 59984 162734 59996
rect 237374 59984 237380 59996
rect 237432 59984 237438 60036
rect 317230 59984 317236 60036
rect 317288 60024 317294 60036
rect 460934 60024 460940 60036
rect 317288 59996 460940 60024
rect 317288 59984 317294 59996
rect 460934 59984 460940 59996
rect 460992 59984 460998 60036
rect 234430 58760 234436 58812
rect 234488 58800 234494 58812
rect 340874 58800 340880 58812
rect 234488 58772 340880 58800
rect 234488 58760 234494 58772
rect 340874 58760 340880 58772
rect 340932 58760 340938 58812
rect 319990 58692 319996 58744
rect 320048 58732 320054 58744
rect 465074 58732 465080 58744
rect 320048 58704 465080 58732
rect 320048 58692 320054 58704
rect 465074 58692 465080 58704
rect 465132 58692 465138 58744
rect 107562 58624 107568 58676
rect 107620 58664 107626 58676
rect 158714 58664 158720 58676
rect 107620 58636 158720 58664
rect 107620 58624 107626 58636
rect 158714 58624 158720 58636
rect 158772 58624 158778 58676
rect 159910 58624 159916 58676
rect 159968 58664 159974 58676
rect 234614 58664 234620 58676
rect 159968 58636 234620 58664
rect 159968 58624 159974 58636
rect 234614 58624 234620 58636
rect 234672 58624 234678 58676
rect 340690 58624 340696 58676
rect 340748 58664 340754 58676
rect 495434 58664 495440 58676
rect 340748 58636 495440 58664
rect 340748 58624 340754 58636
rect 495434 58624 495440 58636
rect 495492 58624 495498 58676
rect 197722 57944 197728 57996
rect 197780 57984 197786 57996
rect 197998 57984 198004 57996
rect 197780 57956 198004 57984
rect 197780 57944 197786 57956
rect 197998 57944 198004 57956
rect 198056 57944 198062 57996
rect 239674 57944 239680 57996
rect 239732 57984 239738 57996
rect 239861 57987 239919 57993
rect 239861 57984 239873 57987
rect 239732 57956 239873 57984
rect 239732 57944 239738 57956
rect 239861 57953 239873 57956
rect 239907 57953 239919 57987
rect 267090 57984 267096 57996
rect 267051 57956 267096 57984
rect 239861 57947 239919 57953
rect 267090 57944 267096 57956
rect 267148 57944 267154 57996
rect 92109 57919 92167 57925
rect 92109 57885 92121 57919
rect 92155 57916 92167 57919
rect 92198 57916 92204 57928
rect 92155 57888 92204 57916
rect 92155 57885 92167 57888
rect 92109 57879 92167 57885
rect 92198 57876 92204 57888
rect 92256 57876 92262 57928
rect 286870 57332 286876 57384
rect 286928 57372 286934 57384
rect 416866 57372 416872 57384
rect 286928 57344 416872 57372
rect 286928 57332 286934 57344
rect 416866 57332 416872 57344
rect 416924 57332 416930 57384
rect 193030 57264 193036 57316
rect 193088 57304 193094 57316
rect 281534 57304 281540 57316
rect 193088 57276 281540 57304
rect 193088 57264 193094 57276
rect 281534 57264 281540 57276
rect 281592 57264 281598 57316
rect 299382 57264 299388 57316
rect 299440 57304 299446 57316
rect 436094 57304 436100 57316
rect 299440 57276 436100 57304
rect 299440 57264 299446 57276
rect 436094 57264 436100 57276
rect 436152 57264 436158 57316
rect 104526 57196 104532 57248
rect 104584 57236 104590 57248
rect 155954 57236 155960 57248
rect 104584 57208 155960 57236
rect 104584 57196 104590 57208
rect 155954 57196 155960 57208
rect 156012 57196 156018 57248
rect 157242 57196 157248 57248
rect 157300 57236 157306 57248
rect 230474 57236 230480 57248
rect 157300 57208 230480 57236
rect 157300 57196 157306 57208
rect 230474 57196 230480 57208
rect 230532 57196 230538 57248
rect 231118 57196 231124 57248
rect 231176 57236 231182 57248
rect 324314 57236 324320 57248
rect 231176 57208 324320 57236
rect 231176 57196 231182 57208
rect 324314 57196 324320 57208
rect 324372 57196 324378 57248
rect 394602 57196 394608 57248
rect 394660 57236 394666 57248
rect 572714 57236 572720 57248
rect 394660 57208 572720 57236
rect 394660 57196 394666 57208
rect 572714 57196 572720 57208
rect 572772 57196 572778 57248
rect 96246 56624 96252 56636
rect 96207 56596 96252 56624
rect 96246 56584 96252 56596
rect 96304 56584 96310 56636
rect 200114 56624 200120 56636
rect 200075 56596 200120 56624
rect 200114 56584 200120 56596
rect 200172 56584 200178 56636
rect 341889 56627 341947 56633
rect 341889 56593 341901 56627
rect 341935 56624 341947 56627
rect 342070 56624 342076 56636
rect 341935 56596 342076 56624
rect 341935 56593 341947 56596
rect 341889 56587 341947 56593
rect 342070 56584 342076 56596
rect 342128 56584 342134 56636
rect 518894 56624 518900 56636
rect 518855 56596 518900 56624
rect 518894 56584 518900 56596
rect 518952 56584 518958 56636
rect 532694 56624 532700 56636
rect 532655 56596 532700 56624
rect 532694 56584 532700 56596
rect 532752 56584 532758 56636
rect 569954 56624 569960 56636
rect 569915 56596 569960 56624
rect 569954 56584 569960 56596
rect 570012 56584 570018 56636
rect 96246 56488 96252 56500
rect 96207 56460 96252 56488
rect 96246 56448 96252 56460
rect 96304 56448 96310 56500
rect 286962 55972 286968 56024
rect 287020 56012 287026 56024
rect 418154 56012 418160 56024
rect 287020 55984 418160 56012
rect 287020 55972 287026 55984
rect 418154 55972 418160 55984
rect 418212 55972 418218 56024
rect 191098 55904 191104 55956
rect 191156 55944 191162 55956
rect 278774 55944 278780 55956
rect 191156 55916 278780 55944
rect 191156 55904 191162 55916
rect 278774 55904 278780 55916
rect 278832 55904 278838 55956
rect 296622 55904 296628 55956
rect 296680 55944 296686 55956
rect 431954 55944 431960 55956
rect 296680 55916 431960 55944
rect 296680 55904 296686 55916
rect 431954 55904 431960 55916
rect 432012 55904 432018 55956
rect 103330 55836 103336 55888
rect 103388 55876 103394 55888
rect 151814 55876 151820 55888
rect 103388 55848 151820 55876
rect 103388 55836 103394 55848
rect 151814 55836 151820 55848
rect 151872 55836 151878 55888
rect 154390 55836 154396 55888
rect 154448 55876 154454 55888
rect 227806 55876 227812 55888
rect 154448 55848 227812 55876
rect 154448 55836 154454 55848
rect 227806 55836 227812 55848
rect 227864 55836 227870 55888
rect 230290 55836 230296 55888
rect 230348 55876 230354 55888
rect 335354 55876 335360 55888
rect 230348 55848 335360 55876
rect 230348 55836 230354 55848
rect 335354 55836 335360 55848
rect 335412 55836 335418 55888
rect 403618 55836 403624 55888
rect 403676 55876 403682 55888
rect 552014 55876 552020 55888
rect 403676 55848 552020 55876
rect 403676 55836 403682 55848
rect 552014 55836 552020 55848
rect 552072 55836 552078 55888
rect 274358 54612 274364 54664
rect 274416 54652 274422 54664
rect 400214 54652 400220 54664
rect 274416 54624 400220 54652
rect 274416 54612 274422 54624
rect 400214 54612 400220 54624
rect 400272 54612 400278 54664
rect 151446 54544 151452 54596
rect 151504 54584 151510 54596
rect 223574 54584 223580 54596
rect 151504 54556 223580 54584
rect 151504 54544 151510 54556
rect 223574 54544 223580 54556
rect 223632 54544 223638 54596
rect 281442 54544 281448 54596
rect 281500 54584 281506 54596
rect 409874 54584 409880 54596
rect 281500 54556 409880 54584
rect 281500 54544 281506 54556
rect 409874 54544 409880 54556
rect 409932 54544 409938 54596
rect 194502 54476 194508 54528
rect 194560 54516 194566 54528
rect 285674 54516 285680 54528
rect 194560 54488 285680 54516
rect 194560 54476 194566 54488
rect 285674 54476 285680 54488
rect 285732 54476 285738 54528
rect 369762 54476 369768 54528
rect 369820 54516 369826 54528
rect 536926 54516 536932 54528
rect 369820 54488 536932 54516
rect 369820 54476 369826 54488
rect 536926 54476 536932 54488
rect 536984 54476 536990 54528
rect 182082 53116 182088 53168
rect 182140 53156 182146 53168
rect 267737 53159 267795 53165
rect 267737 53156 267749 53159
rect 182140 53128 267749 53156
rect 182140 53116 182146 53128
rect 267737 53125 267749 53128
rect 267783 53125 267795 53159
rect 267737 53119 267795 53125
rect 273162 53116 273168 53168
rect 273220 53156 273226 53168
rect 397454 53156 397460 53168
rect 273220 53128 397460 53156
rect 273220 53116 273226 53128
rect 397454 53116 397460 53128
rect 397512 53116 397518 53168
rect 100570 53048 100576 53100
rect 100628 53088 100634 53100
rect 149054 53088 149060 53100
rect 100628 53060 149060 53088
rect 100628 53048 100634 53060
rect 149054 53048 149060 53060
rect 149112 53048 149118 53100
rect 150342 53048 150348 53100
rect 150400 53088 150406 53100
rect 219434 53088 219440 53100
rect 150400 53060 219440 53088
rect 150400 53048 150406 53060
rect 219434 53048 219440 53060
rect 219492 53048 219498 53100
rect 249610 53048 249616 53100
rect 249668 53088 249674 53100
rect 364334 53088 364340 53100
rect 249668 53060 364340 53088
rect 249668 53048 249674 53060
rect 364334 53048 364340 53060
rect 364392 53048 364398 53100
rect 367002 53048 367008 53100
rect 367060 53088 367066 53100
rect 534074 53088 534080 53100
rect 367060 53060 534080 53088
rect 367060 53048 367066 53060
rect 534074 53048 534080 53060
rect 534132 53048 534138 53100
rect 180702 51756 180708 51808
rect 180760 51796 180766 51808
rect 263594 51796 263600 51808
rect 180760 51768 263600 51796
rect 180760 51756 180766 51768
rect 263594 51756 263600 51768
rect 263652 51756 263658 51808
rect 270310 51756 270316 51808
rect 270368 51796 270374 51808
rect 393314 51796 393320 51808
rect 270368 51768 393320 51796
rect 270368 51756 270374 51768
rect 393314 51756 393320 51768
rect 393372 51756 393378 51808
rect 97902 51688 97908 51740
rect 97960 51728 97966 51740
rect 144914 51728 144920 51740
rect 97960 51700 144920 51728
rect 97960 51688 97966 51700
rect 144914 51688 144920 51700
rect 144972 51688 144978 51740
rect 147582 51688 147588 51740
rect 147640 51728 147646 51740
rect 216674 51728 216680 51740
rect 147640 51700 216680 51728
rect 147640 51688 147646 51700
rect 216674 51688 216680 51700
rect 216732 51688 216738 51740
rect 246942 51688 246948 51740
rect 247000 51728 247006 51740
rect 360194 51728 360200 51740
rect 247000 51700 360200 51728
rect 247000 51688 247006 51700
rect 360194 51688 360200 51700
rect 360252 51688 360258 51740
rect 367738 51688 367744 51740
rect 367796 51728 367802 51740
rect 529934 51728 529940 51740
rect 367796 51700 529940 51728
rect 367796 51688 367802 51700
rect 529934 51688 529940 51700
rect 529992 51688 529998 51740
rect 239674 51116 239680 51128
rect 239635 51088 239680 51116
rect 239674 51076 239680 51088
rect 239732 51076 239738 51128
rect 267090 51116 267096 51128
rect 267051 51088 267096 51116
rect 267090 51076 267096 51088
rect 267148 51076 267154 51128
rect 342070 51076 342076 51128
rect 342128 51076 342134 51128
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 79502 51048 79508 51060
rect 3476 51020 79508 51048
rect 3476 51008 3482 51020
rect 79502 51008 79508 51020
rect 79560 51008 79566 51060
rect 342088 50992 342116 51076
rect 342070 50940 342076 50992
rect 342128 50940 342134 50992
rect 144822 50396 144828 50448
rect 144880 50436 144886 50448
rect 212534 50436 212540 50448
rect 144880 50408 212540 50436
rect 144880 50396 144886 50408
rect 212534 50396 212540 50408
rect 212592 50396 212598 50448
rect 231762 50396 231768 50448
rect 231820 50436 231826 50448
rect 339494 50436 339500 50448
rect 231820 50408 339500 50436
rect 231820 50396 231826 50408
rect 339494 50396 339500 50408
rect 339552 50396 339558 50448
rect 362770 50396 362776 50448
rect 362828 50436 362834 50448
rect 527174 50436 527180 50448
rect 362828 50408 527180 50436
rect 362828 50396 362834 50408
rect 527174 50396 527180 50408
rect 527232 50396 527238 50448
rect 177850 50328 177856 50380
rect 177908 50368 177914 50380
rect 260834 50368 260840 50380
rect 177908 50340 260840 50368
rect 177908 50328 177914 50340
rect 260834 50328 260840 50340
rect 260892 50328 260898 50380
rect 267642 50328 267648 50380
rect 267700 50368 267706 50380
rect 390554 50368 390560 50380
rect 267700 50340 390560 50368
rect 267700 50328 267706 50340
rect 390554 50328 390560 50340
rect 390612 50328 390618 50380
rect 397362 50328 397368 50380
rect 397420 50368 397426 50380
rect 567930 50368 567936 50380
rect 397420 50340 567936 50368
rect 397420 50328 397426 50340
rect 567930 50328 567936 50340
rect 567988 50328 567994 50380
rect 197262 49036 197268 49088
rect 197320 49076 197326 49088
rect 288434 49076 288440 49088
rect 197320 49048 288440 49076
rect 197320 49036 197326 49048
rect 288434 49036 288440 49048
rect 288492 49036 288498 49088
rect 353110 49036 353116 49088
rect 353168 49076 353174 49088
rect 511994 49076 512000 49088
rect 353168 49048 512000 49076
rect 353168 49036 353174 49048
rect 511994 49036 512000 49048
rect 512052 49036 512058 49088
rect 95142 48968 95148 49020
rect 95200 49008 95206 49020
rect 140774 49008 140780 49020
rect 95200 48980 140780 49008
rect 95200 48968 95206 48980
rect 140774 48968 140780 48980
rect 140832 48968 140838 49020
rect 141970 48968 141976 49020
rect 142028 49008 142034 49020
rect 209866 49008 209872 49020
rect 142028 48980 209872 49008
rect 142028 48968 142034 48980
rect 209866 48968 209872 48980
rect 209924 48968 209930 49020
rect 252370 48968 252376 49020
rect 252428 49008 252434 49020
rect 368474 49008 368480 49020
rect 252428 48980 368480 49008
rect 252428 48968 252434 48980
rect 368474 48968 368480 48980
rect 368532 48968 368538 49020
rect 378042 48968 378048 49020
rect 378100 49008 378106 49020
rect 549254 49008 549260 49020
rect 378100 48980 549260 49008
rect 378100 48968 378106 48980
rect 549254 48968 549260 48980
rect 549312 48968 549318 49020
rect 92106 48328 92112 48340
rect 92067 48300 92112 48328
rect 92106 48288 92112 48300
rect 92164 48288 92170 48340
rect 239674 48328 239680 48340
rect 239635 48300 239680 48328
rect 239674 48288 239680 48300
rect 239732 48288 239738 48340
rect 267090 48328 267096 48340
rect 267051 48300 267096 48328
rect 267090 48288 267096 48300
rect 267148 48288 267154 48340
rect 567841 48263 567899 48269
rect 567841 48229 567853 48263
rect 567887 48260 567899 48263
rect 567930 48260 567936 48272
rect 567887 48232 567936 48260
rect 567887 48229 567899 48232
rect 567841 48223 567899 48229
rect 567930 48220 567936 48232
rect 567988 48220 567994 48272
rect 170950 47608 170956 47660
rect 171008 47648 171014 47660
rect 249794 47648 249800 47660
rect 171008 47620 249800 47648
rect 171008 47608 171014 47620
rect 249794 47608 249800 47620
rect 249852 47608 249858 47660
rect 350350 47608 350356 47660
rect 350408 47648 350414 47660
rect 509234 47648 509240 47660
rect 350408 47620 509240 47648
rect 350408 47608 350414 47620
rect 509234 47608 509240 47620
rect 509292 47608 509298 47660
rect 92106 47540 92112 47592
rect 92164 47580 92170 47592
rect 138014 47580 138020 47592
rect 92164 47552 138020 47580
rect 92164 47540 92170 47552
rect 138014 47540 138020 47552
rect 138072 47540 138078 47592
rect 139210 47540 139216 47592
rect 139268 47580 139274 47592
rect 205634 47580 205640 47592
rect 139268 47552 205640 47580
rect 139268 47540 139274 47552
rect 205634 47540 205640 47552
rect 205692 47540 205698 47592
rect 249702 47540 249708 47592
rect 249760 47580 249766 47592
rect 365714 47580 365720 47592
rect 249760 47552 365720 47580
rect 249760 47540 249766 47552
rect 365714 47540 365720 47552
rect 365772 47540 365778 47592
rect 373810 47540 373816 47592
rect 373868 47580 373874 47592
rect 542354 47580 542360 47592
rect 373868 47552 542360 47580
rect 373868 47540 373874 47552
rect 542354 47540 542360 47552
rect 542412 47540 542418 47592
rect 96249 46971 96307 46977
rect 96249 46937 96261 46971
rect 96295 46968 96307 46971
rect 96338 46968 96344 46980
rect 96295 46940 96344 46968
rect 96295 46937 96307 46940
rect 96249 46931 96307 46937
rect 96338 46928 96344 46940
rect 96396 46928 96402 46980
rect 267734 46968 267740 46980
rect 267695 46940 267740 46968
rect 267734 46928 267740 46940
rect 267792 46928 267798 46980
rect 138014 46900 138020 46912
rect 137975 46872 138020 46900
rect 138014 46860 138020 46872
rect 138072 46860 138078 46912
rect 200114 46900 200120 46912
rect 200075 46872 200120 46900
rect 200114 46860 200120 46872
rect 200172 46860 200178 46912
rect 509234 46900 509240 46912
rect 509195 46872 509240 46900
rect 509234 46860 509240 46872
rect 509292 46860 509298 46912
rect 518894 46900 518900 46912
rect 518855 46872 518900 46900
rect 518894 46860 518900 46872
rect 518952 46860 518958 46912
rect 527174 46900 527180 46912
rect 527135 46872 527180 46900
rect 527174 46860 527180 46872
rect 527232 46860 527238 46912
rect 532694 46900 532700 46912
rect 532655 46872 532700 46900
rect 532694 46860 532700 46872
rect 532752 46860 532758 46912
rect 569954 46900 569960 46912
rect 569915 46872 569960 46900
rect 569954 46860 569960 46872
rect 570012 46860 570018 46912
rect 137922 46248 137928 46300
rect 137980 46288 137986 46300
rect 201494 46288 201500 46300
rect 137980 46260 201500 46288
rect 137980 46248 137986 46260
rect 201494 46248 201500 46260
rect 201552 46248 201558 46300
rect 347682 46248 347688 46300
rect 347740 46288 347746 46300
rect 505094 46288 505100 46300
rect 347740 46260 505100 46288
rect 347740 46248 347746 46260
rect 505094 46248 505100 46260
rect 505152 46248 505158 46300
rect 169018 46180 169024 46232
rect 169076 46220 169082 46232
rect 242894 46220 242900 46232
rect 169076 46192 242900 46220
rect 169076 46180 169082 46192
rect 242894 46180 242900 46192
rect 242952 46180 242958 46232
rect 245562 46180 245568 46232
rect 245620 46220 245626 46232
rect 357434 46220 357440 46232
rect 245620 46192 357440 46220
rect 245620 46180 245626 46192
rect 357434 46180 357440 46192
rect 357492 46180 357498 46232
rect 371142 46180 371148 46232
rect 371200 46220 371206 46232
rect 538214 46220 538220 46232
rect 371200 46192 538220 46220
rect 371200 46180 371206 46192
rect 538214 46180 538220 46192
rect 538272 46180 538278 46232
rect 114370 44888 114376 44940
rect 114428 44928 114434 44940
rect 168374 44928 168380 44940
rect 114428 44900 168380 44928
rect 114428 44888 114434 44900
rect 168374 44888 168380 44900
rect 168432 44888 168438 44940
rect 344922 44888 344928 44940
rect 344980 44928 344986 44940
rect 502334 44928 502340 44940
rect 344980 44900 502340 44928
rect 344980 44888 344986 44900
rect 502334 44888 502340 44900
rect 502392 44888 502398 44940
rect 164878 44820 164884 44872
rect 164936 44860 164942 44872
rect 241514 44860 241520 44872
rect 164936 44832 241520 44860
rect 164936 44820 164942 44832
rect 241514 44820 241520 44832
rect 241572 44820 241578 44872
rect 242802 44820 242808 44872
rect 242860 44860 242866 44872
rect 354674 44860 354680 44872
rect 242860 44832 354680 44860
rect 242860 44820 242866 44832
rect 354674 44820 354680 44832
rect 354732 44820 354738 44872
rect 368382 44820 368388 44872
rect 368440 44860 368446 44872
rect 535454 44860 535460 44872
rect 368440 44832 535460 44860
rect 368440 44820 368446 44832
rect 535454 44820 535460 44832
rect 535512 44820 535518 44872
rect 168190 43460 168196 43512
rect 168248 43500 168254 43512
rect 245654 43500 245660 43512
rect 168248 43472 245660 43500
rect 168248 43460 168254 43472
rect 245654 43460 245660 43472
rect 245712 43460 245718 43512
rect 342070 43460 342076 43512
rect 342128 43500 342134 43512
rect 498194 43500 498200 43512
rect 342128 43472 498200 43500
rect 342128 43460 342134 43472
rect 498194 43460 498200 43472
rect 498252 43460 498258 43512
rect 135162 43392 135168 43444
rect 135220 43432 135226 43444
rect 198734 43432 198740 43444
rect 135220 43404 198740 43432
rect 135220 43392 135226 43404
rect 198734 43392 198740 43404
rect 198792 43392 198798 43444
rect 239674 43392 239680 43444
rect 239732 43432 239738 43444
rect 350534 43432 350540 43444
rect 239732 43404 350540 43432
rect 239732 43392 239738 43404
rect 350534 43392 350540 43404
rect 350592 43392 350598 43444
rect 365622 43392 365628 43444
rect 365680 43432 365686 43444
rect 531314 43432 531320 43444
rect 365680 43404 531320 43432
rect 365680 43392 365686 43404
rect 531314 43392 531320 43404
rect 531372 43392 531378 43444
rect 132402 42100 132408 42152
rect 132460 42140 132466 42152
rect 194594 42140 194600 42152
rect 132460 42112 194600 42140
rect 132460 42100 132466 42112
rect 194594 42100 194600 42112
rect 194652 42100 194658 42152
rect 340782 42100 340788 42152
rect 340840 42140 340846 42152
rect 494054 42140 494060 42152
rect 340840 42112 494060 42140
rect 340840 42100 340846 42112
rect 494054 42100 494060 42112
rect 494112 42100 494118 42152
rect 160002 42032 160008 42084
rect 160060 42072 160066 42084
rect 235994 42072 236000 42084
rect 160060 42044 236000 42072
rect 160060 42032 160066 42044
rect 235994 42032 236000 42044
rect 236052 42032 236058 42084
rect 238662 42032 238668 42084
rect 238720 42072 238726 42084
rect 347774 42072 347780 42084
rect 238720 42044 347780 42072
rect 238720 42032 238726 42044
rect 347774 42032 347780 42044
rect 347832 42032 347838 42084
rect 355962 42032 355968 42084
rect 356020 42072 356026 42084
rect 517514 42072 517520 42084
rect 356020 42044 517520 42072
rect 356020 42032 356026 42044
rect 517514 42032 517520 42044
rect 517572 42032 517578 42084
rect 267001 41531 267059 41537
rect 267001 41497 267013 41531
rect 267047 41528 267059 41531
rect 267090 41528 267096 41540
rect 267047 41500 267096 41528
rect 267047 41497 267059 41500
rect 267001 41491 267059 41497
rect 267090 41488 267096 41500
rect 267148 41488 267154 41540
rect 96338 41460 96344 41472
rect 96264 41432 96344 41460
rect 96264 41404 96292 41432
rect 96338 41420 96344 41432
rect 96396 41420 96402 41472
rect 214926 41420 214932 41472
rect 214984 41420 214990 41472
rect 227254 41420 227260 41472
rect 227312 41420 227318 41472
rect 96246 41352 96252 41404
rect 96304 41352 96310 41404
rect 214944 41324 214972 41420
rect 215018 41324 215024 41336
rect 214944 41296 215024 41324
rect 215018 41284 215024 41296
rect 215076 41284 215082 41336
rect 227272 41324 227300 41420
rect 402330 41352 402336 41404
rect 402388 41392 402394 41404
rect 580166 41392 580172 41404
rect 402388 41364 580172 41392
rect 402388 41352 402394 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 227346 41324 227352 41336
rect 227272 41296 227352 41324
rect 227346 41284 227352 41296
rect 227404 41284 227410 41336
rect 226242 40808 226248 40860
rect 226300 40848 226306 40860
rect 329834 40848 329840 40860
rect 226300 40820 329840 40848
rect 226300 40808 226306 40820
rect 329834 40808 329840 40820
rect 329892 40808 329898 40860
rect 270402 40740 270408 40792
rect 270460 40780 270466 40792
rect 394694 40780 394700 40792
rect 270460 40752 394700 40780
rect 270460 40740 270466 40752
rect 394694 40740 394700 40752
rect 394752 40740 394758 40792
rect 129550 40672 129556 40724
rect 129608 40712 129614 40724
rect 191834 40712 191840 40724
rect 129608 40684 191840 40712
rect 129608 40672 129614 40684
rect 191834 40672 191840 40684
rect 191892 40672 191898 40724
rect 284202 40672 284208 40724
rect 284260 40712 284266 40724
rect 414014 40712 414020 40724
rect 284260 40684 414020 40712
rect 284260 40672 284266 40684
rect 414014 40672 414020 40684
rect 414072 40672 414078 40724
rect 184842 39380 184848 39432
rect 184900 39420 184906 39432
rect 270586 39420 270592 39432
rect 184900 39392 270592 39420
rect 184900 39380 184906 39392
rect 270586 39380 270592 39392
rect 270644 39380 270650 39432
rect 326982 39380 326988 39432
rect 327040 39420 327046 39432
rect 476114 39420 476120 39432
rect 327040 39392 476120 39420
rect 327040 39380 327046 39392
rect 476114 39380 476120 39392
rect 476172 39380 476178 39432
rect 126790 39312 126796 39364
rect 126848 39352 126854 39364
rect 187694 39352 187700 39364
rect 126848 39324 187700 39352
rect 126848 39312 126854 39324
rect 187694 39312 187700 39324
rect 187752 39312 187758 39364
rect 223390 39312 223396 39364
rect 223448 39352 223454 39364
rect 325694 39352 325700 39364
rect 223448 39324 325700 39352
rect 223448 39312 223454 39324
rect 325694 39312 325700 39324
rect 325752 39312 325758 39364
rect 346302 39312 346308 39364
rect 346360 39352 346366 39364
rect 502426 39352 502432 39364
rect 346360 39324 502432 39352
rect 346360 39312 346366 39324
rect 502426 39312 502432 39324
rect 502484 39312 502490 39364
rect 266998 38672 267004 38684
rect 266959 38644 267004 38672
rect 266998 38632 267004 38644
rect 267056 38632 267062 38684
rect 567838 38672 567844 38684
rect 567799 38644 567844 38672
rect 567838 38632 567844 38644
rect 567896 38632 567902 38684
rect 198550 38564 198556 38616
rect 198608 38604 198614 38616
rect 198734 38604 198740 38616
rect 198608 38576 198740 38604
rect 198608 38564 198614 38576
rect 198734 38564 198740 38576
rect 198792 38564 198798 38616
rect 162762 38020 162768 38072
rect 162820 38060 162826 38072
rect 238754 38060 238760 38072
rect 162820 38032 238760 38060
rect 162820 38020 162826 38032
rect 238754 38020 238760 38032
rect 238812 38020 238818 38072
rect 220722 37952 220728 38004
rect 220780 37992 220786 38004
rect 321646 37992 321652 38004
rect 220780 37964 321652 37992
rect 220780 37952 220786 37964
rect 321646 37952 321652 37964
rect 321704 37952 321710 38004
rect 331858 37952 331864 38004
rect 331916 37992 331922 38004
rect 478874 37992 478880 38004
rect 331916 37964 478880 37992
rect 331916 37952 331922 37964
rect 478874 37952 478880 37964
rect 478932 37952 478938 38004
rect 122742 37884 122748 37936
rect 122800 37924 122806 37936
rect 180794 37924 180800 37936
rect 122800 37896 180800 37924
rect 122800 37884 122806 37896
rect 180794 37884 180800 37896
rect 180852 37884 180858 37936
rect 237282 37884 237288 37936
rect 237340 37924 237346 37936
rect 346394 37924 346400 37936
rect 237340 37896 346400 37924
rect 237340 37884 237346 37896
rect 346394 37884 346400 37896
rect 346452 37884 346458 37936
rect 348970 37884 348976 37936
rect 349028 37924 349034 37936
rect 506474 37924 506480 37936
rect 349028 37896 506480 37924
rect 349028 37884 349034 37896
rect 506474 37884 506480 37896
rect 506532 37884 506538 37936
rect 138014 37312 138020 37324
rect 137975 37284 138020 37312
rect 138014 37272 138020 37284
rect 138072 37272 138078 37324
rect 200114 37312 200120 37324
rect 200075 37284 200120 37312
rect 200114 37272 200120 37284
rect 200172 37272 200178 37324
rect 509234 37312 509240 37324
rect 509195 37284 509240 37312
rect 509234 37272 509240 37284
rect 509292 37272 509298 37324
rect 518894 37312 518900 37324
rect 518855 37284 518900 37312
rect 518894 37272 518900 37284
rect 518952 37272 518958 37324
rect 527174 37312 527180 37324
rect 527135 37284 527180 37312
rect 527174 37272 527180 37284
rect 527232 37272 527238 37324
rect 532694 37312 532700 37324
rect 532655 37284 532700 37312
rect 532694 37272 532700 37284
rect 532752 37272 532758 37324
rect 569954 37312 569960 37324
rect 569915 37284 569960 37312
rect 569954 37272 569960 37284
rect 570012 37272 570018 37324
rect 215018 37244 215024 37256
rect 214979 37216 215024 37244
rect 215018 37204 215024 37216
rect 215076 37204 215082 37256
rect 227346 37244 227352 37256
rect 227307 37216 227352 37244
rect 227346 37204 227352 37216
rect 227404 37204 227410 37256
rect 314562 36592 314568 36644
rect 314620 36632 314626 36644
rect 458174 36632 458180 36644
rect 314620 36604 458180 36632
rect 314620 36592 314626 36604
rect 458174 36592 458180 36604
rect 458232 36592 458238 36644
rect 119982 36524 119988 36576
rect 120040 36564 120046 36576
rect 176654 36564 176660 36576
rect 120040 36536 176660 36564
rect 120040 36524 120046 36536
rect 176654 36524 176660 36536
rect 176712 36524 176718 36576
rect 213822 36524 213828 36576
rect 213880 36564 213886 36576
rect 311894 36564 311900 36576
rect 213880 36536 311900 36564
rect 213880 36524 213886 36536
rect 311894 36524 311900 36536
rect 311952 36524 311958 36576
rect 328270 36524 328276 36576
rect 328328 36564 328334 36576
rect 477586 36564 477592 36576
rect 328328 36536 477592 36564
rect 328328 36524 328334 36536
rect 477586 36524 477592 36536
rect 477644 36524 477650 36576
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 21358 35884 21364 35896
rect 3476 35856 21364 35884
rect 3476 35844 3482 35856
rect 21358 35844 21364 35856
rect 21416 35844 21422 35896
rect 190362 35232 190368 35284
rect 190420 35272 190426 35284
rect 278866 35272 278872 35284
rect 190420 35244 278872 35272
rect 190420 35232 190426 35244
rect 278866 35232 278872 35244
rect 278924 35232 278930 35284
rect 280062 35232 280068 35284
rect 280120 35272 280126 35284
rect 408586 35272 408592 35284
rect 280120 35244 408592 35272
rect 280120 35232 280126 35244
rect 408586 35232 408592 35244
rect 408644 35232 408650 35284
rect 117130 35164 117136 35216
rect 117188 35204 117194 35216
rect 173894 35204 173900 35216
rect 117188 35176 173900 35204
rect 117188 35164 117194 35176
rect 173894 35164 173900 35176
rect 173952 35164 173958 35216
rect 252462 35164 252468 35216
rect 252520 35204 252526 35216
rect 367094 35204 367100 35216
rect 252520 35176 367100 35204
rect 252520 35164 252526 35176
rect 367094 35164 367100 35176
rect 367152 35164 367158 35216
rect 372522 35164 372528 35216
rect 372580 35204 372586 35216
rect 540974 35204 540980 35216
rect 372580 35176 540980 35204
rect 372580 35164 372586 35176
rect 540974 35164 540980 35176
rect 541032 35164 541038 35216
rect 360102 33804 360108 33856
rect 360160 33844 360166 33856
rect 523034 33844 523040 33856
rect 360160 33816 523040 33844
rect 360160 33804 360166 33816
rect 523034 33804 523040 33816
rect 523092 33804 523098 33856
rect 114462 33736 114468 33788
rect 114520 33776 114526 33788
rect 169754 33776 169760 33788
rect 114520 33748 169760 33776
rect 114520 33736 114526 33748
rect 169754 33736 169760 33748
rect 169812 33736 169818 33788
rect 177942 33736 177948 33788
rect 178000 33776 178006 33788
rect 262306 33776 262312 33788
rect 178000 33748 262312 33776
rect 178000 33736 178006 33748
rect 262306 33736 262312 33748
rect 262364 33736 262370 33788
rect 264882 33736 264888 33788
rect 264940 33776 264946 33788
rect 386414 33776 386420 33788
rect 264940 33748 386420 33776
rect 264940 33736 264946 33748
rect 386414 33736 386420 33748
rect 386472 33736 386478 33788
rect 387702 33736 387708 33788
rect 387760 33776 387766 33788
rect 563146 33776 563152 33788
rect 387760 33748 563152 33776
rect 387760 33736 387766 33748
rect 563146 33736 563152 33748
rect 563204 33736 563210 33788
rect 357342 32444 357348 32496
rect 357400 32484 357406 32496
rect 520274 32484 520280 32496
rect 357400 32456 520280 32484
rect 357400 32444 357406 32456
rect 520274 32444 520280 32456
rect 520332 32444 520338 32496
rect 115198 32376 115204 32428
rect 115256 32416 115262 32428
rect 167086 32416 167092 32428
rect 115256 32388 167092 32416
rect 115256 32376 115262 32388
rect 167086 32376 167092 32388
rect 167144 32376 167150 32428
rect 176562 32376 176568 32428
rect 176620 32416 176626 32428
rect 258074 32416 258080 32428
rect 176620 32388 258080 32416
rect 176620 32376 176626 32388
rect 258074 32376 258080 32388
rect 258132 32376 258138 32428
rect 260742 32376 260748 32428
rect 260800 32416 260806 32428
rect 379514 32416 379520 32428
rect 260800 32388 379520 32416
rect 260800 32376 260806 32388
rect 379514 32376 379520 32388
rect 379572 32376 379578 32428
rect 384942 32376 384948 32428
rect 385000 32416 385006 32428
rect 560294 32416 560300 32428
rect 385000 32388 560300 32416
rect 385000 32376 385006 32388
rect 560294 32376 560300 32388
rect 560352 32376 560358 32428
rect 96246 31804 96252 31816
rect 96172 31776 96252 31804
rect 96172 31748 96200 31776
rect 96246 31764 96252 31776
rect 96304 31764 96310 31816
rect 96154 31696 96160 31748
rect 96212 31696 96218 31748
rect 197998 31696 198004 31748
rect 198056 31736 198062 31748
rect 198182 31736 198188 31748
rect 198056 31708 198188 31736
rect 198056 31696 198062 31708
rect 198182 31696 198188 31708
rect 198240 31696 198246 31748
rect 266998 31696 267004 31748
rect 267056 31736 267062 31748
rect 267182 31736 267188 31748
rect 267056 31708 267188 31736
rect 267056 31696 267062 31708
rect 267182 31696 267188 31708
rect 267240 31696 267246 31748
rect 567838 31696 567844 31748
rect 567896 31736 567902 31748
rect 568022 31736 568028 31748
rect 567896 31708 568028 31736
rect 567896 31696 567902 31708
rect 568022 31696 568028 31708
rect 568080 31696 568086 31748
rect 354582 31084 354588 31136
rect 354640 31124 354646 31136
rect 516134 31124 516140 31136
rect 354640 31096 516140 31124
rect 354640 31084 354646 31096
rect 516134 31084 516140 31096
rect 516192 31084 516198 31136
rect 111058 31016 111064 31068
rect 111116 31056 111122 31068
rect 162854 31056 162860 31068
rect 111116 31028 162860 31056
rect 111116 31016 111122 31028
rect 162854 31016 162860 31028
rect 162912 31016 162918 31068
rect 173802 31016 173808 31068
rect 173860 31056 173866 31068
rect 253934 31056 253940 31068
rect 173860 31028 253940 31056
rect 173860 31016 173866 31028
rect 253934 31016 253940 31028
rect 253992 31016 253998 31068
rect 255222 31016 255228 31068
rect 255280 31056 255286 31068
rect 372614 31056 372620 31068
rect 255280 31028 372620 31056
rect 255280 31016 255286 31028
rect 372614 31016 372620 31028
rect 372672 31016 372678 31068
rect 380710 31016 380716 31068
rect 380768 31056 380774 31068
rect 553394 31056 553400 31068
rect 380768 31028 553400 31056
rect 380768 31016 380774 31028
rect 553394 31016 553400 31028
rect 553452 31016 553458 31068
rect 402238 30268 402244 30320
rect 402296 30308 402302 30320
rect 580166 30308 580172 30320
rect 402296 30280 580172 30308
rect 402296 30268 402302 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 248230 29656 248236 29708
rect 248288 29696 248294 29708
rect 361574 29696 361580 29708
rect 248288 29668 361580 29696
rect 248288 29656 248294 29668
rect 361574 29656 361580 29668
rect 361632 29656 361638 29708
rect 106090 29588 106096 29640
rect 106148 29628 106154 29640
rect 158806 29628 158812 29640
rect 106148 29600 158812 29628
rect 106148 29588 106154 29600
rect 158806 29588 158812 29600
rect 158864 29588 158870 29640
rect 168282 29588 168288 29640
rect 168340 29628 168346 29640
rect 247034 29628 247040 29640
rect 168340 29600 247040 29628
rect 168340 29588 168346 29600
rect 247034 29588 247040 29600
rect 247092 29588 247098 29640
rect 288342 29588 288348 29640
rect 288400 29628 288406 29640
rect 419534 29628 419540 29640
rect 288400 29600 419540 29628
rect 288400 29588 288406 29600
rect 419534 29588 419540 29600
rect 419592 29588 419598 29640
rect 198093 28951 198151 28957
rect 198093 28917 198105 28951
rect 198139 28948 198151 28951
rect 198182 28948 198188 28960
rect 198139 28920 198188 28948
rect 198139 28917 198151 28920
rect 198093 28911 198151 28917
rect 198182 28908 198188 28920
rect 198240 28908 198246 28960
rect 267093 28951 267151 28957
rect 267093 28917 267105 28951
rect 267139 28948 267151 28951
rect 267182 28948 267188 28960
rect 267139 28920 267188 28948
rect 267139 28917 267151 28920
rect 267093 28911 267151 28917
rect 267182 28908 267188 28920
rect 267240 28908 267246 28960
rect 337930 28296 337936 28348
rect 337988 28336 337994 28348
rect 491294 28336 491300 28348
rect 337988 28308 491300 28336
rect 337988 28296 337994 28308
rect 491294 28296 491300 28308
rect 491352 28296 491358 28348
rect 90910 28228 90916 28280
rect 90968 28268 90974 28280
rect 133874 28268 133880 28280
rect 90968 28240 133880 28268
rect 90968 28228 90974 28240
rect 133874 28228 133880 28240
rect 133932 28228 133938 28280
rect 158622 28228 158628 28280
rect 158680 28268 158686 28280
rect 233234 28268 233240 28280
rect 158680 28240 233240 28268
rect 158680 28228 158686 28240
rect 233234 28228 233240 28240
rect 233292 28228 233298 28280
rect 236638 28228 236644 28280
rect 236696 28268 236702 28280
rect 343634 28268 343640 28280
rect 236696 28240 343640 28268
rect 236696 28228 236702 28240
rect 343634 28228 343640 28240
rect 343692 28228 343698 28280
rect 361482 28228 361488 28280
rect 361540 28268 361546 28280
rect 524506 28268 524512 28280
rect 361540 28240 524512 28268
rect 361540 28228 361546 28240
rect 524506 28228 524512 28240
rect 524564 28228 524570 28280
rect 215021 27659 215079 27665
rect 215021 27625 215033 27659
rect 215067 27656 215079 27659
rect 215110 27656 215116 27668
rect 215067 27628 215116 27656
rect 215067 27625 215079 27628
rect 215021 27619 215079 27625
rect 215110 27616 215116 27628
rect 215168 27616 215174 27668
rect 227349 27659 227407 27665
rect 227349 27625 227361 27659
rect 227395 27656 227407 27659
rect 227438 27656 227444 27668
rect 227395 27628 227444 27656
rect 227395 27625 227407 27628
rect 227349 27619 227407 27625
rect 227438 27616 227444 27628
rect 227496 27616 227502 27668
rect 138014 27548 138020 27600
rect 138072 27588 138078 27600
rect 138474 27588 138480 27600
rect 138072 27560 138480 27588
rect 138072 27548 138078 27560
rect 138474 27548 138480 27560
rect 138532 27548 138538 27600
rect 198734 27548 198740 27600
rect 198792 27548 198798 27600
rect 509234 27588 509240 27600
rect 509195 27560 509240 27588
rect 509234 27548 509240 27560
rect 509292 27548 509298 27600
rect 518894 27588 518900 27600
rect 518855 27560 518900 27588
rect 518894 27548 518900 27560
rect 518952 27548 518958 27600
rect 527174 27588 527180 27600
rect 527135 27560 527180 27588
rect 527174 27548 527180 27560
rect 527232 27548 527238 27600
rect 532694 27588 532700 27600
rect 532655 27560 532700 27588
rect 532694 27548 532700 27560
rect 532752 27548 532758 27600
rect 568022 27588 568028 27600
rect 567983 27560 568028 27588
rect 568022 27548 568028 27560
rect 568080 27548 568086 27600
rect 569954 27588 569960 27600
rect 569915 27560 569960 27588
rect 569954 27548 569960 27560
rect 570012 27548 570018 27600
rect 198752 27461 198780 27548
rect 198737 27455 198795 27461
rect 198737 27421 198749 27455
rect 198783 27421 198795 27455
rect 198737 27415 198795 27421
rect 335262 26936 335268 26988
rect 335320 26976 335326 26988
rect 487154 26976 487160 26988
rect 335320 26948 487160 26976
rect 335320 26936 335326 26948
rect 487154 26936 487160 26948
rect 487212 26936 487218 26988
rect 104802 26868 104808 26920
rect 104860 26908 104866 26920
rect 154574 26908 154580 26920
rect 104860 26880 154580 26908
rect 104860 26868 104866 26880
rect 154574 26868 154580 26880
rect 154632 26868 154638 26920
rect 155862 26868 155868 26920
rect 155920 26908 155926 26920
rect 229094 26908 229100 26920
rect 155920 26880 229100 26908
rect 155920 26868 155926 26880
rect 229094 26868 229100 26880
rect 229152 26868 229158 26920
rect 230382 26868 230388 26920
rect 230440 26908 230446 26920
rect 336734 26908 336740 26920
rect 230440 26880 336740 26908
rect 230440 26868 230446 26880
rect 336734 26868 336740 26880
rect 336792 26868 336798 26920
rect 353202 26868 353208 26920
rect 353260 26908 353266 26920
rect 513374 26908 513380 26920
rect 353260 26880 513380 26908
rect 353260 26868 353266 26880
rect 513374 26868 513380 26880
rect 513432 26868 513438 26920
rect 332502 25576 332508 25628
rect 332560 25616 332566 25628
rect 484394 25616 484400 25628
rect 332560 25588 484400 25616
rect 332560 25576 332566 25588
rect 484394 25576 484400 25588
rect 484452 25576 484458 25628
rect 102042 25508 102048 25560
rect 102100 25548 102106 25560
rect 150526 25548 150532 25560
rect 102100 25520 150532 25548
rect 102100 25508 102106 25520
rect 150526 25508 150532 25520
rect 150584 25508 150590 25560
rect 154482 25508 154488 25560
rect 154540 25548 154546 25560
rect 226334 25548 226340 25560
rect 154540 25520 226340 25548
rect 154540 25508 154546 25520
rect 226334 25508 226340 25520
rect 226392 25508 226398 25560
rect 227438 25508 227444 25560
rect 227496 25548 227502 25560
rect 332594 25548 332600 25560
rect 227496 25520 332600 25548
rect 227496 25508 227502 25520
rect 332594 25508 332600 25520
rect 332652 25508 332658 25560
rect 350442 25508 350448 25560
rect 350500 25548 350506 25560
rect 510706 25548 510712 25560
rect 350500 25520 510712 25548
rect 350500 25508 350506 25520
rect 510706 25508 510712 25520
rect 510764 25508 510770 25560
rect 224218 24148 224224 24200
rect 224276 24188 224282 24200
rect 318794 24188 318800 24200
rect 224276 24160 318800 24188
rect 224276 24148 224282 24160
rect 318794 24148 318800 24160
rect 318852 24148 318858 24200
rect 324130 24148 324136 24200
rect 324188 24188 324194 24200
rect 471974 24188 471980 24200
rect 324188 24160 471980 24188
rect 324188 24148 324194 24160
rect 471974 24148 471980 24160
rect 472032 24148 472038 24200
rect 99190 24080 99196 24132
rect 99248 24120 99254 24132
rect 147674 24120 147680 24132
rect 99248 24092 147680 24120
rect 99248 24080 99254 24092
rect 147674 24080 147680 24092
rect 147732 24080 147738 24132
rect 151722 24080 151728 24132
rect 151780 24120 151786 24132
rect 222194 24120 222200 24132
rect 151780 24092 222200 24120
rect 151780 24080 151786 24092
rect 222194 24080 222200 24092
rect 222252 24080 222258 24132
rect 234522 24080 234528 24132
rect 234580 24120 234586 24132
rect 342254 24120 342260 24132
rect 234580 24092 342260 24120
rect 234580 24080 234586 24092
rect 342254 24080 342260 24092
rect 342312 24080 342318 24132
rect 343542 24080 343548 24132
rect 343600 24120 343606 24132
rect 499574 24120 499580 24132
rect 343600 24092 499580 24120
rect 343600 24080 343606 24092
rect 499574 24080 499580 24092
rect 499632 24080 499638 24132
rect 200114 22828 200120 22840
rect 200075 22800 200120 22828
rect 200114 22788 200120 22800
rect 200172 22788 200178 22840
rect 215110 22788 215116 22840
rect 215168 22828 215174 22840
rect 314654 22828 314660 22840
rect 215168 22800 314660 22828
rect 215168 22788 215174 22800
rect 314654 22788 314660 22800
rect 314712 22788 314718 22840
rect 321370 22788 321376 22840
rect 321428 22828 321434 22840
rect 467926 22828 467932 22840
rect 321428 22800 467932 22828
rect 321428 22788 321434 22800
rect 467926 22788 467932 22800
rect 467984 22788 467990 22840
rect 96154 22720 96160 22772
rect 96212 22760 96218 22772
rect 143534 22760 143540 22772
rect 96212 22732 143540 22760
rect 96212 22720 96218 22732
rect 143534 22720 143540 22732
rect 143592 22720 143598 22772
rect 148962 22720 148968 22772
rect 149020 22760 149026 22772
rect 218146 22760 218152 22772
rect 149020 22732 218152 22760
rect 149020 22720 149026 22732
rect 218146 22720 218152 22732
rect 218204 22720 218210 22772
rect 227622 22720 227628 22772
rect 227680 22760 227686 22772
rect 331306 22760 331312 22772
rect 227680 22732 331312 22760
rect 227680 22720 227686 22732
rect 331306 22720 331312 22732
rect 331364 22720 331370 22772
rect 338022 22720 338028 22772
rect 338080 22760 338086 22772
rect 492674 22760 492680 22772
rect 338080 22732 492680 22760
rect 338080 22720 338086 22732
rect 492674 22720 492680 22732
rect 492732 22720 492738 22772
rect 267734 22692 267740 22704
rect 267695 22664 267740 22692
rect 267734 22652 267740 22664
rect 267792 22652 267798 22704
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 79410 22080 79416 22092
rect 3200 22052 79416 22080
rect 3200 22040 3206 22052
rect 79410 22040 79416 22052
rect 79468 22040 79474 22092
rect 208302 21428 208308 21480
rect 208360 21468 208366 21480
rect 305086 21468 305092 21480
rect 208360 21440 305092 21468
rect 208360 21428 208366 21440
rect 305086 21428 305092 21440
rect 305144 21428 305150 21480
rect 318058 21428 318064 21480
rect 318116 21468 318122 21480
rect 454034 21468 454040 21480
rect 318116 21440 454040 21468
rect 318116 21428 318122 21440
rect 454034 21428 454040 21440
rect 454092 21428 454098 21480
rect 88978 21360 88984 21412
rect 89036 21400 89042 21412
rect 131114 21400 131120 21412
rect 89036 21372 131120 21400
rect 89036 21360 89042 21372
rect 131114 21360 131120 21372
rect 131172 21360 131178 21412
rect 143442 21360 143448 21412
rect 143500 21400 143506 21412
rect 211154 21400 211160 21412
rect 143500 21372 211160 21400
rect 143500 21360 143506 21372
rect 211154 21360 211160 21372
rect 211212 21360 211218 21412
rect 217962 21360 217968 21412
rect 218020 21400 218026 21412
rect 317414 21400 317420 21412
rect 218020 21372 317420 21400
rect 218020 21360 218026 21372
rect 317414 21360 317420 21372
rect 317472 21360 317478 21412
rect 326338 21360 326344 21412
rect 326396 21400 326402 21412
rect 473354 21400 473360 21412
rect 326396 21372 473360 21400
rect 326396 21360 326402 21372
rect 473354 21360 473360 21372
rect 473412 21360 473418 21412
rect 142062 20000 142068 20052
rect 142120 20040 142126 20052
rect 208394 20040 208400 20052
rect 142120 20012 208400 20040
rect 142120 20000 142126 20012
rect 208394 20000 208400 20012
rect 208452 20000 208458 20052
rect 304902 20000 304908 20052
rect 304960 20040 304966 20052
rect 443086 20040 443092 20052
rect 304960 20012 443092 20040
rect 304960 20000 304966 20012
rect 443086 20000 443092 20012
rect 443144 20000 443150 20052
rect 446398 20000 446404 20052
rect 446456 20040 446462 20052
rect 571426 20040 571432 20052
rect 446456 20012 571432 20040
rect 446456 20000 446462 20012
rect 571426 20000 571432 20012
rect 571484 20000 571490 20052
rect 97258 19932 97264 19984
rect 97316 19972 97322 19984
rect 140866 19972 140872 19984
rect 97316 19944 140872 19972
rect 97316 19932 97322 19944
rect 140866 19932 140872 19944
rect 140924 19932 140930 19984
rect 205542 19932 205548 19984
rect 205600 19972 205606 19984
rect 300854 19972 300860 19984
rect 205600 19944 300860 19972
rect 205600 19932 205606 19944
rect 300854 19932 300860 19944
rect 300912 19932 300918 19984
rect 320082 19932 320088 19984
rect 320140 19972 320146 19984
rect 466454 19972 466460 19984
rect 320140 19944 466460 19972
rect 320140 19932 320146 19944
rect 466454 19932 466460 19944
rect 466512 19932 466518 19984
rect 198090 19360 198096 19372
rect 198051 19332 198096 19360
rect 198090 19320 198096 19332
rect 198148 19320 198154 19372
rect 267090 19360 267096 19372
rect 267051 19332 267096 19360
rect 267090 19320 267096 19332
rect 267148 19320 267154 19372
rect 491294 19292 491300 19304
rect 491255 19264 491300 19292
rect 491294 19252 491300 19264
rect 491352 19252 491358 19304
rect 492674 19252 492680 19304
rect 492732 19292 492738 19304
rect 510614 19292 510620 19304
rect 492732 19264 492777 19292
rect 510575 19264 510620 19292
rect 492732 19252 492738 19264
rect 510614 19252 510620 19264
rect 510672 19252 510678 19304
rect 516134 19292 516140 19304
rect 516095 19264 516140 19292
rect 516134 19252 516140 19264
rect 516192 19252 516198 19304
rect 547874 19252 547880 19304
rect 547932 19292 547938 19304
rect 548886 19292 548892 19304
rect 547932 19264 548892 19292
rect 547932 19252 547938 19264
rect 548886 19252 548892 19264
rect 548944 19252 548950 19304
rect 550634 19252 550640 19304
rect 550692 19292 550698 19304
rect 553394 19292 553400 19304
rect 550692 19264 550737 19292
rect 553355 19264 553400 19292
rect 550692 19252 550698 19264
rect 553394 19252 553400 19264
rect 553452 19252 553458 19304
rect 560294 19252 560300 19304
rect 560352 19292 560358 19304
rect 560754 19292 560760 19304
rect 560352 19264 560760 19292
rect 560352 19252 560358 19264
rect 560754 19252 560760 19264
rect 560812 19252 560818 19304
rect 283558 18708 283564 18760
rect 283616 18748 283622 18760
rect 400306 18748 400312 18760
rect 283616 18720 400312 18748
rect 283616 18708 283622 18720
rect 400306 18708 400312 18720
rect 400364 18708 400370 18760
rect 269022 18640 269028 18692
rect 269080 18680 269086 18692
rect 390646 18680 390652 18692
rect 269080 18652 390652 18680
rect 269080 18640 269086 18652
rect 390646 18640 390652 18652
rect 390704 18640 390710 18692
rect 92382 18572 92388 18624
rect 92440 18612 92446 18624
rect 136634 18612 136640 18624
rect 92440 18584 136640 18612
rect 92440 18572 92446 18584
rect 136634 18572 136640 18584
rect 136692 18572 136698 18624
rect 139302 18572 139308 18624
rect 139360 18612 139366 18624
rect 204254 18612 204260 18624
rect 139360 18584 204260 18612
rect 139360 18572 139366 18584
rect 204254 18572 204260 18584
rect 204312 18572 204318 18624
rect 207658 18572 207664 18624
rect 207716 18612 207722 18624
rect 296806 18612 296812 18624
rect 207716 18584 296812 18612
rect 207716 18572 207722 18584
rect 296806 18572 296812 18584
rect 296864 18572 296870 18624
rect 380802 18572 380808 18624
rect 380860 18612 380866 18624
rect 554866 18612 554872 18624
rect 380860 18584 554872 18612
rect 380860 18572 380866 18584
rect 554866 18572 554872 18584
rect 554924 18572 554930 18624
rect 518894 18000 518900 18012
rect 518855 17972 518900 18000
rect 518894 17960 518900 17972
rect 518952 17960 518958 18012
rect 527174 18000 527180 18012
rect 527135 17972 527180 18000
rect 527174 17960 527180 17972
rect 527232 17960 527238 18012
rect 568022 18000 568028 18012
rect 567983 17972 568028 18000
rect 568022 17960 568028 17972
rect 568080 17960 568086 18012
rect 555418 17892 555424 17944
rect 555476 17932 555482 17944
rect 579798 17932 579804 17944
rect 555476 17904 579804 17932
rect 555476 17892 555482 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 257982 17348 257988 17400
rect 258040 17388 258046 17400
rect 376754 17388 376760 17400
rect 258040 17360 376760 17388
rect 258040 17348 258046 17360
rect 376754 17348 376760 17360
rect 376812 17348 376818 17400
rect 136542 17280 136548 17332
rect 136600 17320 136606 17332
rect 201586 17320 201592 17332
rect 136600 17292 201592 17320
rect 136600 17280 136606 17292
rect 201586 17280 201592 17292
rect 201644 17280 201650 17332
rect 272518 17280 272524 17332
rect 272576 17320 272582 17332
rect 396074 17320 396080 17332
rect 272576 17292 396080 17320
rect 272576 17280 272582 17292
rect 396074 17280 396080 17292
rect 396132 17280 396138 17332
rect 89622 17212 89628 17264
rect 89680 17252 89686 17264
rect 132586 17252 132592 17264
rect 89680 17224 132592 17252
rect 89680 17212 89686 17224
rect 132586 17212 132592 17224
rect 132644 17212 132650 17264
rect 201402 17212 201408 17264
rect 201460 17252 201466 17264
rect 293954 17252 293960 17264
rect 201460 17224 293960 17252
rect 201460 17212 201466 17224
rect 293954 17212 293960 17224
rect 294012 17212 294018 17264
rect 376662 17212 376668 17264
rect 376720 17252 376726 17264
rect 546494 17252 546500 17264
rect 376720 17224 546500 17252
rect 376720 17212 376726 17224
rect 546494 17212 546500 17224
rect 546552 17212 546558 17264
rect 344278 15988 344284 16040
rect 344336 16028 344342 16040
rect 451366 16028 451372 16040
rect 344336 16000 451372 16028
rect 344336 15988 344342 16000
rect 451366 15988 451372 16000
rect 451424 15988 451430 16040
rect 195882 15920 195888 15972
rect 195940 15960 195946 15972
rect 287146 15960 287152 15972
rect 195940 15932 287152 15960
rect 195940 15920 195946 15932
rect 287146 15920 287152 15932
rect 287204 15920 287210 15972
rect 291102 15920 291108 15972
rect 291160 15960 291166 15972
rect 425146 15960 425152 15972
rect 291160 15932 425152 15960
rect 291160 15920 291166 15932
rect 425146 15920 425152 15932
rect 425204 15920 425210 15972
rect 86862 15852 86868 15904
rect 86920 15892 86926 15904
rect 129734 15892 129740 15904
rect 86920 15864 129740 15892
rect 86920 15852 86926 15864
rect 129734 15852 129740 15864
rect 129792 15852 129798 15904
rect 131758 15852 131764 15904
rect 131816 15892 131822 15904
rect 193306 15892 193312 15904
rect 131816 15864 193312 15892
rect 131816 15852 131822 15864
rect 193306 15852 193312 15864
rect 193364 15852 193370 15904
rect 261478 15852 261484 15904
rect 261536 15892 261542 15904
rect 374086 15892 374092 15904
rect 261536 15864 374092 15892
rect 261536 15852 261542 15864
rect 374086 15852 374092 15864
rect 374144 15852 374150 15904
rect 398742 15852 398748 15904
rect 398800 15892 398806 15904
rect 578970 15892 578976 15904
rect 398800 15864 578976 15892
rect 398800 15852 398806 15864
rect 578970 15852 578976 15864
rect 579028 15852 579034 15904
rect 527174 14832 527180 14884
rect 527232 14872 527238 14884
rect 527358 14872 527364 14884
rect 527232 14844 527364 14872
rect 527232 14832 527238 14844
rect 527358 14832 527364 14844
rect 527416 14832 527422 14884
rect 193122 14492 193128 14544
rect 193180 14532 193186 14544
rect 282914 14532 282920 14544
rect 193180 14504 282920 14532
rect 193180 14492 193186 14504
rect 282914 14492 282920 14504
rect 282972 14492 282978 14544
rect 333790 14492 333796 14544
rect 333848 14532 333854 14544
rect 485866 14532 485872 14544
rect 333848 14504 485872 14532
rect 333848 14492 333854 14504
rect 485866 14492 485872 14504
rect 485924 14492 485930 14544
rect 85482 14424 85488 14476
rect 85540 14464 85546 14476
rect 126974 14464 126980 14476
rect 85540 14436 126980 14464
rect 85540 14424 85546 14436
rect 126974 14424 126980 14436
rect 127032 14424 127038 14476
rect 129642 14424 129648 14476
rect 129700 14464 129706 14476
rect 190454 14464 190460 14476
rect 129700 14436 190460 14464
rect 129700 14424 129706 14436
rect 190454 14424 190460 14436
rect 190512 14424 190518 14476
rect 251082 14424 251088 14476
rect 251140 14464 251146 14476
rect 365806 14464 365812 14476
rect 251140 14436 365812 14464
rect 251140 14424 251146 14436
rect 365806 14424 365812 14436
rect 365864 14424 365870 14476
rect 386322 14424 386328 14476
rect 386380 14464 386386 14476
rect 561950 14464 561956 14476
rect 386380 14436 561956 14464
rect 386380 14424 386386 14436
rect 561950 14424 561956 14436
rect 562008 14424 562014 14476
rect 106918 13132 106924 13184
rect 106976 13172 106982 13184
rect 128354 13172 128360 13184
rect 106976 13144 128360 13172
rect 106976 13132 106982 13144
rect 128354 13132 128360 13144
rect 128412 13132 128418 13184
rect 188982 13132 188988 13184
rect 189040 13172 189046 13184
rect 276014 13172 276020 13184
rect 189040 13144 276020 13172
rect 189040 13132 189046 13144
rect 276014 13132 276020 13144
rect 276072 13132 276078 13184
rect 294598 13132 294604 13184
rect 294656 13172 294662 13184
rect 382274 13172 382280 13184
rect 294656 13144 382280 13172
rect 294656 13132 294662 13144
rect 382274 13132 382280 13144
rect 382332 13132 382338 13184
rect 126882 13064 126888 13116
rect 126940 13104 126946 13116
rect 186314 13104 186320 13116
rect 126940 13076 186320 13104
rect 126940 13064 126946 13076
rect 186314 13064 186320 13076
rect 186372 13064 186378 13116
rect 248322 13064 248328 13116
rect 248380 13104 248386 13116
rect 362954 13104 362960 13116
rect 248380 13076 362960 13104
rect 248380 13064 248386 13076
rect 362954 13064 362960 13076
rect 363012 13064 363018 13116
rect 373902 13064 373908 13116
rect 373960 13104 373966 13116
rect 544102 13104 544108 13116
rect 373960 13076 544108 13104
rect 373960 13064 373966 13076
rect 544102 13064 544108 13076
rect 544160 13064 544166 13116
rect 517514 12452 517520 12504
rect 517572 12452 517578 12504
rect 518894 12452 518900 12504
rect 518952 12452 518958 12504
rect 524414 12452 524420 12504
rect 524472 12452 524478 12504
rect 545114 12452 545120 12504
rect 545172 12452 545178 12504
rect 568574 12452 568580 12504
rect 568632 12452 568638 12504
rect 133874 12384 133880 12436
rect 133932 12424 133938 12436
rect 134794 12424 134800 12436
rect 133932 12396 134800 12424
rect 133932 12384 133938 12396
rect 134794 12384 134800 12396
rect 134852 12384 134858 12436
rect 136634 12384 136640 12436
rect 136692 12424 136698 12436
rect 137186 12424 137192 12436
rect 136692 12396 137192 12424
rect 136692 12384 136698 12396
rect 137186 12384 137192 12396
rect 137244 12384 137250 12436
rect 143534 12384 143540 12436
rect 143592 12424 143598 12436
rect 144454 12424 144460 12436
rect 143592 12396 144460 12424
rect 143592 12384 143598 12396
rect 144454 12384 144460 12396
rect 144512 12384 144518 12436
rect 144914 12384 144920 12436
rect 144972 12424 144978 12436
rect 145650 12424 145656 12436
rect 144972 12396 145656 12424
rect 144972 12384 144978 12396
rect 145650 12384 145656 12396
rect 145708 12384 145714 12436
rect 195974 12384 195980 12436
rect 196032 12424 196038 12436
rect 196802 12424 196808 12436
rect 196032 12396 196808 12424
rect 196032 12384 196038 12396
rect 196802 12384 196808 12396
rect 196860 12384 196866 12436
rect 202874 12384 202880 12436
rect 202932 12424 202938 12436
rect 203886 12424 203892 12436
rect 202932 12396 203892 12424
rect 202932 12384 202938 12396
rect 203886 12384 203892 12396
rect 203944 12384 203950 12436
rect 204254 12384 204260 12436
rect 204312 12424 204318 12436
rect 205082 12424 205088 12436
rect 204312 12396 205088 12424
rect 204312 12384 204318 12396
rect 205082 12384 205088 12396
rect 205140 12384 205146 12436
rect 263594 12384 263600 12436
rect 263652 12424 263658 12436
rect 264606 12424 264612 12436
rect 263652 12396 264612 12424
rect 263652 12384 263658 12396
rect 264606 12384 264612 12396
rect 264664 12384 264670 12436
rect 266354 12384 266360 12436
rect 266412 12424 266418 12436
rect 266998 12424 267004 12436
rect 266412 12396 267004 12424
rect 266412 12384 266418 12396
rect 266998 12384 267004 12396
rect 267056 12384 267062 12436
rect 270586 12384 270592 12436
rect 270644 12424 270650 12436
rect 271690 12424 271696 12436
rect 270644 12396 271696 12424
rect 270644 12384 270650 12396
rect 271690 12384 271696 12396
rect 271748 12384 271754 12436
rect 487154 12384 487160 12436
rect 487212 12424 487218 12436
rect 488166 12424 488172 12436
rect 487212 12396 488172 12424
rect 487212 12384 487218 12396
rect 488166 12384 488172 12396
rect 488224 12384 488230 12436
rect 488534 12384 488540 12436
rect 488592 12424 488598 12436
rect 489362 12424 489368 12436
rect 488592 12396 489368 12424
rect 488592 12384 488598 12396
rect 489362 12384 489368 12396
rect 489420 12384 489426 12436
rect 505094 12384 505100 12436
rect 505152 12424 505158 12436
rect 506014 12424 506020 12436
rect 505152 12396 506020 12424
rect 505152 12384 505158 12396
rect 506014 12384 506020 12396
rect 506072 12384 506078 12436
rect 506474 12384 506480 12436
rect 506532 12424 506538 12436
rect 507210 12424 507216 12436
rect 506532 12396 507216 12424
rect 506532 12384 506538 12396
rect 507210 12384 507216 12396
rect 507268 12384 507274 12436
rect 513374 12384 513380 12436
rect 513432 12424 513438 12436
rect 514386 12424 514392 12436
rect 513432 12396 514392 12424
rect 513432 12384 513438 12396
rect 514386 12384 514392 12396
rect 514444 12384 514450 12436
rect 514754 12384 514760 12436
rect 514812 12424 514818 12436
rect 515582 12424 515588 12436
rect 514812 12396 515588 12424
rect 514812 12384 514818 12396
rect 515582 12384 515588 12396
rect 515640 12384 515646 12436
rect 517532 12356 517560 12452
rect 517882 12356 517888 12368
rect 517532 12328 517888 12356
rect 517882 12316 517888 12328
rect 517940 12316 517946 12368
rect 518912 12356 518940 12452
rect 521654 12384 521660 12436
rect 521712 12424 521718 12436
rect 522666 12424 522672 12436
rect 521712 12396 522672 12424
rect 521712 12384 521718 12396
rect 522666 12384 522672 12396
rect 522724 12384 522730 12436
rect 523034 12384 523040 12436
rect 523092 12424 523098 12436
rect 523862 12424 523868 12436
rect 523092 12396 523868 12424
rect 523092 12384 523098 12396
rect 523862 12384 523868 12396
rect 523920 12384 523926 12436
rect 519078 12356 519084 12368
rect 518912 12328 519084 12356
rect 519078 12316 519084 12328
rect 519136 12316 519142 12368
rect 524432 12356 524460 12452
rect 529934 12384 529940 12436
rect 529992 12424 529998 12436
rect 531038 12424 531044 12436
rect 529992 12396 531044 12424
rect 529992 12384 529998 12396
rect 531038 12384 531044 12396
rect 531096 12384 531102 12436
rect 531314 12384 531320 12436
rect 531372 12424 531378 12436
rect 532234 12424 532240 12436
rect 531372 12396 532240 12424
rect 531372 12384 531378 12396
rect 532234 12384 532240 12396
rect 532292 12384 532298 12436
rect 525058 12356 525064 12368
rect 524432 12328 525064 12356
rect 525058 12316 525064 12328
rect 525116 12316 525122 12368
rect 545132 12356 545160 12452
rect 549254 12384 549260 12436
rect 549312 12424 549318 12436
rect 550082 12424 550088 12436
rect 549312 12396 550088 12424
rect 549312 12384 549318 12396
rect 550082 12384 550088 12396
rect 550140 12384 550146 12436
rect 557534 12384 557540 12436
rect 557592 12424 557598 12436
rect 558362 12424 558368 12436
rect 557592 12396 558368 12424
rect 557592 12384 557598 12396
rect 558362 12384 558368 12396
rect 558420 12384 558426 12436
rect 564434 12384 564440 12436
rect 564492 12424 564498 12436
rect 565538 12424 565544 12436
rect 564492 12396 565544 12424
rect 564492 12384 564498 12396
rect 565538 12384 565544 12396
rect 565596 12384 565602 12436
rect 565814 12384 565820 12436
rect 565872 12424 565878 12436
rect 566734 12424 566740 12436
rect 565872 12396 566740 12424
rect 565872 12384 565878 12396
rect 566734 12384 566740 12396
rect 566792 12384 566798 12436
rect 568592 12424 568620 12452
rect 569034 12424 569040 12436
rect 568592 12396 569040 12424
rect 569034 12384 569040 12396
rect 569092 12384 569098 12436
rect 545298 12356 545304 12368
rect 545132 12328 545304 12356
rect 545298 12316 545304 12328
rect 545356 12316 545362 12368
rect 550637 12359 550695 12365
rect 550637 12325 550649 12359
rect 550683 12356 550695 12359
rect 551186 12356 551192 12368
rect 550683 12328 551192 12356
rect 550683 12325 550695 12328
rect 550637 12319 550695 12325
rect 551186 12316 551192 12328
rect 551244 12316 551250 12368
rect 552106 12316 552112 12368
rect 552164 12356 552170 12368
rect 552382 12356 552388 12368
rect 552164 12328 552388 12356
rect 552164 12316 552170 12328
rect 552382 12316 552388 12328
rect 552440 12316 552446 12368
rect 186222 11840 186228 11892
rect 186280 11880 186286 11892
rect 272886 11880 272892 11892
rect 186280 11852 272892 11880
rect 186280 11840 186286 11852
rect 272886 11840 272892 11852
rect 272944 11840 272950 11892
rect 241422 11772 241428 11824
rect 241480 11812 241486 11824
rect 351914 11812 351920 11824
rect 241480 11784 351920 11812
rect 241480 11772 241486 11784
rect 351914 11772 351920 11784
rect 351972 11772 351978 11824
rect 363598 11772 363604 11824
rect 363656 11812 363662 11824
rect 526254 11812 526260 11824
rect 363656 11784 526260 11812
rect 363656 11772 363662 11784
rect 526254 11772 526260 11784
rect 526312 11772 526318 11824
rect 124122 11704 124128 11756
rect 124180 11744 124186 11756
rect 183554 11744 183560 11756
rect 124180 11716 183560 11744
rect 124180 11704 124186 11716
rect 183554 11704 183560 11716
rect 183612 11704 183618 11756
rect 259362 11704 259368 11756
rect 259420 11744 259426 11756
rect 378134 11744 378140 11756
rect 259420 11716 378140 11744
rect 259420 11704 259426 11716
rect 378134 11704 378140 11716
rect 378192 11704 378198 11756
rect 390462 11704 390468 11756
rect 390520 11744 390526 11756
rect 567838 11744 567844 11756
rect 390520 11716 567844 11744
rect 390520 11704 390526 11716
rect 567838 11704 567844 11716
rect 567896 11704 567902 11756
rect 266262 10412 266268 10464
rect 266320 10452 266326 10464
rect 389174 10452 389180 10464
rect 266320 10424 389180 10452
rect 266320 10412 266326 10424
rect 389174 10412 389180 10424
rect 389232 10412 389238 10464
rect 183462 10344 183468 10396
rect 183520 10384 183526 10396
rect 269298 10384 269304 10396
rect 183520 10356 269304 10384
rect 183520 10344 183526 10356
rect 269298 10344 269304 10356
rect 269356 10344 269362 10396
rect 351822 10344 351828 10396
rect 351880 10384 351886 10396
rect 512086 10384 512092 10396
rect 351880 10356 512092 10384
rect 351880 10344 351886 10356
rect 512086 10344 512092 10356
rect 512144 10344 512150 10396
rect 121362 10276 121368 10328
rect 121420 10316 121426 10328
rect 179414 10316 179420 10328
rect 121420 10288 179420 10316
rect 121420 10276 121426 10288
rect 179414 10276 179420 10288
rect 179472 10276 179478 10328
rect 246298 10276 246304 10328
rect 246356 10316 246362 10328
rect 347866 10316 347872 10328
rect 246356 10288 347872 10316
rect 246356 10276 246362 10288
rect 347866 10276 347872 10288
rect 347924 10276 347930 10328
rect 383562 10276 383568 10328
rect 383620 10316 383626 10328
rect 557166 10316 557172 10328
rect 383620 10288 557172 10316
rect 383620 10276 383626 10288
rect 557166 10276 557172 10288
rect 557224 10276 557230 10328
rect 198737 9707 198795 9713
rect 198737 9673 198749 9707
rect 198783 9704 198795 9707
rect 199194 9704 199200 9716
rect 198783 9676 199200 9704
rect 198783 9673 198795 9676
rect 198737 9667 198795 9673
rect 199194 9664 199200 9676
rect 199252 9664 199258 9716
rect 200117 9707 200175 9713
rect 200117 9673 200129 9707
rect 200163 9704 200175 9707
rect 200390 9704 200396 9716
rect 200163 9676 200396 9704
rect 200163 9673 200175 9676
rect 200117 9667 200175 9673
rect 200390 9664 200396 9676
rect 200448 9664 200454 9716
rect 267737 9707 267795 9713
rect 267737 9673 267749 9707
rect 267783 9704 267795 9707
rect 268102 9704 268108 9716
rect 267783 9676 268108 9704
rect 267783 9673 267795 9676
rect 267737 9667 267795 9673
rect 268102 9664 268108 9676
rect 268160 9664 268166 9716
rect 491297 9707 491355 9713
rect 491297 9673 491309 9707
rect 491343 9704 491355 9707
rect 491754 9704 491760 9716
rect 491343 9676 491760 9704
rect 491343 9673 491355 9676
rect 491297 9667 491355 9673
rect 491754 9664 491760 9676
rect 491812 9664 491818 9716
rect 492677 9707 492735 9713
rect 492677 9673 492689 9707
rect 492723 9704 492735 9707
rect 492950 9704 492956 9716
rect 492723 9676 492956 9704
rect 492723 9673 492735 9676
rect 492677 9667 492735 9673
rect 492950 9664 492956 9676
rect 493008 9664 493014 9716
rect 509237 9707 509295 9713
rect 509237 9673 509249 9707
rect 509283 9704 509295 9707
rect 509602 9704 509608 9716
rect 509283 9676 509608 9704
rect 509283 9673 509295 9676
rect 509237 9667 509295 9673
rect 509602 9664 509608 9676
rect 509660 9664 509666 9716
rect 510617 9707 510675 9713
rect 510617 9673 510629 9707
rect 510663 9704 510675 9707
rect 510798 9704 510804 9716
rect 510663 9676 510804 9704
rect 510663 9673 510675 9676
rect 510617 9667 510675 9673
rect 510798 9664 510804 9676
rect 510856 9664 510862 9716
rect 516137 9707 516195 9713
rect 516137 9673 516149 9707
rect 516183 9704 516195 9707
rect 516778 9704 516784 9716
rect 516183 9676 516784 9704
rect 516183 9673 516195 9676
rect 516137 9667 516195 9673
rect 516778 9664 516784 9676
rect 516836 9664 516842 9716
rect 532697 9707 532755 9713
rect 532697 9673 532709 9707
rect 532743 9704 532755 9707
rect 533430 9704 533436 9716
rect 532743 9676 533436 9704
rect 532743 9673 532755 9676
rect 532697 9667 532755 9673
rect 533430 9664 533436 9676
rect 533488 9664 533494 9716
rect 553397 9707 553455 9713
rect 553397 9673 553409 9707
rect 553443 9704 553455 9707
rect 553578 9704 553584 9716
rect 553443 9676 553584 9704
rect 553443 9673 553455 9676
rect 553397 9667 553455 9673
rect 553578 9664 553584 9676
rect 553636 9664 553642 9716
rect 569957 9707 570015 9713
rect 569957 9673 569969 9707
rect 570003 9704 570015 9707
rect 570230 9704 570236 9716
rect 570003 9676 570236 9704
rect 570003 9673 570015 9676
rect 569957 9667 570015 9673
rect 570230 9664 570236 9676
rect 570288 9664 570294 9716
rect 517882 9636 517888 9648
rect 517843 9608 517888 9636
rect 517882 9596 517888 9608
rect 517940 9596 517946 9648
rect 519078 9636 519084 9648
rect 519039 9608 519084 9636
rect 519078 9596 519084 9608
rect 519136 9596 519142 9648
rect 525058 9596 525064 9648
rect 525116 9596 525122 9648
rect 527450 9596 527456 9648
rect 527508 9596 527514 9648
rect 545298 9636 545304 9648
rect 545259 9608 545304 9636
rect 545298 9596 545304 9608
rect 545356 9596 545362 9648
rect 548886 9636 548892 9648
rect 548847 9608 548892 9636
rect 548886 9596 548892 9608
rect 548944 9596 548950 9648
rect 550082 9636 550088 9648
rect 550043 9608 550088 9636
rect 550082 9596 550088 9608
rect 550140 9596 550146 9648
rect 525076 9512 525104 9596
rect 527468 9512 527496 9596
rect 525058 9460 525064 9512
rect 525116 9460 525122 9512
rect 527450 9460 527456 9512
rect 527508 9460 527514 9512
rect 171042 9052 171048 9104
rect 171100 9092 171106 9104
rect 251450 9092 251456 9104
rect 171100 9064 251456 9092
rect 171100 9052 171106 9064
rect 251450 9052 251456 9064
rect 251508 9052 251514 9104
rect 223482 8984 223488 9036
rect 223540 9024 223546 9036
rect 327626 9024 327632 9036
rect 223540 8996 327632 9024
rect 223540 8984 223546 8996
rect 327626 8984 327632 8996
rect 327684 8984 327690 9036
rect 349062 8984 349068 9036
rect 349120 9024 349126 9036
rect 508406 9024 508412 9036
rect 349120 8996 508412 9024
rect 349120 8984 349126 8996
rect 508406 8984 508412 8996
rect 508464 8984 508470 9036
rect 118602 8916 118608 8968
rect 118660 8956 118666 8968
rect 176562 8956 176568 8968
rect 118660 8928 176568 8956
rect 118660 8916 118666 8928
rect 176562 8916 176568 8928
rect 176620 8916 176626 8968
rect 244182 8916 244188 8968
rect 244240 8956 244246 8968
rect 357342 8956 357348 8968
rect 244240 8928 357348 8956
rect 244240 8916 244246 8928
rect 357342 8916 357348 8928
rect 357400 8916 357406 8968
rect 375282 8916 375288 8968
rect 375340 8956 375346 8968
rect 546586 8956 546592 8968
rect 375340 8928 546592 8956
rect 375340 8916 375346 8928
rect 546586 8916 546592 8928
rect 546644 8916 546650 8968
rect 135898 8644 135904 8696
rect 135956 8684 135962 8696
rect 144825 8687 144883 8693
rect 144825 8684 144837 8687
rect 135956 8656 144837 8684
rect 135956 8644 135962 8656
rect 144825 8653 144837 8656
rect 144871 8653 144883 8687
rect 144825 8647 144883 8653
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 79318 8276 79324 8288
rect 3476 8248 79324 8276
rect 3476 8236 3482 8248
rect 79318 8236 79324 8248
rect 79376 8236 79382 8288
rect 174538 7692 174544 7744
rect 174596 7732 174602 7744
rect 244366 7732 244372 7744
rect 174596 7704 244372 7732
rect 174596 7692 174602 7704
rect 244366 7692 244372 7704
rect 244424 7692 244430 7744
rect 494146 7732 494152 7744
rect 489932 7704 494152 7732
rect 132586 7624 132592 7676
rect 132644 7664 132650 7676
rect 133782 7664 133788 7676
rect 132644 7636 133788 7664
rect 132644 7624 132650 7636
rect 133782 7624 133788 7636
rect 133840 7624 133846 7676
rect 140774 7624 140780 7676
rect 140832 7664 140838 7676
rect 142062 7664 142068 7676
rect 140832 7636 142068 7664
rect 140832 7624 140838 7636
rect 142062 7624 142068 7636
rect 142120 7624 142126 7676
rect 222102 7624 222108 7676
rect 222160 7664 222166 7676
rect 324038 7664 324044 7676
rect 222160 7636 324044 7664
rect 222160 7624 222166 7636
rect 324038 7624 324044 7636
rect 324096 7624 324102 7676
rect 339402 7624 339408 7676
rect 339460 7664 339466 7676
rect 489932 7664 489960 7704
rect 494146 7692 494152 7704
rect 494204 7692 494210 7744
rect 339460 7636 489960 7664
rect 339460 7624 339466 7636
rect 494054 7624 494060 7676
rect 494112 7664 494118 7676
rect 495342 7664 495348 7676
rect 494112 7636 495348 7664
rect 494112 7624 494118 7636
rect 495342 7624 495348 7636
rect 495400 7624 495406 7676
rect 511994 7624 512000 7676
rect 512052 7664 512058 7676
rect 513190 7664 513196 7676
rect 512052 7636 513196 7664
rect 512052 7624 512058 7636
rect 513190 7624 513196 7636
rect 513248 7624 513254 7676
rect 117222 7556 117228 7608
rect 117280 7596 117286 7608
rect 172974 7596 172980 7608
rect 117280 7568 172980 7596
rect 117280 7556 117286 7568
rect 172974 7556 172980 7568
rect 173032 7556 173038 7608
rect 201494 7556 201500 7608
rect 201552 7596 201558 7608
rect 202690 7596 202696 7608
rect 201552 7568 202696 7596
rect 201552 7556 201558 7568
rect 202690 7556 202696 7568
rect 202748 7556 202754 7608
rect 240042 7556 240048 7608
rect 240100 7596 240106 7608
rect 350258 7596 350264 7608
rect 240100 7568 350264 7596
rect 240100 7556 240106 7568
rect 350258 7556 350264 7568
rect 350316 7556 350322 7608
rect 362862 7556 362868 7608
rect 362920 7596 362926 7608
rect 362920 7568 525748 7596
rect 362920 7556 362926 7568
rect 485774 7488 485780 7540
rect 485832 7528 485838 7540
rect 486970 7528 486976 7540
rect 485832 7500 486976 7528
rect 485832 7488 485838 7500
rect 486970 7488 486976 7500
rect 487028 7488 487034 7540
rect 525720 7528 525748 7568
rect 528554 7556 528560 7608
rect 528612 7596 528618 7608
rect 529842 7596 529848 7608
rect 528612 7568 529848 7596
rect 528612 7556 528618 7568
rect 529842 7556 529848 7568
rect 529900 7556 529906 7608
rect 546494 7556 546500 7608
rect 546552 7596 546558 7608
rect 547690 7596 547696 7608
rect 546552 7568 547696 7596
rect 546552 7556 546558 7568
rect 547690 7556 547696 7568
rect 547748 7556 547754 7608
rect 554774 7556 554780 7608
rect 554832 7596 554838 7608
rect 555970 7596 555976 7608
rect 554832 7568 555976 7596
rect 554832 7556 554838 7568
rect 555970 7556 555976 7568
rect 556028 7556 556034 7608
rect 563146 7556 563152 7608
rect 563204 7596 563210 7608
rect 564342 7596 564348 7608
rect 563204 7568 564348 7596
rect 563204 7556 563210 7568
rect 564342 7556 564348 7568
rect 564400 7556 564406 7608
rect 571334 7556 571340 7608
rect 571392 7596 571398 7608
rect 572622 7596 572628 7608
rect 571392 7568 572628 7596
rect 571392 7556 571398 7568
rect 572622 7556 572628 7568
rect 572680 7556 572686 7608
rect 528646 7528 528652 7540
rect 525720 7500 528652 7528
rect 528646 7488 528652 7500
rect 528704 7488 528710 7540
rect 482186 7284 482192 7336
rect 482244 7324 482250 7336
rect 486513 7327 486571 7333
rect 486513 7324 486525 7327
rect 482244 7296 486525 7324
rect 482244 7284 482250 7296
rect 486513 7293 486525 7296
rect 486559 7293 486571 7327
rect 486513 7287 486571 7293
rect 161382 6196 161388 6248
rect 161440 6236 161446 6248
rect 237190 6236 237196 6248
rect 161440 6208 237196 6236
rect 161440 6196 161446 6208
rect 237190 6196 237196 6208
rect 237248 6196 237254 6248
rect 336642 6196 336648 6248
rect 336700 6236 336706 6248
rect 490558 6236 490564 6248
rect 336700 6208 490564 6236
rect 336700 6196 336706 6208
rect 490558 6196 490564 6208
rect 490616 6196 490622 6248
rect 111702 6128 111708 6180
rect 111760 6168 111766 6180
rect 165890 6168 165896 6180
rect 111760 6140 165896 6168
rect 111760 6128 111766 6140
rect 165890 6128 165896 6140
rect 165948 6128 165954 6180
rect 233142 6128 233148 6180
rect 233200 6168 233206 6180
rect 340690 6168 340696 6180
rect 233200 6140 340696 6168
rect 233200 6128 233206 6140
rect 340690 6128 340696 6140
rect 340748 6128 340754 6180
rect 358722 6128 358728 6180
rect 358780 6168 358786 6180
rect 521470 6168 521476 6180
rect 358780 6140 521476 6168
rect 358780 6128 358786 6140
rect 521470 6128 521476 6140
rect 521528 6128 521534 6180
rect 84102 4836 84108 4888
rect 84160 4876 84166 4888
rect 126606 4876 126612 4888
rect 84160 4848 126612 4876
rect 84160 4836 84166 4848
rect 126606 4836 126612 4848
rect 126664 4836 126670 4888
rect 144825 4879 144883 4885
rect 144825 4845 144837 4879
rect 144871 4876 144883 4879
rect 154577 4879 154635 4885
rect 154577 4876 154589 4879
rect 144871 4848 154589 4876
rect 144871 4845 144883 4848
rect 144825 4839 144883 4845
rect 154577 4845 154589 4848
rect 154623 4845 154635 4879
rect 154577 4839 154635 4845
rect 178678 4836 178684 4888
rect 178736 4876 178742 4888
rect 197998 4876 198004 4888
rect 178736 4848 198004 4876
rect 178736 4836 178742 4848
rect 197998 4836 198004 4848
rect 198056 4836 198062 4888
rect 198182 4836 198188 4888
rect 198240 4876 198246 4888
rect 253842 4876 253848 4888
rect 198240 4848 253848 4876
rect 198240 4836 198246 4848
rect 253842 4836 253848 4848
rect 253900 4836 253906 4888
rect 291838 4836 291844 4888
rect 291896 4876 291902 4888
rect 383562 4876 383568 4888
rect 291896 4848 383568 4876
rect 291896 4836 291902 4848
rect 383562 4836 383568 4848
rect 383620 4836 383626 4888
rect 420178 4836 420184 4888
rect 420236 4876 420242 4888
rect 483474 4876 483480 4888
rect 420236 4848 483480 4876
rect 420236 4836 420242 4848
rect 483474 4836 483480 4848
rect 483532 4836 483538 4888
rect 125502 4768 125508 4820
rect 125560 4808 125566 4820
rect 144914 4808 144920 4820
rect 125560 4780 144920 4808
rect 125560 4768 125566 4780
rect 144914 4768 144920 4780
rect 144972 4768 144978 4820
rect 145006 4768 145012 4820
rect 145064 4808 145070 4820
rect 184842 4808 184848 4820
rect 145064 4780 184848 4808
rect 145064 4768 145070 4780
rect 184842 4768 184848 4780
rect 184900 4768 184906 4820
rect 203518 4768 203524 4820
rect 203576 4808 203582 4820
rect 265802 4808 265808 4820
rect 203576 4780 265808 4808
rect 203576 4768 203582 4780
rect 265802 4768 265808 4780
rect 265860 4768 265866 4820
rect 267182 4768 267188 4820
rect 267240 4808 267246 4820
rect 290734 4808 290740 4820
rect 267240 4780 290740 4808
rect 267240 4768 267246 4780
rect 290734 4768 290740 4780
rect 290792 4768 290798 4820
rect 298002 4768 298008 4820
rect 298060 4808 298066 4820
rect 434622 4808 434628 4820
rect 298060 4780 434628 4808
rect 298060 4768 298066 4780
rect 434622 4768 434628 4780
rect 434680 4768 434686 4820
rect 493318 4768 493324 4820
rect 493376 4808 493382 4820
rect 559558 4808 559564 4820
rect 493376 4780 559564 4808
rect 493376 4768 493382 4780
rect 559558 4768 559564 4780
rect 559616 4768 559622 4820
rect 347866 4156 347872 4208
rect 347924 4196 347930 4208
rect 349062 4196 349068 4208
rect 347924 4168 349068 4196
rect 347924 4156 347930 4168
rect 349062 4156 349068 4168
rect 349120 4156 349126 4208
rect 400214 4156 400220 4208
rect 400272 4196 400278 4208
rect 401318 4196 401324 4208
rect 400272 4168 401324 4196
rect 400272 4156 400278 4168
rect 401318 4156 401324 4168
rect 401376 4156 401382 4208
rect 408494 4156 408500 4208
rect 408552 4196 408558 4208
rect 409690 4196 409696 4208
rect 408552 4168 409696 4196
rect 408552 4156 408558 4168
rect 409690 4156 409696 4168
rect 409748 4156 409754 4208
rect 306282 4088 306288 4140
rect 306340 4128 306346 4140
rect 446582 4128 446588 4140
rect 306340 4100 446588 4128
rect 306340 4088 306346 4100
rect 446582 4088 446588 4100
rect 446640 4088 446646 4140
rect 309042 4020 309048 4072
rect 309100 4060 309106 4072
rect 450170 4060 450176 4072
rect 309100 4032 450176 4060
rect 309100 4020 309106 4032
rect 450170 4020 450176 4032
rect 450228 4020 450234 4072
rect 88242 3952 88248 4004
rect 88300 3992 88306 4004
rect 132586 3992 132592 4004
rect 88300 3964 132592 3992
rect 88300 3952 88306 3964
rect 132586 3952 132592 3964
rect 132644 3952 132650 4004
rect 311802 3952 311808 4004
rect 311860 3992 311866 4004
rect 453666 3992 453672 4004
rect 311860 3964 453672 3992
rect 311860 3952 311866 3964
rect 453666 3952 453672 3964
rect 453724 3952 453730 4004
rect 91002 3884 91008 3936
rect 91060 3924 91066 3936
rect 136082 3924 136088 3936
rect 91060 3896 136088 3924
rect 91060 3884 91066 3896
rect 136082 3884 136088 3896
rect 136140 3884 136146 3936
rect 154577 3927 154635 3933
rect 154577 3893 154589 3927
rect 154623 3924 154635 3927
rect 162302 3924 162308 3936
rect 154623 3896 162308 3924
rect 154623 3893 154635 3896
rect 154577 3887 154635 3893
rect 162302 3884 162308 3896
rect 162360 3884 162366 3936
rect 315942 3884 315948 3936
rect 316000 3924 316006 3936
rect 460842 3924 460848 3936
rect 316000 3896 460848 3924
rect 316000 3884 316006 3896
rect 460842 3884 460848 3896
rect 460900 3884 460906 3936
rect 93762 3816 93768 3868
rect 93820 3856 93826 3868
rect 139670 3856 139676 3868
rect 93820 3828 139676 3856
rect 93820 3816 93826 3828
rect 139670 3816 139676 3828
rect 139728 3816 139734 3868
rect 313182 3816 313188 3868
rect 313240 3856 313246 3868
rect 457254 3856 457260 3868
rect 313240 3828 457260 3856
rect 313240 3816 313246 3828
rect 457254 3816 457260 3828
rect 457312 3816 457318 3868
rect 96522 3748 96528 3800
rect 96580 3788 96586 3800
rect 143258 3788 143264 3800
rect 96580 3760 143264 3788
rect 96580 3748 96586 3760
rect 143258 3748 143264 3760
rect 143316 3748 143322 3800
rect 318702 3748 318708 3800
rect 318760 3788 318766 3800
rect 464430 3788 464436 3800
rect 318760 3760 464436 3788
rect 318760 3748 318766 3760
rect 464430 3748 464436 3760
rect 464488 3748 464494 3800
rect 99282 3680 99288 3732
rect 99340 3720 99346 3732
rect 146846 3720 146852 3732
rect 99340 3692 146852 3720
rect 99340 3680 99346 3692
rect 146846 3680 146852 3692
rect 146904 3680 146910 3732
rect 321462 3680 321468 3732
rect 321520 3720 321526 3732
rect 467834 3720 467840 3732
rect 321520 3692 467840 3720
rect 321520 3680 321526 3692
rect 467834 3680 467840 3692
rect 467892 3680 467898 3732
rect 103422 3612 103428 3664
rect 103480 3652 103486 3664
rect 153930 3652 153936 3664
rect 103480 3624 153936 3652
rect 103480 3612 103486 3624
rect 153930 3612 153936 3624
rect 153988 3612 153994 3664
rect 324222 3612 324228 3664
rect 324280 3652 324286 3664
rect 471514 3652 471520 3664
rect 324280 3624 471520 3652
rect 324280 3612 324286 3624
rect 471514 3612 471520 3624
rect 471572 3612 471578 3664
rect 100662 3544 100668 3596
rect 100720 3584 100726 3596
rect 150434 3584 150440 3596
rect 100720 3556 150440 3584
rect 100720 3544 100726 3556
rect 150434 3544 150440 3556
rect 150492 3544 150498 3596
rect 218146 3544 218152 3596
rect 218204 3584 218210 3596
rect 219342 3584 219348 3596
rect 218204 3556 219348 3584
rect 218204 3544 218210 3556
rect 219342 3544 219348 3556
rect 219400 3544 219406 3596
rect 227714 3544 227720 3596
rect 227772 3584 227778 3596
rect 228910 3584 228916 3596
rect 227772 3556 228916 3584
rect 227772 3544 227778 3556
rect 228910 3544 228916 3556
rect 228968 3544 228974 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 263410 3584 263416 3596
rect 262272 3556 263416 3584
rect 262272 3544 262278 3556
rect 263410 3544 263416 3556
rect 263468 3544 263474 3596
rect 278866 3544 278872 3596
rect 278924 3584 278930 3596
rect 280062 3584 280068 3596
rect 278924 3556 280068 3584
rect 278924 3544 278930 3556
rect 280062 3544 280068 3556
rect 280120 3544 280126 3596
rect 304994 3544 305000 3596
rect 305052 3584 305058 3596
rect 306190 3584 306196 3596
rect 305052 3556 306196 3584
rect 305052 3544 305058 3556
rect 306190 3544 306196 3556
rect 306248 3544 306254 3596
rect 313366 3544 313372 3596
rect 313424 3584 313430 3596
rect 314562 3584 314568 3596
rect 313424 3556 314568 3584
rect 313424 3544 313430 3556
rect 314562 3544 314568 3556
rect 314620 3544 314626 3596
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 325602 3544 325608 3596
rect 325660 3584 325666 3596
rect 475102 3584 475108 3596
rect 325660 3556 475108 3584
rect 325660 3544 325666 3556
rect 475102 3544 475108 3556
rect 475160 3544 475166 3596
rect 502426 3544 502432 3596
rect 502484 3584 502490 3596
rect 503622 3584 503628 3596
rect 502484 3556 503628 3584
rect 502484 3544 502490 3556
rect 503622 3544 503628 3556
rect 503680 3544 503686 3596
rect 518897 3587 518955 3593
rect 518897 3553 518909 3587
rect 518943 3584 518955 3587
rect 528465 3587 528523 3593
rect 528465 3584 528477 3587
rect 518943 3556 528477 3584
rect 518943 3553 518955 3556
rect 518897 3547 518955 3553
rect 528465 3553 528477 3556
rect 528511 3553 528523 3587
rect 528465 3547 528523 3553
rect 536926 3544 536932 3596
rect 536984 3584 536990 3596
rect 538122 3584 538128 3596
rect 536984 3556 538128 3584
rect 536984 3544 536990 3556
rect 538122 3544 538128 3556
rect 538180 3544 538186 3596
rect 568206 3544 568212 3596
rect 568264 3584 568270 3596
rect 568264 3556 572760 3584
rect 568264 3544 568270 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 81434 3516 81440 3528
rect 624 3488 81440 3516
rect 624 3476 630 3488
rect 81434 3476 81440 3488
rect 81492 3476 81498 3528
rect 106182 3476 106188 3528
rect 106240 3516 106246 3528
rect 157518 3516 157524 3528
rect 106240 3488 157524 3516
rect 106240 3476 106246 3488
rect 157518 3476 157524 3488
rect 157576 3476 157582 3528
rect 158714 3476 158720 3528
rect 158772 3516 158778 3528
rect 159910 3516 159916 3528
rect 158772 3488 159916 3516
rect 158772 3476 158778 3488
rect 159910 3476 159916 3488
rect 159968 3476 159974 3528
rect 166994 3476 167000 3528
rect 167052 3516 167058 3528
rect 168190 3516 168196 3528
rect 167052 3488 168196 3516
rect 167052 3476 167058 3488
rect 168190 3476 168196 3488
rect 168248 3476 168254 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 211062 3516 211068 3528
rect 209832 3488 211068 3516
rect 209832 3476 209838 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 328362 3476 328368 3528
rect 328420 3516 328426 3528
rect 478690 3516 478696 3528
rect 328420 3488 478696 3516
rect 328420 3476 328426 3488
rect 478690 3476 478696 3488
rect 478748 3476 478754 3528
rect 509145 3519 509203 3525
rect 509145 3485 509157 3519
rect 509191 3516 509203 3519
rect 511905 3519 511963 3525
rect 511905 3516 511917 3519
rect 509191 3488 511917 3516
rect 509191 3485 509203 3488
rect 509145 3479 509203 3485
rect 511905 3485 511917 3488
rect 511951 3485 511963 3519
rect 559009 3519 559067 3525
rect 559009 3516 559021 3519
rect 511905 3479 511963 3485
rect 529860 3488 559021 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 82906 3448 82912 3460
rect 1728 3420 82912 3448
rect 1728 3408 1734 3420
rect 82906 3408 82912 3420
rect 82964 3408 82970 3460
rect 108942 3408 108948 3460
rect 109000 3448 109006 3460
rect 161106 3448 161112 3460
rect 109000 3420 161112 3448
rect 109000 3408 109006 3420
rect 161106 3408 161112 3420
rect 161164 3408 161170 3460
rect 331122 3408 331128 3460
rect 331180 3448 331186 3460
rect 482278 3448 482284 3460
rect 331180 3420 482284 3448
rect 331180 3408 331186 3420
rect 482278 3408 482284 3420
rect 482336 3408 482342 3460
rect 486513 3451 486571 3457
rect 486513 3417 486525 3451
rect 486559 3448 486571 3451
rect 499577 3451 499635 3457
rect 499577 3448 499589 3451
rect 486559 3420 499589 3448
rect 486559 3417 486571 3420
rect 486513 3411 486571 3417
rect 499577 3417 499589 3420
rect 499623 3417 499635 3451
rect 499577 3411 499635 3417
rect 511997 3451 512055 3457
rect 511997 3417 512009 3451
rect 512043 3448 512055 3451
rect 518897 3451 518955 3457
rect 518897 3448 518909 3451
rect 512043 3420 518909 3448
rect 512043 3417 512055 3420
rect 511997 3411 512055 3417
rect 518897 3417 518909 3420
rect 518943 3417 518955 3451
rect 518897 3411 518955 3417
rect 528465 3451 528523 3457
rect 528465 3417 528477 3451
rect 528511 3448 528523 3451
rect 529860 3448 529888 3488
rect 559009 3485 559021 3488
rect 559055 3485 559067 3519
rect 572732 3516 572760 3556
rect 578602 3516 578608 3528
rect 572732 3488 578608 3516
rect 559009 3479 559067 3485
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 578970 3476 578976 3528
rect 579028 3516 579034 3528
rect 579798 3516 579804 3528
rect 579028 3488 579804 3516
rect 579028 3476 579034 3488
rect 579798 3476 579804 3488
rect 579856 3476 579862 3528
rect 528511 3420 529888 3448
rect 528511 3417 528523 3420
rect 528465 3411 528523 3417
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375190 3380 375196 3392
rect 374052 3352 375196 3380
rect 374052 3340 374058 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 425054 3340 425060 3392
rect 425112 3380 425118 3392
rect 426342 3380 426348 3392
rect 425112 3352 426348 3380
rect 425112 3340 425118 3352
rect 426342 3340 426348 3352
rect 426400 3340 426406 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 499577 3315 499635 3321
rect 499577 3281 499589 3315
rect 499623 3312 499635 3315
rect 509145 3315 509203 3321
rect 509145 3312 509157 3315
rect 499623 3284 509157 3312
rect 499623 3281 499635 3284
rect 499577 3275 499635 3281
rect 509145 3281 509157 3284
rect 509191 3281 509203 3315
rect 509145 3275 509203 3281
rect 559009 3315 559067 3321
rect 559009 3281 559021 3315
rect 559055 3312 559067 3315
rect 582190 3312 582196 3324
rect 559055 3284 582196 3312
rect 559055 3281 559067 3284
rect 559009 3275 559067 3281
rect 582190 3272 582196 3284
rect 582248 3272 582254 3324
rect 578878 3136 578884 3188
rect 578936 3176 578942 3188
rect 580994 3176 581000 3188
rect 578936 3148 581000 3176
rect 578936 3136 578942 3148
rect 580994 3136 581000 3148
rect 581052 3136 581058 3188
rect 287054 1368 287060 1420
rect 287112 1408 287118 1420
rect 288342 1408 288348 1420
rect 287112 1380 288348 1408
rect 287112 1368 287118 1380
rect 288342 1368 288348 1380
rect 288400 1368 288406 1420
rect 126974 552 126980 604
rect 127032 592 127038 604
rect 127802 592 127808 604
rect 127032 564 127808 592
rect 127032 552 127038 564
rect 127802 552 127808 564
rect 127860 552 127866 604
rect 128354 552 128360 604
rect 128412 592 128418 604
rect 128998 592 129004 604
rect 128412 564 129004 592
rect 128412 552 128418 564
rect 128998 552 129004 564
rect 129056 552 129062 604
rect 131114 552 131120 604
rect 131172 592 131178 604
rect 131390 592 131396 604
rect 131172 564 131396 592
rect 131172 552 131178 564
rect 131390 552 131396 564
rect 131448 552 131454 604
rect 200390 552 200396 604
rect 200448 592 200454 604
rect 200482 592 200488 604
rect 200448 564 200488 592
rect 200448 552 200454 564
rect 200482 552 200488 564
rect 200540 552 200546 604
rect 306374 552 306380 604
rect 306432 592 306438 604
rect 307386 592 307392 604
rect 306432 564 307392 592
rect 306432 552 306438 564
rect 307386 552 307392 564
rect 307444 552 307450 604
rect 307754 552 307760 604
rect 307812 592 307818 604
rect 308582 592 308588 604
rect 307812 564 308588 592
rect 307812 552 307818 564
rect 308582 552 308588 564
rect 308640 552 308646 604
rect 309134 552 309140 604
rect 309192 592 309198 604
rect 309778 592 309784 604
rect 309192 564 309784 592
rect 309192 552 309198 564
rect 309778 552 309784 564
rect 309836 552 309842 604
rect 310514 552 310520 604
rect 310572 592 310578 604
rect 310974 592 310980 604
rect 310572 564 310980 592
rect 310572 552 310578 564
rect 310974 552 310980 564
rect 311032 552 311038 604
rect 314654 552 314660 604
rect 314712 592 314718 604
rect 315758 592 315764 604
rect 314712 564 315764 592
rect 314712 552 314718 564
rect 315758 552 315764 564
rect 315816 552 315822 604
rect 517882 592 517888 604
rect 517843 564 517888 592
rect 517882 552 517888 564
rect 517940 552 517946 604
rect 519078 592 519084 604
rect 519039 564 519084 592
rect 519078 552 519084 564
rect 519136 552 519142 604
rect 545298 592 545304 604
rect 545259 564 545304 592
rect 545298 552 545304 564
rect 545356 552 545362 604
rect 548886 592 548892 604
rect 548847 564 548892 592
rect 548886 552 548892 564
rect 548944 552 548950 604
rect 550082 592 550088 604
rect 550043 564 550088 592
rect 550082 552 550088 564
rect 550140 552 550146 604
rect 576854 552 576860 604
rect 576912 592 576918 604
rect 577406 592 577412 604
rect 576912 564 577412 592
rect 576912 552 576918 564
rect 577406 552 577412 564
rect 577464 552 577470 604
<< via1 >>
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 283288 698232 283340 698284
rect 283932 698232 283984 698284
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 201500 697552 201552 697604
rect 202788 697552 202840 697604
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 331220 697552 331272 697604
rect 332508 697552 332560 697604
rect 567844 696940 567896 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 72700 694084 72752 694136
rect 283104 694084 283156 694136
rect 283288 694084 283340 694136
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 218060 692792 218112 692844
rect 219072 692792 219124 692844
rect 234620 692792 234672 692844
rect 235264 692792 235316 692844
rect 347780 692792 347832 692844
rect 348884 692792 348936 692844
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 283104 692724 283156 692776
rect 283288 692724 283340 692776
rect 412824 692724 412876 692776
rect 542544 692724 542596 692776
rect 542728 692724 542780 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 154396 685788 154448 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 299480 684428 299532 684480
rect 300124 684428 300176 684480
rect 429200 684428 429252 684480
rect 429844 684428 429896 684480
rect 558920 684428 558972 684480
rect 559656 684428 559708 684480
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 282920 683068 282972 683120
rect 299480 683068 299532 683120
rect 412640 683068 412692 683120
rect 429200 683068 429252 683120
rect 542360 683068 542412 683120
rect 558920 683068 558972 683120
rect 3516 681708 3568 681760
rect 8944 681708 8996 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 218060 673480 218112 673532
rect 218244 673480 218296 673532
rect 234620 673480 234672 673532
rect 234804 673480 234856 673532
rect 347780 673480 347832 673532
rect 347964 673480 348016 673532
rect 364340 673480 364392 673532
rect 364524 673480 364576 673532
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 494060 673480 494112 673532
rect 494244 673480 494296 673532
rect 558184 673480 558236 673532
rect 580172 673480 580224 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 283380 666544 283432 666596
rect 299940 666544 299992 666596
rect 413100 666544 413152 666596
rect 429660 666544 429712 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 73068 656820 73120 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 218060 654100 218112 654152
rect 218244 654100 218296 654152
rect 234620 654100 234672 654152
rect 234804 654100 234856 654152
rect 347780 654100 347832 654152
rect 347964 654100 348016 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 14464 652740 14516 652792
rect 566464 650020 566516 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 283104 647232 283156 647284
rect 283196 647232 283248 647284
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 72976 640364 73028 640416
rect 283104 640364 283156 640416
rect 283196 640364 283248 640416
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 72792 640228 72844 640280
rect 573364 638936 573416 638988
rect 580172 638936 580224 638988
rect 72792 637508 72844 637560
rect 72884 637508 72936 637560
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 218060 634788 218112 634840
rect 218244 634788 218296 634840
rect 234620 634788 234672 634840
rect 234804 634788 234856 634840
rect 347780 634788 347832 634840
rect 347964 634788 348016 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 283012 630640 283064 630692
rect 283196 630640 283248 630692
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 556804 626560 556856 626612
rect 580172 626560 580224 626612
rect 73068 626535 73120 626544
rect 73068 626501 73077 626535
rect 73077 626501 73111 626535
rect 73111 626501 73120 626535
rect 73068 626492 73120 626501
rect 3240 623772 3292 623824
rect 29644 623772 29696 623824
rect 73068 616879 73120 616888
rect 73068 616845 73077 616879
rect 73077 616845 73111 616879
rect 73111 616845 73120 616879
rect 73068 616836 73120 616845
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 218060 615476 218112 615528
rect 218244 615476 218296 615528
rect 234620 615476 234672 615528
rect 234804 615476 234856 615528
rect 347780 615476 347832 615528
rect 347964 615476 348016 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 477500 615476 477552 615528
rect 477684 615476 477736 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 73068 611396 73120 611448
rect 283012 611328 283064 611380
rect 283196 611328 283248 611380
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 72884 611260 72936 611312
rect 283104 608583 283156 608592
rect 283104 608549 283113 608583
rect 283113 608549 283147 608583
rect 283147 608549 283156 608583
rect 283104 608540 283156 608549
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 412824 608583 412876 608592
rect 412824 608549 412833 608583
rect 412833 608549 412867 608583
rect 412867 608549 412876 608583
rect 412824 608540 412876 608549
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 542544 608583 542596 608592
rect 542544 608549 542553 608583
rect 542553 608549 542587 608583
rect 542587 608549 542596 608583
rect 542544 608540 542596 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 565084 603100 565136 603152
rect 580172 603100 580224 603152
rect 283288 601672 283340 601724
rect 299848 601672 299900 601724
rect 413008 601672 413060 601724
rect 429568 601672 429620 601724
rect 542728 601672 542780 601724
rect 559288 601672 559340 601724
rect 72976 601536 73028 601588
rect 73160 601536 73212 601588
rect 72976 598884 73028 598936
rect 283288 598927 283340 598936
rect 283288 598893 283297 598927
rect 283297 598893 283331 598927
rect 283331 598893 283340 598927
rect 283288 598884 283340 598893
rect 299848 598927 299900 598936
rect 299848 598893 299857 598927
rect 299857 598893 299891 598927
rect 299891 598893 299900 598927
rect 299848 598884 299900 598893
rect 413008 598927 413060 598936
rect 413008 598893 413017 598927
rect 413017 598893 413051 598927
rect 413051 598893 413060 598927
rect 413008 598884 413060 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 542728 598927 542780 598936
rect 542728 598893 542737 598927
rect 542737 598893 542771 598927
rect 542771 598893 542780 598927
rect 542728 598884 542780 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 137744 596164 137796 596216
rect 137928 596164 137980 596216
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 218060 596164 218112 596216
rect 218244 596164 218296 596216
rect 234620 596164 234672 596216
rect 234804 596164 234856 596216
rect 347780 596164 347832 596216
rect 347964 596164 348016 596216
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 477500 596164 477552 596216
rect 477684 596164 477736 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3332 594804 3384 594856
rect 44824 594804 44876 594856
rect 570604 592016 570656 592068
rect 580172 592016 580224 592068
rect 72884 589339 72936 589348
rect 72884 589305 72893 589339
rect 72893 589305 72927 589339
rect 72927 589305 72936 589339
rect 72884 589296 72936 589305
rect 283380 589296 283432 589348
rect 299940 589296 299992 589348
rect 413100 589296 413152 589348
rect 429660 589296 429712 589348
rect 542820 589296 542872 589348
rect 559380 589296 559432 589348
rect 8024 589271 8076 589280
rect 8024 589237 8033 589271
rect 8033 589237 8067 589271
rect 8067 589237 8076 589271
rect 8024 589228 8076 589237
rect 137744 589271 137796 589280
rect 137744 589237 137753 589271
rect 137753 589237 137787 589271
rect 137787 589237 137796 589271
rect 137744 589228 137796 589237
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 218152 589228 218204 589280
rect 234712 589228 234764 589280
rect 347872 589228 347924 589280
rect 364432 589228 364484 589280
rect 477592 589228 477644 589280
rect 494152 589228 494204 589280
rect 72700 582360 72752 582412
rect 72884 582360 72936 582412
rect 283380 582428 283432 582480
rect 299940 582428 299992 582480
rect 413100 582428 413152 582480
rect 429660 582428 429712 582480
rect 542820 582428 542872 582480
rect 559380 582428 559432 582480
rect 283288 582292 283340 582344
rect 299848 582292 299900 582344
rect 413008 582292 413060 582344
rect 429568 582292 429620 582344
rect 542728 582292 542780 582344
rect 559288 582292 559340 582344
rect 8024 579751 8076 579760
rect 8024 579717 8033 579751
rect 8033 579717 8067 579751
rect 8067 579717 8076 579751
rect 8024 579708 8076 579717
rect 137744 579751 137796 579760
rect 137744 579717 137753 579751
rect 137753 579717 137787 579751
rect 137787 579717 137796 579751
rect 137744 579708 137796 579717
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 218060 579683 218112 579692
rect 218060 579649 218069 579683
rect 218069 579649 218103 579683
rect 218103 579649 218112 579683
rect 218060 579640 218112 579649
rect 234620 579683 234672 579692
rect 234620 579649 234629 579683
rect 234629 579649 234663 579683
rect 234663 579649 234672 579683
rect 234620 579640 234672 579649
rect 347780 579683 347832 579692
rect 347780 579649 347789 579683
rect 347789 579649 347823 579683
rect 347823 579649 347832 579683
rect 364340 579683 364392 579692
rect 347780 579640 347832 579649
rect 364340 579649 364349 579683
rect 364349 579649 364383 579683
rect 364383 579649 364392 579683
rect 364340 579640 364392 579649
rect 477500 579683 477552 579692
rect 477500 579649 477509 579683
rect 477509 579649 477543 579683
rect 477543 579649 477552 579683
rect 477500 579640 477552 579649
rect 494060 579683 494112 579692
rect 494060 579649 494069 579683
rect 494069 579649 494103 579683
rect 494103 579649 494112 579683
rect 494060 579640 494112 579649
rect 555424 579640 555476 579692
rect 580172 579640 580224 579692
rect 7932 579572 7984 579624
rect 8116 579572 8168 579624
rect 72700 579572 72752 579624
rect 137652 579572 137704 579624
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 72608 569959 72660 569968
rect 72608 569925 72617 569959
rect 72617 569925 72651 569959
rect 72651 569925 72660 569959
rect 72608 569916 72660 569925
rect 137560 569959 137612 569968
rect 137560 569925 137569 569959
rect 137569 569925 137603 569959
rect 137603 569925 137612 569959
rect 137560 569916 137612 569925
rect 218152 569891 218204 569900
rect 218152 569857 218161 569891
rect 218161 569857 218195 569891
rect 218195 569857 218204 569891
rect 218152 569848 218204 569857
rect 234712 569891 234764 569900
rect 234712 569857 234721 569891
rect 234721 569857 234755 569891
rect 234755 569857 234764 569891
rect 234712 569848 234764 569857
rect 347872 569891 347924 569900
rect 347872 569857 347881 569891
rect 347881 569857 347915 569891
rect 347915 569857 347924 569891
rect 347872 569848 347924 569857
rect 364432 569891 364484 569900
rect 364432 569857 364441 569891
rect 364441 569857 364475 569891
rect 364475 569857 364484 569891
rect 364432 569848 364484 569857
rect 477592 569891 477644 569900
rect 477592 569857 477601 569891
rect 477601 569857 477635 569891
rect 477635 569857 477644 569891
rect 477592 569848 477644 569857
rect 494152 569891 494204 569900
rect 494152 569857 494161 569891
rect 494161 569857 494195 569891
rect 494195 569857 494204 569891
rect 494152 569848 494204 569857
rect 4068 567196 4120 567248
rect 13084 567196 13136 567248
rect 283012 563116 283064 563168
rect 412732 563116 412784 563168
rect 429292 563116 429344 563168
rect 542452 563116 542504 563168
rect 559012 563116 559064 563168
rect 72608 563048 72660 563100
rect 137560 563048 137612 563100
rect 218336 563048 218388 563100
rect 234896 563048 234948 563100
rect 7932 562912 7984 562964
rect 8116 562912 8168 562964
rect 72700 562912 72752 562964
rect 348056 563048 348108 563100
rect 364616 563048 364668 563100
rect 477776 563048 477828 563100
rect 494336 563048 494388 563100
rect 283012 562980 283064 563032
rect 412732 562980 412784 563032
rect 429292 562980 429344 563032
rect 542452 562980 542504 563032
rect 559012 562980 559064 563032
rect 137652 562912 137704 562964
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 137652 560235 137704 560244
rect 137652 560201 137661 560235
rect 137661 560201 137695 560235
rect 137695 560201 137704 560235
rect 137652 560192 137704 560201
rect 283012 560235 283064 560244
rect 283012 560201 283021 560235
rect 283021 560201 283055 560235
rect 283055 560201 283064 560235
rect 283012 560192 283064 560201
rect 412732 560235 412784 560244
rect 412732 560201 412741 560235
rect 412741 560201 412775 560235
rect 412775 560201 412784 560235
rect 412732 560192 412784 560201
rect 429292 560235 429344 560244
rect 429292 560201 429301 560235
rect 429301 560201 429335 560235
rect 429335 560201 429344 560235
rect 429292 560192 429344 560201
rect 542452 560235 542504 560244
rect 542452 560201 542461 560235
rect 542461 560201 542495 560235
rect 542495 560201 542504 560235
rect 542452 560192 542504 560201
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 563704 556180 563756 556232
rect 580172 556180 580224 556232
rect 72608 553435 72660 553444
rect 72608 553401 72617 553435
rect 72617 553401 72651 553435
rect 72651 553401 72660 553435
rect 72608 553392 72660 553401
rect 72608 550647 72660 550656
rect 72608 550613 72617 550647
rect 72617 550613 72651 550647
rect 72651 550613 72660 550647
rect 72608 550604 72660 550613
rect 137836 550604 137888 550656
rect 218152 550604 218204 550656
rect 218428 550604 218480 550656
rect 234712 550604 234764 550656
rect 234988 550604 235040 550656
rect 283196 550604 283248 550656
rect 299480 550604 299532 550656
rect 299756 550604 299808 550656
rect 347872 550604 347924 550656
rect 348148 550604 348200 550656
rect 364432 550604 364484 550656
rect 364708 550604 364760 550656
rect 412916 550604 412968 550656
rect 429476 550604 429528 550656
rect 477592 550604 477644 550656
rect 477868 550604 477920 550656
rect 494152 550604 494204 550656
rect 494428 550604 494480 550656
rect 542636 550604 542688 550656
rect 559196 550604 559248 550656
rect 8024 550579 8076 550588
rect 8024 550545 8033 550579
rect 8033 550545 8067 550579
rect 8067 550545 8076 550579
rect 8024 550536 8076 550545
rect 552664 545096 552716 545148
rect 580172 545096 580224 545148
rect 72608 543736 72660 543788
rect 218428 543804 218480 543856
rect 234988 543804 235040 543856
rect 299480 543736 299532 543788
rect 218336 543668 218388 543720
rect 234896 543668 234948 543720
rect 72700 543600 72752 543652
rect 137652 543600 137704 543652
rect 137836 543600 137888 543652
rect 283012 543600 283064 543652
rect 283196 543600 283248 543652
rect 348148 543804 348200 543856
rect 364708 543804 364760 543856
rect 477868 543804 477920 543856
rect 494428 543804 494480 543856
rect 348056 543668 348108 543720
rect 364616 543668 364668 543720
rect 477776 543668 477828 543720
rect 494336 543668 494388 543720
rect 299572 543600 299624 543652
rect 412732 543600 412784 543652
rect 412916 543600 412968 543652
rect 429292 543600 429344 543652
rect 429476 543600 429528 543652
rect 542452 543600 542504 543652
rect 542636 543600 542688 543652
rect 559012 543600 559064 543652
rect 559196 543600 559248 543652
rect 8208 540948 8260 541000
rect 4068 538228 4120 538280
rect 17224 538228 17276 538280
rect 72608 534123 72660 534132
rect 72608 534089 72617 534123
rect 72617 534089 72651 534123
rect 72651 534089 72660 534123
rect 72608 534080 72660 534089
rect 137652 534012 137704 534064
rect 137836 534012 137888 534064
rect 283012 534012 283064 534064
rect 283196 534012 283248 534064
rect 299572 534012 299624 534064
rect 299756 534012 299808 534064
rect 412732 534012 412784 534064
rect 412916 534012 412968 534064
rect 429292 534012 429344 534064
rect 429476 534012 429528 534064
rect 542452 534012 542504 534064
rect 542636 534012 542688 534064
rect 559012 534012 559064 534064
rect 559196 534012 559248 534064
rect 72608 531335 72660 531344
rect 72608 531301 72617 531335
rect 72617 531301 72651 531335
rect 72651 531301 72660 531335
rect 72608 531292 72660 531301
rect 218152 531292 218204 531344
rect 218428 531292 218480 531344
rect 234712 531292 234764 531344
rect 234988 531292 235040 531344
rect 347872 531292 347924 531344
rect 348148 531292 348200 531344
rect 364432 531292 364484 531344
rect 364708 531292 364760 531344
rect 477592 531292 477644 531344
rect 477868 531292 477920 531344
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 218428 524492 218480 524544
rect 234988 524492 235040 524544
rect 283196 524424 283248 524476
rect 299756 524424 299808 524476
rect 218336 524356 218388 524408
rect 234896 524356 234948 524408
rect 283288 524356 283340 524408
rect 348148 524492 348200 524544
rect 364708 524492 364760 524544
rect 412916 524424 412968 524476
rect 429476 524424 429528 524476
rect 299848 524356 299900 524408
rect 348056 524356 348108 524408
rect 364616 524356 364668 524408
rect 413008 524356 413060 524408
rect 477868 524492 477920 524544
rect 494428 524492 494480 524544
rect 542636 524424 542688 524476
rect 559196 524424 559248 524476
rect 429568 524356 429620 524408
rect 477776 524356 477828 524408
rect 494336 524356 494388 524408
rect 542728 524356 542780 524408
rect 559288 524356 559340 524408
rect 72700 524288 72752 524340
rect 72884 524288 72936 524340
rect 8208 521636 8260 521688
rect 8392 521636 8444 521688
rect 137928 521636 137980 521688
rect 138112 521636 138164 521688
rect 154488 521636 154540 521688
rect 218152 511980 218204 512032
rect 218428 511980 218480 512032
rect 234712 511980 234764 512032
rect 234988 511980 235040 512032
rect 283104 511980 283156 512032
rect 283380 511980 283432 512032
rect 299664 511980 299716 512032
rect 299940 511980 299992 512032
rect 347872 511980 347924 512032
rect 348148 511980 348200 512032
rect 364432 511980 364484 512032
rect 364708 511980 364760 512032
rect 412824 511980 412876 512032
rect 413100 511980 413152 512032
rect 429384 511980 429436 512032
rect 429660 511980 429712 512032
rect 477592 511980 477644 512032
rect 477868 511980 477920 512032
rect 494152 511980 494204 512032
rect 494428 511980 494480 512032
rect 542544 511980 542596 512032
rect 542820 511980 542872 512032
rect 559104 511980 559156 512032
rect 559380 511980 559432 512032
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 3884 509260 3936 509312
rect 39304 509260 39356 509312
rect 551284 509260 551336 509312
rect 580172 509260 580224 509312
rect 8208 502324 8260 502376
rect 8392 502324 8444 502376
rect 72608 502324 72660 502376
rect 73068 502324 73120 502376
rect 137928 502324 137980 502376
rect 138112 502324 138164 502376
rect 154488 502324 154540 502376
rect 218244 502324 218296 502376
rect 218428 502324 218480 502376
rect 234804 502324 234856 502376
rect 234988 502324 235040 502376
rect 283196 502324 283248 502376
rect 283380 502324 283432 502376
rect 299756 502324 299808 502376
rect 299940 502324 299992 502376
rect 347964 502324 348016 502376
rect 348148 502324 348200 502376
rect 364524 502324 364576 502376
rect 364708 502324 364760 502376
rect 412916 502324 412968 502376
rect 413100 502324 413152 502376
rect 429476 502324 429528 502376
rect 429660 502324 429712 502376
rect 477684 502324 477736 502376
rect 477868 502324 477920 502376
rect 494244 502324 494296 502376
rect 494428 502324 494480 502376
rect 542636 502324 542688 502376
rect 542820 502324 542872 502376
rect 559196 502324 559248 502376
rect 559380 502324 559432 502376
rect 569224 498176 569276 498228
rect 580172 498176 580224 498228
rect 7932 492600 7984 492652
rect 8116 492600 8168 492652
rect 137652 492600 137704 492652
rect 137836 492600 137888 492652
rect 154212 492600 154264 492652
rect 154396 492600 154448 492652
rect 283104 492643 283156 492652
rect 283104 492609 283113 492643
rect 283113 492609 283147 492643
rect 283147 492609 283156 492643
rect 283104 492600 283156 492609
rect 299664 492643 299716 492652
rect 299664 492609 299673 492643
rect 299673 492609 299707 492643
rect 299707 492609 299716 492643
rect 299664 492600 299716 492609
rect 412824 492643 412876 492652
rect 412824 492609 412833 492643
rect 412833 492609 412867 492643
rect 412867 492609 412876 492643
rect 412824 492600 412876 492609
rect 429384 492643 429436 492652
rect 429384 492609 429393 492643
rect 429393 492609 429427 492643
rect 429427 492609 429436 492643
rect 429384 492600 429436 492609
rect 542544 492643 542596 492652
rect 542544 492609 542553 492643
rect 542553 492609 542587 492643
rect 542587 492609 542596 492643
rect 542544 492600 542596 492609
rect 559104 492643 559156 492652
rect 559104 492609 559113 492643
rect 559113 492609 559147 492643
rect 559147 492609 559156 492643
rect 559104 492600 559156 492609
rect 554044 485800 554096 485852
rect 579896 485800 579948 485852
rect 283104 485775 283156 485784
rect 283104 485741 283113 485775
rect 283113 485741 283147 485775
rect 283147 485741 283156 485775
rect 283104 485732 283156 485741
rect 299664 485775 299716 485784
rect 299664 485741 299673 485775
rect 299673 485741 299707 485775
rect 299707 485741 299716 485775
rect 299664 485732 299716 485741
rect 412824 485775 412876 485784
rect 412824 485741 412833 485775
rect 412833 485741 412867 485775
rect 412867 485741 412876 485775
rect 412824 485732 412876 485741
rect 429384 485775 429436 485784
rect 429384 485741 429393 485775
rect 429393 485741 429427 485775
rect 429427 485741 429436 485775
rect 429384 485732 429436 485741
rect 542544 485775 542596 485784
rect 542544 485741 542553 485775
rect 542553 485741 542587 485775
rect 542587 485741 542596 485775
rect 542544 485732 542596 485741
rect 559104 485775 559156 485784
rect 559104 485741 559113 485775
rect 559113 485741 559147 485775
rect 559147 485741 559156 485775
rect 559104 485732 559156 485741
rect 3148 480224 3200 480276
rect 10324 480224 10376 480276
rect 72884 480224 72936 480276
rect 73068 480224 73120 480276
rect 218060 480224 218112 480276
rect 218244 480224 218296 480276
rect 234620 480224 234672 480276
rect 234804 480224 234856 480276
rect 347780 480224 347832 480276
rect 347964 480224 348016 480276
rect 364340 480224 364392 480276
rect 364524 480224 364576 480276
rect 477500 480224 477552 480276
rect 477684 480224 477736 480276
rect 494060 480224 494112 480276
rect 494244 480224 494296 480276
rect 283012 476076 283064 476128
rect 283196 476076 283248 476128
rect 299572 476076 299624 476128
rect 299756 476076 299808 476128
rect 412732 476076 412784 476128
rect 412916 476076 412968 476128
rect 429292 476076 429344 476128
rect 429476 476076 429528 476128
rect 542452 476076 542504 476128
rect 542636 476076 542688 476128
rect 559012 476076 559064 476128
rect 559196 476076 559248 476128
rect 8024 473288 8076 473340
rect 8116 473288 8168 473340
rect 137468 473288 137520 473340
rect 137744 473288 137796 473340
rect 283104 473331 283156 473340
rect 283104 473297 283113 473331
rect 283113 473297 283147 473331
rect 283147 473297 283156 473331
rect 283104 473288 283156 473297
rect 299664 473331 299716 473340
rect 299664 473297 299673 473331
rect 299673 473297 299707 473331
rect 299707 473297 299716 473331
rect 299664 473288 299716 473297
rect 412824 473331 412876 473340
rect 412824 473297 412833 473331
rect 412833 473297 412867 473331
rect 412867 473297 412876 473331
rect 412824 473288 412876 473297
rect 429384 473331 429436 473340
rect 429384 473297 429393 473331
rect 429393 473297 429427 473331
rect 429427 473297 429436 473331
rect 429384 473288 429436 473297
rect 542544 473331 542596 473340
rect 542544 473297 542553 473331
rect 542553 473297 542587 473331
rect 542587 473297 542596 473331
rect 542544 473288 542596 473297
rect 559104 473331 559156 473340
rect 559104 473297 559113 473331
rect 559113 473297 559147 473331
rect 559147 473297 559156 473331
rect 559104 473288 559156 473297
rect 154304 466420 154356 466472
rect 154488 466420 154540 466472
rect 283104 466395 283156 466404
rect 283104 466361 283113 466395
rect 283113 466361 283147 466395
rect 283147 466361 283156 466395
rect 283104 466352 283156 466361
rect 299664 466395 299716 466404
rect 299664 466361 299673 466395
rect 299673 466361 299707 466395
rect 299707 466361 299716 466395
rect 299664 466352 299716 466361
rect 412824 466395 412876 466404
rect 412824 466361 412833 466395
rect 412833 466361 412867 466395
rect 412867 466361 412876 466395
rect 412824 466352 412876 466361
rect 429384 466395 429436 466404
rect 429384 466361 429393 466395
rect 429393 466361 429427 466395
rect 429427 466361 429436 466395
rect 429384 466352 429436 466361
rect 542544 466395 542596 466404
rect 542544 466361 542553 466395
rect 542553 466361 542587 466395
rect 542587 466361 542596 466395
rect 542544 466352 542596 466361
rect 559104 466395 559156 466404
rect 559104 466361 559113 466395
rect 559113 466361 559147 466395
rect 559147 466361 559156 466395
rect 559104 466352 559156 466361
rect 571984 462340 572036 462392
rect 580172 462340 580224 462392
rect 72884 460912 72936 460964
rect 73068 460912 73120 460964
rect 218060 460912 218112 460964
rect 218244 460912 218296 460964
rect 234620 460912 234672 460964
rect 234804 460912 234856 460964
rect 347780 460912 347832 460964
rect 347964 460912 348016 460964
rect 364340 460912 364392 460964
rect 364524 460912 364576 460964
rect 477500 460912 477552 460964
rect 477684 460912 477736 460964
rect 494060 460912 494112 460964
rect 494244 460912 494296 460964
rect 299572 453951 299624 453960
rect 299572 453917 299581 453951
rect 299581 453917 299615 453951
rect 299615 453917 299624 453951
rect 299572 453908 299624 453917
rect 3056 451256 3108 451308
rect 6184 451256 6236 451308
rect 8024 447108 8076 447160
rect 137744 447108 137796 447160
rect 154304 447108 154356 447160
rect 282920 447108 282972 447160
rect 412640 447108 412692 447160
rect 429200 447108 429252 447160
rect 542360 447108 542412 447160
rect 558920 447108 558972 447160
rect 8116 447040 8168 447092
rect 137836 447040 137888 447092
rect 154396 447040 154448 447092
rect 283012 447040 283064 447092
rect 299572 447083 299624 447092
rect 299572 447049 299581 447083
rect 299581 447049 299615 447083
rect 299615 447049 299624 447083
rect 299572 447040 299624 447049
rect 412732 447040 412784 447092
rect 429292 447040 429344 447092
rect 542452 447040 542504 447092
rect 559012 447040 559064 447092
rect 8116 444363 8168 444372
rect 8116 444329 8125 444363
rect 8125 444329 8159 444363
rect 8159 444329 8168 444363
rect 8116 444320 8168 444329
rect 137836 444363 137888 444372
rect 137836 444329 137845 444363
rect 137845 444329 137879 444363
rect 137879 444329 137888 444363
rect 137836 444320 137888 444329
rect 154396 444363 154448 444372
rect 154396 444329 154405 444363
rect 154405 444329 154439 444363
rect 154439 444329 154448 444363
rect 154396 444320 154448 444329
rect 218060 441600 218112 441652
rect 218244 441600 218296 441652
rect 234620 441600 234672 441652
rect 234804 441600 234856 441652
rect 347780 441600 347832 441652
rect 347964 441600 348016 441652
rect 364340 441600 364392 441652
rect 364524 441600 364576 441652
rect 477500 441600 477552 441652
rect 477684 441600 477736 441652
rect 494060 441600 494112 441652
rect 494244 441600 494296 441652
rect 560944 438880 560996 438932
rect 580172 438880 580224 438932
rect 72792 437452 72844 437504
rect 72976 437452 73028 437504
rect 8116 437427 8168 437436
rect 8116 437393 8125 437427
rect 8125 437393 8159 437427
rect 8159 437393 8168 437427
rect 8116 437384 8168 437393
rect 137836 437427 137888 437436
rect 137836 437393 137845 437427
rect 137845 437393 137879 437427
rect 137879 437393 137888 437427
rect 137836 437384 137888 437393
rect 154396 437427 154448 437436
rect 154396 437393 154405 437427
rect 154405 437393 154439 437427
rect 154439 437393 154448 437427
rect 154396 437384 154448 437393
rect 283104 434707 283156 434716
rect 283104 434673 283113 434707
rect 283113 434673 283147 434707
rect 283147 434673 283156 434707
rect 283104 434664 283156 434673
rect 299664 434707 299716 434716
rect 299664 434673 299673 434707
rect 299673 434673 299707 434707
rect 299707 434673 299716 434707
rect 299664 434664 299716 434673
rect 412824 434707 412876 434716
rect 412824 434673 412833 434707
rect 412833 434673 412867 434707
rect 412867 434673 412876 434707
rect 412824 434664 412876 434673
rect 429384 434707 429436 434716
rect 429384 434673 429393 434707
rect 429393 434673 429427 434707
rect 429427 434673 429436 434707
rect 429384 434664 429436 434673
rect 542544 434707 542596 434716
rect 542544 434673 542553 434707
rect 542553 434673 542587 434707
rect 542587 434673 542596 434707
rect 542544 434664 542596 434673
rect 559104 434707 559156 434716
rect 559104 434673 559113 434707
rect 559113 434673 559147 434707
rect 559147 434673 559156 434707
rect 559104 434664 559156 434673
rect 283104 427771 283156 427780
rect 283104 427737 283113 427771
rect 283113 427737 283147 427771
rect 283147 427737 283156 427771
rect 283104 427728 283156 427737
rect 299664 427771 299716 427780
rect 299664 427737 299673 427771
rect 299673 427737 299707 427771
rect 299707 427737 299716 427771
rect 299664 427728 299716 427737
rect 412824 427771 412876 427780
rect 412824 427737 412833 427771
rect 412833 427737 412867 427771
rect 412867 427737 412876 427771
rect 412824 427728 412876 427737
rect 429384 427771 429436 427780
rect 429384 427737 429393 427771
rect 429393 427737 429427 427771
rect 429427 427737 429436 427771
rect 429384 427728 429436 427737
rect 542544 427771 542596 427780
rect 542544 427737 542553 427771
rect 542553 427737 542587 427771
rect 542587 427737 542596 427771
rect 542544 427728 542596 427737
rect 559104 427771 559156 427780
rect 559104 427737 559113 427771
rect 559113 427737 559147 427771
rect 559147 427737 559156 427771
rect 559104 427728 559156 427737
rect 8024 425076 8076 425128
rect 8208 425076 8260 425128
rect 137744 425076 137796 425128
rect 137928 425076 137980 425128
rect 154304 425076 154356 425128
rect 154488 425076 154540 425128
rect 300032 424872 300084 424924
rect 397460 424872 397512 424924
rect 311808 424804 311860 424856
rect 412916 424804 412968 424856
rect 323584 424736 323636 424788
rect 429476 424736 429528 424788
rect 335452 424668 335504 424720
rect 462320 424668 462372 424720
rect 347228 424600 347280 424652
rect 477684 424600 477736 424652
rect 72792 424532 72844 424584
rect 123208 424532 123260 424584
rect 252928 424532 252980 424584
rect 299756 424532 299808 424584
rect 359004 424532 359056 424584
rect 494244 424532 494296 424584
rect 41328 424464 41380 424516
rect 111432 424464 111484 424516
rect 264704 424464 264756 424516
rect 331220 424464 331272 424516
rect 370780 424464 370832 424516
rect 527180 424464 527232 424516
rect 24768 424396 24820 424448
rect 99656 424396 99708 424448
rect 106188 424396 106240 424448
rect 146760 424396 146812 424448
rect 154304 424396 154356 424448
rect 170404 424396 170456 424448
rect 205732 424396 205784 424448
rect 218244 424396 218296 424448
rect 229284 424396 229336 424448
rect 266360 424396 266412 424448
rect 276480 424396 276532 424448
rect 347964 424396 348016 424448
rect 382556 424396 382608 424448
rect 542636 424396 542688 424448
rect 8024 424328 8076 424380
rect 87880 424328 87932 424380
rect 89628 424328 89680 424380
rect 134984 424328 135036 424380
rect 137744 424328 137796 424380
rect 158536 424328 158588 424380
rect 171048 424328 171100 424380
rect 182180 424328 182232 424380
rect 217508 424328 217560 424380
rect 234804 424328 234856 424380
rect 241060 424328 241112 424380
rect 283196 424328 283248 424380
rect 288256 424328 288308 424380
rect 364524 424328 364576 424380
rect 394332 424328 394384 424380
rect 559196 424328 559248 424380
rect 3332 423648 3384 423700
rect 7564 423648 7616 423700
rect 193956 423648 194008 423700
rect 201500 423648 201552 423700
rect 8944 419432 8996 419484
rect 78680 419432 78732 419484
rect 401600 419432 401652 419484
rect 567844 419432 567896 419484
rect 425704 415420 425756 415472
rect 580172 415420 580224 415472
rect 401600 412564 401652 412616
rect 580264 412564 580316 412616
rect 3424 411204 3476 411256
rect 78680 411204 78732 411256
rect 401600 405628 401652 405680
rect 558184 405628 558236 405680
rect 14464 404268 14516 404320
rect 78680 404268 78732 404320
rect 401600 398760 401652 398812
rect 566464 398760 566516 398812
rect 29644 395972 29696 396024
rect 78680 395972 78732 396024
rect 3148 394680 3200 394732
rect 21364 394680 21416 394732
rect 407764 391960 407816 392012
rect 580172 391960 580224 392012
rect 401600 390464 401652 390516
rect 573364 390464 573416 390516
rect 3516 389104 3568 389156
rect 78680 389104 78732 389156
rect 401600 383596 401652 383648
rect 556804 383596 556856 383648
rect 44824 380808 44876 380860
rect 78680 380808 78732 380860
rect 401600 376660 401652 376712
rect 565084 376660 565136 376712
rect 13084 373940 13136 373992
rect 78680 373940 78732 373992
rect 401600 369792 401652 369844
rect 570604 369792 570656 369844
rect 576124 368500 576176 368552
rect 580172 368500 580224 368552
rect 3608 365644 3660 365696
rect 78680 365644 78732 365696
rect 401600 362856 401652 362908
rect 555424 362856 555476 362908
rect 17224 358708 17276 358760
rect 78680 358708 78732 358760
rect 405004 357416 405056 357468
rect 579896 357416 579948 357468
rect 401600 355988 401652 356040
rect 563704 355988 563756 356040
rect 39304 350480 39356 350532
rect 78680 350480 78732 350532
rect 401600 347692 401652 347744
rect 552664 347692 552716 347744
rect 403624 345040 403676 345092
rect 580172 345040 580224 345092
rect 3700 343544 3752 343596
rect 78680 343544 78732 343596
rect 401600 340824 401652 340876
rect 578884 340824 578936 340876
rect 3056 336744 3108 336796
rect 37924 336744 37976 336796
rect 10324 335248 10376 335300
rect 78680 335248 78732 335300
rect 401600 333888 401652 333940
rect 551284 333888 551336 333940
rect 6184 327020 6236 327072
rect 78680 327020 78732 327072
rect 401600 327020 401652 327072
rect 569224 327020 569276 327072
rect 3792 320084 3844 320136
rect 78680 320084 78732 320136
rect 401600 320084 401652 320136
rect 554044 320084 554096 320136
rect 401600 313216 401652 313268
rect 571984 313216 572036 313268
rect 7564 311788 7616 311840
rect 78680 311788 78732 311840
rect 409144 310496 409196 310548
rect 579620 310496 579672 310548
rect 402244 305600 402296 305652
rect 578884 305600 578936 305652
rect 21364 304920 21416 304972
rect 78680 304920 78732 304972
rect 401600 304920 401652 304972
rect 580356 304920 580408 304972
rect 401600 298052 401652 298104
rect 560944 298052 560996 298104
rect 3424 296624 3476 296676
rect 78680 296624 78732 296676
rect 401600 291116 401652 291168
rect 425704 291116 425756 291168
rect 3516 289756 3568 289808
rect 78680 289756 78732 289808
rect 401600 284248 401652 284300
rect 580264 284248 580316 284300
rect 37924 281460 37976 281512
rect 78680 281460 78732 281512
rect 401600 277312 401652 277364
rect 407764 277312 407816 277364
rect 425704 274660 425756 274712
rect 580172 274660 580224 274712
rect 3608 274592 3660 274644
rect 78680 274592 78732 274644
rect 401600 270444 401652 270496
rect 576124 270444 576176 270496
rect 3700 266296 3752 266348
rect 78680 266296 78732 266348
rect 407764 263576 407816 263628
rect 579804 263576 579856 263628
rect 401600 262148 401652 262200
rect 405004 262148 405056 262200
rect 3424 259360 3476 259412
rect 78680 259360 78732 259412
rect 401600 255076 401652 255128
rect 403624 255076 403676 255128
rect 403624 251200 403676 251252
rect 580172 251200 580224 251252
rect 3516 251132 3568 251184
rect 78680 251132 78732 251184
rect 3608 244196 3660 244248
rect 78680 244196 78732 244248
rect 401600 241408 401652 241460
rect 409144 241408 409196 241460
rect 3424 235900 3476 235952
rect 78680 235900 78732 235952
rect 401600 234540 401652 234592
rect 578884 234540 578936 234592
rect 3516 229032 3568 229084
rect 78680 229032 78732 229084
rect 405004 227740 405056 227792
rect 580172 227740 580224 227792
rect 401600 227672 401652 227724
rect 425704 227672 425756 227724
rect 2964 220736 3016 220788
rect 78680 220736 78732 220788
rect 401600 220736 401652 220788
rect 407764 220736 407816 220788
rect 401600 212372 401652 212424
rect 403624 212372 403676 212424
rect 3424 208292 3476 208344
rect 79324 208292 79376 208344
rect 401600 205572 401652 205624
rect 405004 205572 405056 205624
rect 401600 198636 401652 198688
rect 580264 198636 580316 198688
rect 3148 194488 3200 194540
rect 79324 194488 79376 194540
rect 401600 191768 401652 191820
rect 580356 191768 580408 191820
rect 401600 182112 401652 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 79416 180752 79468 180804
rect 402244 171028 402296 171080
rect 580172 171028 580224 171080
rect 21364 165588 21416 165640
rect 78680 165588 78732 165640
rect 3516 165520 3568 165572
rect 79324 165520 79376 165572
rect 402244 158652 402296 158704
rect 579804 158652 579856 158704
rect 3148 151716 3200 151768
rect 79508 151716 79560 151768
rect 8944 143556 8996 143608
rect 78680 143556 78732 143608
rect 3240 136552 3292 136604
rect 79416 136552 79468 136604
rect 402336 135192 402388 135244
rect 580172 135192 580224 135244
rect 401600 125604 401652 125656
rect 578884 125604 578936 125656
rect 402244 124108 402296 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 21364 122748 21416 122800
rect 21364 120096 21416 120148
rect 78680 120096 78732 120148
rect 402612 111732 402664 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 79324 108944 79376 108996
rect 401600 104864 401652 104916
rect 555424 104864 555476 104916
rect 370872 102119 370924 102128
rect 370872 102085 370881 102119
rect 370881 102085 370915 102119
rect 370915 102085 370924 102119
rect 370872 102076 370924 102085
rect 89720 100648 89772 100700
rect 90916 100648 90968 100700
rect 97172 100648 97224 100700
rect 97908 100648 97960 100700
rect 98000 100648 98052 100700
rect 99288 100648 99340 100700
rect 99656 100648 99708 100700
rect 100576 100648 100628 100700
rect 102140 100648 102192 100700
rect 103336 100648 103388 100700
rect 105360 100648 105412 100700
rect 106188 100648 106240 100700
rect 107844 100648 107896 100700
rect 108948 100648 109000 100700
rect 153200 100648 153252 100700
rect 154488 100648 154540 100700
rect 154856 100648 154908 100700
rect 155776 100648 155828 100700
rect 201868 100648 201920 100700
rect 202788 100648 202840 100700
rect 204352 100648 204404 100700
rect 205456 100648 205508 100700
rect 234896 100648 234948 100700
rect 236644 100648 236696 100700
rect 237380 100648 237432 100700
rect 238668 100648 238720 100700
rect 243084 100648 243136 100700
rect 244096 100648 244148 100700
rect 263784 100648 263836 100700
rect 264796 100648 264848 100700
rect 267832 100648 267884 100700
rect 269028 100648 269080 100700
rect 271972 100648 272024 100700
rect 273168 100648 273220 100700
rect 276112 100648 276164 100700
rect 277308 100648 277360 100700
rect 345388 100648 345440 100700
rect 346308 100648 346360 100700
rect 347872 100648 347924 100700
rect 348976 100648 349028 100700
rect 349528 100648 349580 100700
rect 350356 100648 350408 100700
rect 370136 100648 370188 100700
rect 371148 100648 371200 100700
rect 374276 100648 374328 100700
rect 375196 100648 375248 100700
rect 375932 100648 375984 100700
rect 376668 100648 376720 100700
rect 93860 100580 93912 100632
rect 97264 100580 97316 100632
rect 265348 100376 265400 100428
rect 266176 100376 266228 100428
rect 262128 100172 262180 100224
rect 291844 100172 291896 100224
rect 293408 100172 293460 100224
rect 309784 100172 309836 100224
rect 379152 100172 379204 100224
rect 403624 100172 403676 100224
rect 152372 100104 152424 100156
rect 153108 100104 153160 100156
rect 165620 100104 165672 100156
rect 174544 100104 174596 100156
rect 180432 100104 180484 100156
rect 203524 100104 203576 100156
rect 217600 100104 217652 100156
rect 224224 100104 224276 100156
rect 240692 100104 240744 100156
rect 241428 100104 241480 100156
rect 108672 100036 108724 100088
rect 135904 100036 135956 100088
rect 172244 100036 172296 100088
rect 221648 100036 221700 100088
rect 231124 100036 231176 100088
rect 238208 100036 238260 100088
rect 246304 100104 246356 100156
rect 255504 100104 255556 100156
rect 261484 100104 261536 100156
rect 280252 100104 280304 100156
rect 281356 100104 281408 100156
rect 289268 100104 289320 100156
rect 322204 100104 322256 100156
rect 335452 100104 335504 100156
rect 355324 100104 355376 100156
rect 372620 100104 372672 100156
rect 373816 100104 373868 100156
rect 392400 100104 392452 100156
rect 446404 100104 446456 100156
rect 261300 100036 261352 100088
rect 294604 100036 294656 100088
rect 331404 100036 331456 100088
rect 420184 100036 420236 100088
rect 85580 99968 85632 100020
rect 106924 99968 106976 100020
rect 133420 99968 133472 100020
rect 178684 99968 178736 100020
rect 197728 99968 197780 100020
rect 267004 99968 267056 100020
rect 271144 99968 271196 100020
rect 272524 99968 272576 100020
rect 273628 99968 273680 100020
rect 283564 99968 283616 100020
rect 292580 99968 292632 100020
rect 300124 99968 300176 100020
rect 309876 99968 309928 100020
rect 344284 99968 344336 100020
rect 384120 99968 384172 100020
rect 493324 99968 493376 100020
rect 269488 99900 269540 99952
rect 270316 99900 270368 99952
rect 376760 99832 376812 99884
rect 377956 99832 378008 99884
rect 95516 99696 95568 99748
rect 96528 99696 96580 99748
rect 149152 99696 149204 99748
rect 150348 99696 150400 99748
rect 150716 99696 150768 99748
rect 151728 99696 151780 99748
rect 200212 99696 200264 99748
rect 201408 99696 201460 99748
rect 239036 99696 239088 99748
rect 240048 99696 240100 99748
rect 281908 99696 281960 99748
rect 282828 99696 282880 99748
rect 103796 99560 103848 99612
rect 104808 99560 104860 99612
rect 306656 99492 306708 99544
rect 313924 99492 313976 99544
rect 87236 99424 87288 99476
rect 88984 99424 89036 99476
rect 130936 99424 130988 99476
rect 131764 99424 131816 99476
rect 164792 99424 164844 99476
rect 169024 99424 169076 99476
rect 183744 99424 183796 99476
rect 186964 99424 187016 99476
rect 202696 99424 202748 99476
rect 207664 99424 207716 99476
rect 241520 99424 241572 99476
rect 250444 99424 250496 99476
rect 302516 99424 302568 99476
rect 304264 99424 304316 99476
rect 311532 99424 311584 99476
rect 318064 99424 318116 99476
rect 361028 99424 361080 99476
rect 363604 99424 363656 99476
rect 364340 99424 364392 99476
rect 367744 99424 367796 99476
rect 378324 99424 378376 99476
rect 381544 99424 381596 99476
rect 383292 99424 383344 99476
rect 385684 99424 385736 99476
rect 88892 99356 88944 99408
rect 89628 99356 89680 99408
rect 109500 99356 109552 99408
rect 111064 99356 111116 99408
rect 111984 99356 112036 99408
rect 115204 99356 115256 99408
rect 116124 99356 116176 99408
rect 117228 99356 117280 99408
rect 117780 99356 117832 99408
rect 118516 99356 118568 99408
rect 120264 99356 120316 99408
rect 121276 99356 121328 99408
rect 121920 99356 121972 99408
rect 122748 99356 122800 99408
rect 124404 99356 124456 99408
rect 125508 99356 125560 99408
rect 126060 99356 126112 99408
rect 126888 99356 126940 99408
rect 128452 99356 128504 99408
rect 129648 99356 129700 99408
rect 130108 99356 130160 99408
rect 131028 99356 131080 99408
rect 132592 99356 132644 99408
rect 133788 99356 133840 99408
rect 134248 99356 134300 99408
rect 135168 99356 135220 99408
rect 136732 99356 136784 99408
rect 137928 99356 137980 99408
rect 138388 99356 138440 99408
rect 139308 99356 139360 99408
rect 140872 99356 140924 99408
rect 142068 99356 142120 99408
rect 142528 99356 142580 99408
rect 143356 99356 143408 99408
rect 145012 99356 145064 99408
rect 146116 99356 146168 99408
rect 146668 99356 146720 99408
rect 147588 99356 147640 99408
rect 157340 99356 157392 99408
rect 158536 99356 158588 99408
rect 158996 99356 159048 99408
rect 159916 99356 159968 99408
rect 160652 99356 160704 99408
rect 161388 99356 161440 99408
rect 161480 99356 161532 99408
rect 162676 99356 162728 99408
rect 163964 99356 164016 99408
rect 164884 99356 164936 99408
rect 167276 99356 167328 99408
rect 168196 99356 168248 99408
rect 168932 99356 168984 99408
rect 169668 99356 169720 99408
rect 169760 99356 169812 99408
rect 170956 99356 171008 99408
rect 171416 99356 171468 99408
rect 172428 99356 172480 99408
rect 173072 99356 173124 99408
rect 173808 99356 173860 99408
rect 175464 99356 175516 99408
rect 176568 99356 176620 99408
rect 179604 99356 179656 99408
rect 180708 99356 180760 99408
rect 181260 99356 181312 99408
rect 182824 99356 182876 99408
rect 185400 99356 185452 99408
rect 186228 99356 186280 99408
rect 187884 99356 187936 99408
rect 188988 99356 189040 99408
rect 189540 99356 189592 99408
rect 191104 99356 191156 99408
rect 192024 99356 192076 99408
rect 193036 99356 193088 99408
rect 206008 99356 206060 99408
rect 206836 99356 206888 99408
rect 208492 99356 208544 99408
rect 209596 99356 209648 99408
rect 210148 99356 210200 99408
rect 210976 99356 211028 99408
rect 212632 99356 212684 99408
rect 213828 99356 213880 99408
rect 214288 99356 214340 99408
rect 215944 99356 215996 99408
rect 216772 99356 216824 99408
rect 217968 99356 218020 99408
rect 218428 99356 218480 99408
rect 219256 99356 219308 99408
rect 220820 99356 220872 99408
rect 222108 99356 222160 99408
rect 222476 99356 222528 99408
rect 223396 99356 223448 99408
rect 224132 99356 224184 99408
rect 224868 99356 224920 99408
rect 224960 99356 225012 99408
rect 226248 99356 226300 99408
rect 226616 99356 226668 99408
rect 227628 99356 227680 99408
rect 229100 99356 229152 99408
rect 230296 99356 230348 99408
rect 232412 99356 232464 99408
rect 233148 99356 233200 99408
rect 233240 99356 233292 99408
rect 234436 99356 234488 99408
rect 244740 99356 244792 99408
rect 245568 99356 245620 99408
rect 247224 99356 247276 99408
rect 248236 99356 248288 99408
rect 251364 99356 251416 99408
rect 252468 99356 252520 99408
rect 253020 99356 253072 99408
rect 254584 99356 254636 99408
rect 259644 99356 259696 99408
rect 260748 99356 260800 99408
rect 284392 99356 284444 99408
rect 285588 99356 285640 99408
rect 286048 99356 286100 99408
rect 286876 99356 286928 99408
rect 287612 99356 287664 99408
rect 288348 99356 288400 99408
rect 288440 99356 288492 99408
rect 289728 99356 289780 99408
rect 290096 99356 290148 99408
rect 291016 99356 291068 99408
rect 294236 99356 294288 99408
rect 295248 99356 295300 99408
rect 295892 99356 295944 99408
rect 296628 99356 296680 99408
rect 296720 99356 296772 99408
rect 297916 99356 297968 99408
rect 298376 99356 298428 99408
rect 299296 99356 299348 99408
rect 300860 99356 300912 99408
rect 302056 99356 302108 99408
rect 304172 99356 304224 99408
rect 304908 99356 304960 99408
rect 309140 99356 309192 99408
rect 310428 99356 310480 99408
rect 310704 99356 310756 99408
rect 311808 99356 311860 99408
rect 314844 99356 314896 99408
rect 315856 99356 315908 99408
rect 316500 99356 316552 99408
rect 317236 99356 317288 99408
rect 318984 99356 319036 99408
rect 319996 99356 320048 99408
rect 320640 99356 320692 99408
rect 321468 99356 321520 99408
rect 323124 99356 323176 99408
rect 324228 99356 324280 99408
rect 324780 99356 324832 99408
rect 326344 99356 326396 99408
rect 327264 99356 327316 99408
rect 328276 99356 328328 99408
rect 328920 99356 328972 99408
rect 331864 99356 331916 99408
rect 332968 99356 333020 99408
rect 333796 99356 333848 99408
rect 337108 99356 337160 99408
rect 337936 99356 337988 99408
rect 339592 99356 339644 99408
rect 340788 99356 340840 99408
rect 352012 99356 352064 99408
rect 353116 99356 353168 99408
rect 353668 99356 353720 99408
rect 354496 99356 354548 99408
rect 356060 99356 356112 99408
rect 357256 99356 357308 99408
rect 357716 99356 357768 99408
rect 358728 99356 358780 99408
rect 359372 99356 359424 99408
rect 360108 99356 360160 99408
rect 360200 99356 360252 99408
rect 361488 99356 361540 99408
rect 361856 99356 361908 99408
rect 362776 99356 362828 99408
rect 365996 99356 366048 99408
rect 366916 99356 366968 99408
rect 367652 99356 367704 99408
rect 368388 99356 368440 99408
rect 368480 99356 368532 99408
rect 369676 99356 369728 99408
rect 379980 99356 380032 99408
rect 380716 99356 380768 99408
rect 382464 99356 382516 99408
rect 383568 99356 383620 99408
rect 386604 99356 386656 99408
rect 387616 99356 387668 99408
rect 388260 99356 388312 99408
rect 388996 99356 389048 99408
rect 390744 99356 390796 99408
rect 391756 99356 391808 99408
rect 396540 99356 396592 99408
rect 398104 99356 398156 99408
rect 399024 99356 399076 99408
rect 400128 99356 400180 99408
rect 370872 99331 370924 99340
rect 370872 99297 370881 99331
rect 370881 99297 370915 99331
rect 370915 99297 370924 99331
rect 370872 99288 370924 99297
rect 228272 98744 228324 98796
rect 333980 98744 334032 98796
rect 317328 98676 317380 98728
rect 462320 98676 462372 98728
rect 91376 98608 91428 98660
rect 92388 98608 92440 98660
rect 145840 98608 145892 98660
rect 215300 98608 215352 98660
rect 333704 98608 333756 98660
rect 485780 98608 485832 98660
rect 342076 98583 342128 98592
rect 342076 98549 342085 98583
rect 342085 98549 342119 98583
rect 342119 98549 342128 98583
rect 342076 98540 342128 98549
rect 163136 97316 163188 97368
rect 240140 97316 240192 97368
rect 312360 97316 312412 97368
rect 455420 97316 455472 97368
rect 230756 97248 230808 97300
rect 338120 97248 338172 97300
rect 341248 97248 341300 97300
rect 496820 97248 496872 97300
rect 278504 96704 278556 96756
rect 278688 96704 278740 96756
rect 267004 96611 267056 96620
rect 267004 96577 267013 96611
rect 267013 96577 267047 96611
rect 267047 96577 267056 96611
rect 267004 96568 267056 96577
rect 278688 96568 278740 96620
rect 305000 95956 305052 96008
rect 444380 95956 444432 96008
rect 149980 95888 150032 95940
rect 220820 95888 220872 95940
rect 225788 95888 225840 95940
rect 331220 95888 331272 95940
rect 343732 95888 343784 95940
rect 500960 95888 501012 95940
rect 92112 95276 92164 95328
rect 92296 95208 92348 95260
rect 198004 95251 198056 95260
rect 198004 95217 198013 95251
rect 198013 95217 198047 95251
rect 198047 95217 198056 95251
rect 198004 95208 198056 95217
rect 198004 95115 198056 95124
rect 198004 95081 198013 95115
rect 198013 95081 198047 95115
rect 198047 95081 198056 95115
rect 198004 95072 198056 95081
rect 277768 94596 277820 94648
rect 405740 94596 405792 94648
rect 346216 94528 346268 94580
rect 503720 94528 503772 94580
rect 196072 94460 196124 94512
rect 287060 94460 287112 94512
rect 394884 94460 394936 94512
rect 574100 94460 574152 94512
rect 3424 93780 3476 93832
rect 79692 93780 79744 93832
rect 295064 93168 295116 93220
rect 430580 93168 430632 93220
rect 147496 93100 147548 93152
rect 218060 93100 218112 93152
rect 219256 93100 219308 93152
rect 320180 93100 320232 93152
rect 354496 93100 354548 93152
rect 514760 93100 514812 93152
rect 153108 91808 153160 91860
rect 224960 91808 225012 91860
rect 291016 91808 291068 91860
rect 423680 91808 423732 91860
rect 216588 91740 216640 91792
rect 316040 91740 316092 91792
rect 357256 91740 357308 91792
rect 518900 91740 518952 91792
rect 155776 90380 155828 90432
rect 227720 90380 227772 90432
rect 285496 90380 285548 90432
rect 416780 90380 416832 90432
rect 213736 90312 213788 90364
rect 313280 90312 313332 90364
rect 358544 90312 358596 90364
rect 521660 90312 521712 90364
rect 92204 89743 92256 89752
rect 92204 89709 92213 89743
rect 92213 89709 92247 89743
rect 92247 89709 92256 89743
rect 92204 89700 92256 89709
rect 151452 89700 151504 89752
rect 151636 89700 151688 89752
rect 198556 89743 198608 89752
rect 198556 89709 198565 89743
rect 198565 89709 198599 89743
rect 198599 89709 198608 89743
rect 198556 89700 198608 89709
rect 227444 89743 227496 89752
rect 227444 89709 227453 89743
rect 227453 89709 227487 89743
rect 227487 89709 227496 89743
rect 227444 89700 227496 89709
rect 274364 89700 274416 89752
rect 274548 89700 274600 89752
rect 267004 89675 267056 89684
rect 267004 89641 267013 89675
rect 267013 89641 267047 89675
rect 267047 89641 267056 89675
rect 267004 89632 267056 89641
rect 282736 89088 282788 89140
rect 412640 89088 412692 89140
rect 158536 89020 158588 89072
rect 231860 89020 231912 89072
rect 299296 89020 299348 89072
rect 434720 89020 434772 89072
rect 210976 88952 211028 89004
rect 307760 88952 307812 89004
rect 364248 88952 364300 89004
rect 528560 88952 528612 89004
rect 402520 88272 402572 88324
rect 580172 88272 580224 88324
rect 146116 87660 146168 87712
rect 213920 87660 213972 87712
rect 264796 87660 264848 87712
rect 385040 87660 385092 87712
rect 187608 87592 187660 87644
rect 274640 87592 274692 87644
rect 277216 87592 277268 87644
rect 404360 87592 404412 87644
rect 104624 86980 104676 87032
rect 104716 86980 104768 87032
rect 227444 87023 227496 87032
rect 227444 86989 227453 87023
rect 227453 86989 227487 87023
rect 227487 86989 227496 87023
rect 227444 86980 227496 86989
rect 239864 86980 239916 87032
rect 239956 86980 240008 87032
rect 278596 87023 278648 87032
rect 278596 86989 278605 87023
rect 278605 86989 278639 87023
rect 278639 86989 278648 87023
rect 278596 86980 278648 86989
rect 342076 87023 342128 87032
rect 342076 86989 342085 87023
rect 342085 86989 342119 87023
rect 342119 86989 342128 87023
rect 342076 86980 342128 86989
rect 309784 86368 309836 86420
rect 427820 86368 427872 86420
rect 281356 86300 281408 86352
rect 408500 86300 408552 86352
rect 143356 86232 143408 86284
rect 209780 86232 209832 86284
rect 211068 86232 211120 86284
rect 309140 86232 309192 86284
rect 366916 86232 366968 86284
rect 532700 86232 532752 86284
rect 92204 85595 92256 85604
rect 92204 85561 92213 85595
rect 92213 85561 92247 85595
rect 92247 85561 92256 85595
rect 92204 85552 92256 85561
rect 96344 85552 96396 85604
rect 96436 85552 96488 85604
rect 198096 85552 198148 85604
rect 198556 85595 198608 85604
rect 198556 85561 198565 85595
rect 198565 85561 198599 85595
rect 198599 85561 198608 85595
rect 198556 85552 198608 85561
rect 518900 85527 518952 85536
rect 518900 85493 518909 85527
rect 518909 85493 518943 85527
rect 518943 85493 518952 85527
rect 518900 85484 518952 85493
rect 532700 85527 532752 85536
rect 532700 85493 532709 85527
rect 532709 85493 532743 85527
rect 532743 85493 532752 85527
rect 532700 85484 532752 85493
rect 275928 84940 275980 84992
rect 401600 84940 401652 84992
rect 289728 84872 289780 84924
rect 420920 84872 420972 84924
rect 209596 84804 209648 84856
rect 305000 84804 305052 84856
rect 369676 84804 369728 84856
rect 536840 84804 536892 84856
rect 273076 83512 273128 83564
rect 398840 83512 398892 83564
rect 400036 83512 400088 83564
rect 482284 83512 482336 83564
rect 206836 83444 206888 83496
rect 302240 83444 302292 83496
rect 370688 83444 370740 83496
rect 539600 83444 539652 83496
rect 140688 82152 140740 82204
rect 207020 82152 207072 82204
rect 315856 82152 315908 82204
rect 459652 82152 459704 82204
rect 104624 82127 104676 82136
rect 104624 82093 104633 82127
rect 104633 82093 104667 82127
rect 104667 82093 104676 82127
rect 104624 82084 104676 82093
rect 175188 82084 175240 82136
rect 256700 82084 256752 82136
rect 257896 82084 257948 82136
rect 375380 82084 375432 82136
rect 381544 82084 381596 82136
rect 550640 82084 550692 82136
rect 227076 82016 227128 82068
rect 227444 82016 227496 82068
rect 341708 82016 341760 82068
rect 342076 82016 342128 82068
rect 239864 81855 239916 81864
rect 239864 81821 239873 81855
rect 239873 81821 239907 81855
rect 239907 81821 239916 81855
rect 239864 81812 239916 81821
rect 266176 80792 266228 80844
rect 387800 80792 387852 80844
rect 91928 80724 91980 80776
rect 277308 80724 277360 80776
rect 402980 80724 403032 80776
rect 137836 80656 137888 80708
rect 202880 80656 202932 80708
rect 204168 80656 204220 80708
rect 298100 80656 298152 80708
rect 385684 80656 385736 80708
rect 557540 80656 557592 80708
rect 198096 80180 198148 80232
rect 267096 80155 267148 80164
rect 267096 80121 267105 80155
rect 267105 80121 267139 80155
rect 267139 80121 267148 80155
rect 267096 80112 267148 80121
rect 278596 80044 278648 80096
rect 278688 79908 278740 79960
rect 3516 79432 3568 79484
rect 8944 79432 8996 79484
rect 201316 79364 201368 79416
rect 295340 79364 295392 79416
rect 329748 79364 329800 79416
rect 480260 79364 480312 79416
rect 135076 79296 135128 79348
rect 200120 79296 200172 79348
rect 263508 79296 263560 79348
rect 383660 79296 383712 79348
rect 388996 79296 389048 79348
rect 564440 79296 564492 79348
rect 198556 78004 198608 78056
rect 291200 78004 291252 78056
rect 307668 78004 307720 78056
rect 448520 78004 448572 78056
rect 133788 77936 133840 77988
rect 195980 77936 196032 77988
rect 260656 77936 260708 77988
rect 380900 77936 380952 77988
rect 391756 77936 391808 77988
rect 568580 77936 568632 77988
rect 104624 77367 104676 77376
rect 104624 77333 104633 77367
rect 104633 77333 104667 77367
rect 104667 77333 104676 77367
rect 104624 77324 104676 77333
rect 239864 77367 239916 77376
rect 239864 77333 239873 77367
rect 239873 77333 239907 77367
rect 239907 77333 239916 77367
rect 239864 77324 239916 77333
rect 267096 77299 267148 77308
rect 267096 77265 267105 77299
rect 267105 77265 267139 77299
rect 267139 77265 267148 77299
rect 267096 77256 267148 77265
rect 104532 77231 104584 77240
rect 104532 77197 104541 77231
rect 104541 77197 104575 77231
rect 104575 77197 104584 77231
rect 104532 77188 104584 77197
rect 151544 77231 151596 77240
rect 151544 77197 151553 77231
rect 151553 77197 151587 77231
rect 151587 77197 151596 77231
rect 151544 77188 151596 77197
rect 239772 77231 239824 77240
rect 239772 77197 239781 77231
rect 239781 77197 239815 77231
rect 239815 77197 239824 77231
rect 239772 77188 239824 77197
rect 402428 77188 402480 77240
rect 580172 77188 580224 77240
rect 254584 76576 254636 76628
rect 369860 76576 369912 76628
rect 131028 76508 131080 76560
rect 193220 76508 193272 76560
rect 194416 76508 194468 76560
rect 284300 76508 284352 76560
rect 304264 76508 304316 76560
rect 441620 76508 441672 76560
rect 198004 75939 198056 75948
rect 198004 75905 198013 75939
rect 198013 75905 198047 75939
rect 198047 75905 198056 75939
rect 198004 75896 198056 75905
rect 518900 75939 518952 75948
rect 518900 75905 518909 75939
rect 518909 75905 518943 75939
rect 518943 75905 518952 75939
rect 518900 75896 518952 75905
rect 532700 75939 532752 75948
rect 532700 75905 532709 75939
rect 532709 75905 532743 75939
rect 532743 75905 532752 75939
rect 532700 75896 532752 75905
rect 191748 75216 191800 75268
rect 280160 75216 280212 75268
rect 300768 75216 300820 75268
rect 437480 75216 437532 75268
rect 128268 75148 128320 75200
rect 189080 75148 189132 75200
rect 245476 75148 245528 75200
rect 358820 75148 358872 75200
rect 393228 75148 393280 75200
rect 571340 75148 571392 75200
rect 215024 74468 215076 74520
rect 215208 74468 215260 74520
rect 188896 73856 188948 73908
rect 277400 73856 277452 73908
rect 300124 73856 300176 73908
rect 426440 73856 426492 73908
rect 244096 73788 244148 73840
rect 356060 73788 356112 73840
rect 395988 73788 396040 73840
rect 575480 73788 575532 73840
rect 186136 72496 186188 72548
rect 273260 72496 273312 72548
rect 282828 72496 282880 72548
rect 411260 72496 411312 72548
rect 224868 72428 224920 72480
rect 328460 72428 328512 72480
rect 375196 72428 375248 72480
rect 545120 72428 545172 72480
rect 274548 71179 274600 71188
rect 274548 71145 274557 71179
rect 274557 71145 274591 71179
rect 274591 71145 274600 71179
rect 274548 71136 274600 71145
rect 285588 71136 285640 71188
rect 415400 71136 415452 71188
rect 186964 71068 187016 71120
rect 270500 71068 270552 71120
rect 303528 71068 303580 71120
rect 443000 71068 443052 71120
rect 125416 71000 125468 71052
rect 184940 71000 184992 71052
rect 219348 71000 219400 71052
rect 321560 71000 321612 71052
rect 377956 71000 378008 71052
rect 547880 71000 547932 71052
rect 227352 70456 227404 70508
rect 267096 70431 267148 70440
rect 267096 70397 267105 70431
rect 267105 70397 267139 70431
rect 267139 70397 267148 70431
rect 267096 70388 267148 70397
rect 341984 70456 342036 70508
rect 227260 70320 227312 70372
rect 341892 70320 341944 70372
rect 182824 69776 182876 69828
rect 266360 69776 266412 69828
rect 209688 69708 209740 69760
rect 306380 69708 306432 69760
rect 322204 69708 322256 69760
rect 422300 69708 422352 69760
rect 122656 69640 122708 69692
rect 182180 69640 182232 69692
rect 256608 69640 256660 69692
rect 374000 69640 374052 69692
rect 382188 69640 382240 69692
rect 554780 69640 554832 69692
rect 292488 68416 292540 68468
rect 425060 68416 425112 68468
rect 179328 68348 179380 68400
rect 262220 68348 262272 68400
rect 302056 68348 302108 68400
rect 438860 68348 438912 68400
rect 121276 68280 121328 68332
rect 178040 68280 178092 68332
rect 215944 68280 215996 68332
rect 313372 68280 313424 68332
rect 387616 68280 387668 68332
rect 563060 68280 563112 68332
rect 92296 67600 92348 67652
rect 104624 67600 104676 67652
rect 151636 67600 151688 67652
rect 239864 67600 239916 67652
rect 267096 67643 267148 67652
rect 267096 67609 267105 67643
rect 267105 67609 267139 67643
rect 267139 67609 267148 67643
rect 267096 67600 267148 67609
rect 274548 67643 274600 67652
rect 274548 67609 274557 67643
rect 274557 67609 274591 67643
rect 274591 67609 274600 67643
rect 274548 67600 274600 67609
rect 550640 67600 550692 67652
rect 550916 67600 550968 67652
rect 151452 67464 151504 67516
rect 151636 67464 151688 67516
rect 274364 67464 274416 67516
rect 274548 67464 274600 67516
rect 278596 66988 278648 67040
rect 407120 66988 407172 67040
rect 176476 66920 176528 66972
rect 259460 66920 259512 66972
rect 295248 66920 295300 66972
rect 429200 66920 429252 66972
rect 118516 66852 118568 66904
rect 175280 66852 175332 66904
rect 212448 66852 212500 66904
rect 310520 66852 310572 66904
rect 389088 66852 389140 66904
rect 565820 66852 565872 66904
rect 96344 66172 96396 66224
rect 200120 66215 200172 66224
rect 200120 66181 200129 66215
rect 200129 66181 200163 66215
rect 200163 66181 200172 66215
rect 200120 66172 200172 66181
rect 227260 66172 227312 66224
rect 227444 66172 227496 66224
rect 341892 66215 341944 66224
rect 341892 66181 341901 66215
rect 341901 66181 341935 66215
rect 341935 66181 341944 66215
rect 341892 66172 341944 66181
rect 518900 66215 518952 66224
rect 518900 66181 518909 66215
rect 518909 66181 518943 66215
rect 518943 66181 518952 66215
rect 518900 66172 518952 66181
rect 532700 66215 532752 66224
rect 532700 66181 532709 66215
rect 532709 66181 532743 66215
rect 532743 66181 532752 66215
rect 532700 66172 532752 66181
rect 268936 65628 268988 65680
rect 391940 65628 391992 65680
rect 173716 65560 173768 65612
rect 255320 65560 255372 65612
rect 297916 65560 297968 65612
rect 433340 65560 433392 65612
rect 206928 65492 206980 65544
rect 303620 65492 303672 65544
rect 391848 65492 391900 65544
rect 3332 64812 3384 64864
rect 79600 64812 79652 64864
rect 205456 64200 205508 64252
rect 299480 64200 299532 64252
rect 302148 64200 302200 64252
rect 440240 64200 440292 64252
rect 115848 64132 115900 64184
rect 171140 64132 171192 64184
rect 172428 64132 172480 64184
rect 252560 64132 252612 64184
rect 253848 64132 253900 64184
rect 371240 64132 371292 64184
rect 398104 64132 398156 64184
rect 576860 64132 576912 64184
rect 214932 63452 214984 63504
rect 215024 63452 215076 63504
rect 239864 62951 239916 62960
rect 239864 62917 239873 62951
rect 239873 62917 239907 62951
rect 239907 62917 239916 62951
rect 239864 62908 239916 62917
rect 202788 62840 202840 62892
rect 296720 62840 296772 62892
rect 313924 62840 313976 62892
rect 447140 62840 447192 62892
rect 113088 62772 113140 62824
rect 167000 62772 167052 62824
rect 169668 62772 169720 62824
rect 248420 62772 248472 62824
rect 250444 62772 250496 62824
rect 353300 62772 353352 62824
rect 400128 62772 400180 62824
rect 578884 62772 578936 62824
rect 267096 62747 267148 62756
rect 267096 62713 267105 62747
rect 267105 62713 267139 62747
rect 267139 62713 267148 62747
rect 267096 62704 267148 62713
rect 166908 61412 166960 61464
rect 244280 61412 244332 61464
rect 310428 61412 310480 61464
rect 451280 61412 451332 61464
rect 110328 61344 110380 61396
rect 164240 61344 164292 61396
rect 200028 61344 200080 61396
rect 292580 61344 292632 61396
rect 322848 61344 322900 61396
rect 469220 61344 469272 61396
rect 104624 60800 104676 60852
rect 104532 60664 104584 60716
rect 235908 60052 235960 60104
rect 345020 60052 345072 60104
rect 355324 60052 355376 60104
rect 488540 60052 488592 60104
rect 162676 59984 162728 60036
rect 237380 59984 237432 60036
rect 317236 59984 317288 60036
rect 460940 59984 460992 60036
rect 234436 58760 234488 58812
rect 340880 58760 340932 58812
rect 319996 58692 320048 58744
rect 465080 58692 465132 58744
rect 107568 58624 107620 58676
rect 158720 58624 158772 58676
rect 159916 58624 159968 58676
rect 234620 58624 234672 58676
rect 340696 58624 340748 58676
rect 495440 58624 495492 58676
rect 197728 57944 197780 57996
rect 198004 57944 198056 57996
rect 239680 57944 239732 57996
rect 267096 57987 267148 57996
rect 267096 57953 267105 57987
rect 267105 57953 267139 57987
rect 267139 57953 267148 57987
rect 267096 57944 267148 57953
rect 92204 57876 92256 57928
rect 286876 57332 286928 57384
rect 416872 57332 416924 57384
rect 193036 57264 193088 57316
rect 281540 57264 281592 57316
rect 299388 57264 299440 57316
rect 436100 57264 436152 57316
rect 104532 57196 104584 57248
rect 155960 57196 156012 57248
rect 157248 57196 157300 57248
rect 230480 57196 230532 57248
rect 231124 57196 231176 57248
rect 324320 57196 324372 57248
rect 394608 57196 394660 57248
rect 572720 57196 572772 57248
rect 96252 56627 96304 56636
rect 96252 56593 96261 56627
rect 96261 56593 96295 56627
rect 96295 56593 96304 56627
rect 96252 56584 96304 56593
rect 200120 56627 200172 56636
rect 200120 56593 200129 56627
rect 200129 56593 200163 56627
rect 200163 56593 200172 56627
rect 200120 56584 200172 56593
rect 342076 56584 342128 56636
rect 518900 56627 518952 56636
rect 518900 56593 518909 56627
rect 518909 56593 518943 56627
rect 518943 56593 518952 56627
rect 518900 56584 518952 56593
rect 532700 56627 532752 56636
rect 532700 56593 532709 56627
rect 532709 56593 532743 56627
rect 532743 56593 532752 56627
rect 532700 56584 532752 56593
rect 569960 56627 570012 56636
rect 569960 56593 569969 56627
rect 569969 56593 570003 56627
rect 570003 56593 570012 56627
rect 569960 56584 570012 56593
rect 96252 56491 96304 56500
rect 96252 56457 96261 56491
rect 96261 56457 96295 56491
rect 96295 56457 96304 56491
rect 96252 56448 96304 56457
rect 286968 55972 287020 56024
rect 418160 55972 418212 56024
rect 191104 55904 191156 55956
rect 278780 55904 278832 55956
rect 296628 55904 296680 55956
rect 431960 55904 432012 55956
rect 103336 55836 103388 55888
rect 151820 55836 151872 55888
rect 154396 55836 154448 55888
rect 227812 55836 227864 55888
rect 230296 55836 230348 55888
rect 335360 55836 335412 55888
rect 403624 55836 403676 55888
rect 552020 55836 552072 55888
rect 274364 54612 274416 54664
rect 400220 54612 400272 54664
rect 151452 54544 151504 54596
rect 223580 54544 223632 54596
rect 281448 54544 281500 54596
rect 409880 54544 409932 54596
rect 194508 54476 194560 54528
rect 285680 54476 285732 54528
rect 369768 54476 369820 54528
rect 536932 54476 536984 54528
rect 182088 53116 182140 53168
rect 273168 53116 273220 53168
rect 397460 53116 397512 53168
rect 100576 53048 100628 53100
rect 149060 53048 149112 53100
rect 150348 53048 150400 53100
rect 219440 53048 219492 53100
rect 249616 53048 249668 53100
rect 364340 53048 364392 53100
rect 367008 53048 367060 53100
rect 534080 53048 534132 53100
rect 180708 51756 180760 51808
rect 263600 51756 263652 51808
rect 270316 51756 270368 51808
rect 393320 51756 393372 51808
rect 97908 51688 97960 51740
rect 144920 51688 144972 51740
rect 147588 51688 147640 51740
rect 216680 51688 216732 51740
rect 246948 51688 247000 51740
rect 360200 51688 360252 51740
rect 367744 51688 367796 51740
rect 529940 51688 529992 51740
rect 239680 51119 239732 51128
rect 239680 51085 239689 51119
rect 239689 51085 239723 51119
rect 239723 51085 239732 51119
rect 239680 51076 239732 51085
rect 267096 51119 267148 51128
rect 267096 51085 267105 51119
rect 267105 51085 267139 51119
rect 267139 51085 267148 51119
rect 267096 51076 267148 51085
rect 342076 51076 342128 51128
rect 3424 51008 3476 51060
rect 79508 51008 79560 51060
rect 342076 50940 342128 50992
rect 144828 50396 144880 50448
rect 212540 50396 212592 50448
rect 231768 50396 231820 50448
rect 339500 50396 339552 50448
rect 362776 50396 362828 50448
rect 527180 50396 527232 50448
rect 177856 50328 177908 50380
rect 260840 50328 260892 50380
rect 267648 50328 267700 50380
rect 390560 50328 390612 50380
rect 397368 50328 397420 50380
rect 567936 50328 567988 50380
rect 197268 49036 197320 49088
rect 288440 49036 288492 49088
rect 353116 49036 353168 49088
rect 512000 49036 512052 49088
rect 95148 48968 95200 49020
rect 140780 48968 140832 49020
rect 141976 48968 142028 49020
rect 209872 48968 209924 49020
rect 252376 48968 252428 49020
rect 368480 48968 368532 49020
rect 378048 48968 378100 49020
rect 549260 48968 549312 49020
rect 92112 48331 92164 48340
rect 92112 48297 92121 48331
rect 92121 48297 92155 48331
rect 92155 48297 92164 48331
rect 92112 48288 92164 48297
rect 239680 48331 239732 48340
rect 239680 48297 239689 48331
rect 239689 48297 239723 48331
rect 239723 48297 239732 48331
rect 239680 48288 239732 48297
rect 267096 48331 267148 48340
rect 267096 48297 267105 48331
rect 267105 48297 267139 48331
rect 267139 48297 267148 48331
rect 267096 48288 267148 48297
rect 567936 48220 567988 48272
rect 170956 47608 171008 47660
rect 249800 47608 249852 47660
rect 350356 47608 350408 47660
rect 509240 47608 509292 47660
rect 92112 47540 92164 47592
rect 138020 47540 138072 47592
rect 139216 47540 139268 47592
rect 205640 47540 205692 47592
rect 249708 47540 249760 47592
rect 365720 47540 365772 47592
rect 373816 47540 373868 47592
rect 542360 47540 542412 47592
rect 96344 46928 96396 46980
rect 267740 46971 267792 46980
rect 267740 46937 267749 46971
rect 267749 46937 267783 46971
rect 267783 46937 267792 46971
rect 267740 46928 267792 46937
rect 138020 46903 138072 46912
rect 138020 46869 138029 46903
rect 138029 46869 138063 46903
rect 138063 46869 138072 46903
rect 138020 46860 138072 46869
rect 200120 46903 200172 46912
rect 200120 46869 200129 46903
rect 200129 46869 200163 46903
rect 200163 46869 200172 46903
rect 200120 46860 200172 46869
rect 509240 46903 509292 46912
rect 509240 46869 509249 46903
rect 509249 46869 509283 46903
rect 509283 46869 509292 46903
rect 509240 46860 509292 46869
rect 518900 46903 518952 46912
rect 518900 46869 518909 46903
rect 518909 46869 518943 46903
rect 518943 46869 518952 46903
rect 518900 46860 518952 46869
rect 527180 46903 527232 46912
rect 527180 46869 527189 46903
rect 527189 46869 527223 46903
rect 527223 46869 527232 46903
rect 527180 46860 527232 46869
rect 532700 46903 532752 46912
rect 532700 46869 532709 46903
rect 532709 46869 532743 46903
rect 532743 46869 532752 46903
rect 532700 46860 532752 46869
rect 569960 46903 570012 46912
rect 569960 46869 569969 46903
rect 569969 46869 570003 46903
rect 570003 46869 570012 46903
rect 569960 46860 570012 46869
rect 137928 46248 137980 46300
rect 201500 46248 201552 46300
rect 347688 46248 347740 46300
rect 505100 46248 505152 46300
rect 169024 46180 169076 46232
rect 242900 46180 242952 46232
rect 245568 46180 245620 46232
rect 357440 46180 357492 46232
rect 371148 46180 371200 46232
rect 538220 46180 538272 46232
rect 114376 44888 114428 44940
rect 168380 44888 168432 44940
rect 344928 44888 344980 44940
rect 502340 44888 502392 44940
rect 164884 44820 164936 44872
rect 241520 44820 241572 44872
rect 242808 44820 242860 44872
rect 354680 44820 354732 44872
rect 368388 44820 368440 44872
rect 535460 44820 535512 44872
rect 168196 43460 168248 43512
rect 245660 43460 245712 43512
rect 342076 43460 342128 43512
rect 498200 43460 498252 43512
rect 135168 43392 135220 43444
rect 198740 43392 198792 43444
rect 239680 43392 239732 43444
rect 350540 43392 350592 43444
rect 365628 43392 365680 43444
rect 531320 43392 531372 43444
rect 132408 42100 132460 42152
rect 194600 42100 194652 42152
rect 340788 42100 340840 42152
rect 494060 42100 494112 42152
rect 160008 42032 160060 42084
rect 236000 42032 236052 42084
rect 238668 42032 238720 42084
rect 347780 42032 347832 42084
rect 355968 42032 356020 42084
rect 517520 42032 517572 42084
rect 267096 41488 267148 41540
rect 96344 41420 96396 41472
rect 214932 41420 214984 41472
rect 227260 41420 227312 41472
rect 96252 41352 96304 41404
rect 215024 41284 215076 41336
rect 402336 41352 402388 41404
rect 580172 41352 580224 41404
rect 227352 41284 227404 41336
rect 226248 40808 226300 40860
rect 329840 40808 329892 40860
rect 270408 40740 270460 40792
rect 394700 40740 394752 40792
rect 129556 40672 129608 40724
rect 191840 40672 191892 40724
rect 284208 40672 284260 40724
rect 414020 40672 414072 40724
rect 184848 39380 184900 39432
rect 270592 39380 270644 39432
rect 326988 39380 327040 39432
rect 476120 39380 476172 39432
rect 126796 39312 126848 39364
rect 187700 39312 187752 39364
rect 223396 39312 223448 39364
rect 325700 39312 325752 39364
rect 346308 39312 346360 39364
rect 502432 39312 502484 39364
rect 267004 38675 267056 38684
rect 267004 38641 267013 38675
rect 267013 38641 267047 38675
rect 267047 38641 267056 38675
rect 267004 38632 267056 38641
rect 567844 38675 567896 38684
rect 567844 38641 567853 38675
rect 567853 38641 567887 38675
rect 567887 38641 567896 38675
rect 567844 38632 567896 38641
rect 198556 38564 198608 38616
rect 198740 38564 198792 38616
rect 162768 38020 162820 38072
rect 238760 38020 238812 38072
rect 220728 37952 220780 38004
rect 321652 37952 321704 38004
rect 331864 37952 331916 38004
rect 478880 37952 478932 38004
rect 122748 37884 122800 37936
rect 180800 37884 180852 37936
rect 237288 37884 237340 37936
rect 346400 37884 346452 37936
rect 348976 37884 349028 37936
rect 506480 37884 506532 37936
rect 138020 37315 138072 37324
rect 138020 37281 138029 37315
rect 138029 37281 138063 37315
rect 138063 37281 138072 37315
rect 138020 37272 138072 37281
rect 200120 37315 200172 37324
rect 200120 37281 200129 37315
rect 200129 37281 200163 37315
rect 200163 37281 200172 37315
rect 200120 37272 200172 37281
rect 509240 37315 509292 37324
rect 509240 37281 509249 37315
rect 509249 37281 509283 37315
rect 509283 37281 509292 37315
rect 509240 37272 509292 37281
rect 518900 37315 518952 37324
rect 518900 37281 518909 37315
rect 518909 37281 518943 37315
rect 518943 37281 518952 37315
rect 518900 37272 518952 37281
rect 527180 37315 527232 37324
rect 527180 37281 527189 37315
rect 527189 37281 527223 37315
rect 527223 37281 527232 37315
rect 527180 37272 527232 37281
rect 532700 37315 532752 37324
rect 532700 37281 532709 37315
rect 532709 37281 532743 37315
rect 532743 37281 532752 37315
rect 532700 37272 532752 37281
rect 569960 37315 570012 37324
rect 569960 37281 569969 37315
rect 569969 37281 570003 37315
rect 570003 37281 570012 37315
rect 569960 37272 570012 37281
rect 215024 37247 215076 37256
rect 215024 37213 215033 37247
rect 215033 37213 215067 37247
rect 215067 37213 215076 37247
rect 215024 37204 215076 37213
rect 227352 37247 227404 37256
rect 227352 37213 227361 37247
rect 227361 37213 227395 37247
rect 227395 37213 227404 37247
rect 227352 37204 227404 37213
rect 314568 36592 314620 36644
rect 458180 36592 458232 36644
rect 119988 36524 120040 36576
rect 176660 36524 176712 36576
rect 213828 36524 213880 36576
rect 311900 36524 311952 36576
rect 328276 36524 328328 36576
rect 477592 36524 477644 36576
rect 3424 35844 3476 35896
rect 21364 35844 21416 35896
rect 190368 35232 190420 35284
rect 278872 35232 278924 35284
rect 280068 35232 280120 35284
rect 408592 35232 408644 35284
rect 117136 35164 117188 35216
rect 173900 35164 173952 35216
rect 252468 35164 252520 35216
rect 367100 35164 367152 35216
rect 372528 35164 372580 35216
rect 540980 35164 541032 35216
rect 360108 33804 360160 33856
rect 523040 33804 523092 33856
rect 114468 33736 114520 33788
rect 169760 33736 169812 33788
rect 177948 33736 178000 33788
rect 262312 33736 262364 33788
rect 264888 33736 264940 33788
rect 386420 33736 386472 33788
rect 387708 33736 387760 33788
rect 563152 33736 563204 33788
rect 357348 32444 357400 32496
rect 520280 32444 520332 32496
rect 115204 32376 115256 32428
rect 167092 32376 167144 32428
rect 176568 32376 176620 32428
rect 258080 32376 258132 32428
rect 260748 32376 260800 32428
rect 379520 32376 379572 32428
rect 384948 32376 385000 32428
rect 560300 32376 560352 32428
rect 96252 31764 96304 31816
rect 96160 31696 96212 31748
rect 198004 31696 198056 31748
rect 198188 31696 198240 31748
rect 267004 31696 267056 31748
rect 267188 31696 267240 31748
rect 567844 31696 567896 31748
rect 568028 31696 568080 31748
rect 354588 31084 354640 31136
rect 516140 31084 516192 31136
rect 111064 31016 111116 31068
rect 162860 31016 162912 31068
rect 173808 31016 173860 31068
rect 253940 31016 253992 31068
rect 255228 31016 255280 31068
rect 372620 31016 372672 31068
rect 380716 31016 380768 31068
rect 553400 31016 553452 31068
rect 402244 30268 402296 30320
rect 580172 30268 580224 30320
rect 248236 29656 248288 29708
rect 361580 29656 361632 29708
rect 106096 29588 106148 29640
rect 158812 29588 158864 29640
rect 168288 29588 168340 29640
rect 247040 29588 247092 29640
rect 288348 29588 288400 29640
rect 419540 29588 419592 29640
rect 198188 28908 198240 28960
rect 267188 28908 267240 28960
rect 337936 28296 337988 28348
rect 491300 28296 491352 28348
rect 90916 28228 90968 28280
rect 133880 28228 133932 28280
rect 158628 28228 158680 28280
rect 233240 28228 233292 28280
rect 236644 28228 236696 28280
rect 343640 28228 343692 28280
rect 361488 28228 361540 28280
rect 524512 28228 524564 28280
rect 215116 27616 215168 27668
rect 227444 27616 227496 27668
rect 138020 27548 138072 27600
rect 138480 27548 138532 27600
rect 198740 27548 198792 27600
rect 509240 27591 509292 27600
rect 509240 27557 509249 27591
rect 509249 27557 509283 27591
rect 509283 27557 509292 27591
rect 509240 27548 509292 27557
rect 518900 27591 518952 27600
rect 518900 27557 518909 27591
rect 518909 27557 518943 27591
rect 518943 27557 518952 27591
rect 518900 27548 518952 27557
rect 527180 27591 527232 27600
rect 527180 27557 527189 27591
rect 527189 27557 527223 27591
rect 527223 27557 527232 27591
rect 527180 27548 527232 27557
rect 532700 27591 532752 27600
rect 532700 27557 532709 27591
rect 532709 27557 532743 27591
rect 532743 27557 532752 27591
rect 532700 27548 532752 27557
rect 568028 27591 568080 27600
rect 568028 27557 568037 27591
rect 568037 27557 568071 27591
rect 568071 27557 568080 27591
rect 568028 27548 568080 27557
rect 569960 27591 570012 27600
rect 569960 27557 569969 27591
rect 569969 27557 570003 27591
rect 570003 27557 570012 27591
rect 569960 27548 570012 27557
rect 335268 26936 335320 26988
rect 487160 26936 487212 26988
rect 104808 26868 104860 26920
rect 154580 26868 154632 26920
rect 155868 26868 155920 26920
rect 229100 26868 229152 26920
rect 230388 26868 230440 26920
rect 336740 26868 336792 26920
rect 353208 26868 353260 26920
rect 513380 26868 513432 26920
rect 332508 25576 332560 25628
rect 484400 25576 484452 25628
rect 102048 25508 102100 25560
rect 150532 25508 150584 25560
rect 154488 25508 154540 25560
rect 226340 25508 226392 25560
rect 227444 25508 227496 25560
rect 332600 25508 332652 25560
rect 350448 25508 350500 25560
rect 510712 25508 510764 25560
rect 224224 24148 224276 24200
rect 318800 24148 318852 24200
rect 324136 24148 324188 24200
rect 471980 24148 472032 24200
rect 99196 24080 99248 24132
rect 147680 24080 147732 24132
rect 151728 24080 151780 24132
rect 222200 24080 222252 24132
rect 234528 24080 234580 24132
rect 342260 24080 342312 24132
rect 343548 24080 343600 24132
rect 499580 24080 499632 24132
rect 200120 22831 200172 22840
rect 200120 22797 200129 22831
rect 200129 22797 200163 22831
rect 200163 22797 200172 22831
rect 200120 22788 200172 22797
rect 215116 22788 215168 22840
rect 314660 22788 314712 22840
rect 321376 22788 321428 22840
rect 467932 22788 467984 22840
rect 96160 22720 96212 22772
rect 143540 22720 143592 22772
rect 148968 22720 149020 22772
rect 218152 22720 218204 22772
rect 227628 22720 227680 22772
rect 331312 22720 331364 22772
rect 338028 22720 338080 22772
rect 492680 22720 492732 22772
rect 267740 22695 267792 22704
rect 267740 22661 267749 22695
rect 267749 22661 267783 22695
rect 267783 22661 267792 22695
rect 267740 22652 267792 22661
rect 3148 22040 3200 22092
rect 79416 22040 79468 22092
rect 208308 21428 208360 21480
rect 305092 21428 305144 21480
rect 318064 21428 318116 21480
rect 454040 21428 454092 21480
rect 88984 21360 89036 21412
rect 131120 21360 131172 21412
rect 143448 21360 143500 21412
rect 211160 21360 211212 21412
rect 217968 21360 218020 21412
rect 317420 21360 317472 21412
rect 326344 21360 326396 21412
rect 473360 21360 473412 21412
rect 142068 20000 142120 20052
rect 208400 20000 208452 20052
rect 304908 20000 304960 20052
rect 443092 20000 443144 20052
rect 446404 20000 446456 20052
rect 571432 20000 571484 20052
rect 97264 19932 97316 19984
rect 140872 19932 140924 19984
rect 205548 19932 205600 19984
rect 300860 19932 300912 19984
rect 320088 19932 320140 19984
rect 466460 19932 466512 19984
rect 198096 19363 198148 19372
rect 198096 19329 198105 19363
rect 198105 19329 198139 19363
rect 198139 19329 198148 19363
rect 198096 19320 198148 19329
rect 267096 19363 267148 19372
rect 267096 19329 267105 19363
rect 267105 19329 267139 19363
rect 267139 19329 267148 19363
rect 267096 19320 267148 19329
rect 491300 19295 491352 19304
rect 491300 19261 491309 19295
rect 491309 19261 491343 19295
rect 491343 19261 491352 19295
rect 491300 19252 491352 19261
rect 492680 19295 492732 19304
rect 492680 19261 492689 19295
rect 492689 19261 492723 19295
rect 492723 19261 492732 19295
rect 510620 19295 510672 19304
rect 492680 19252 492732 19261
rect 510620 19261 510629 19295
rect 510629 19261 510663 19295
rect 510663 19261 510672 19295
rect 510620 19252 510672 19261
rect 516140 19295 516192 19304
rect 516140 19261 516149 19295
rect 516149 19261 516183 19295
rect 516183 19261 516192 19295
rect 516140 19252 516192 19261
rect 547880 19252 547932 19304
rect 548892 19252 548944 19304
rect 550640 19295 550692 19304
rect 550640 19261 550649 19295
rect 550649 19261 550683 19295
rect 550683 19261 550692 19295
rect 553400 19295 553452 19304
rect 550640 19252 550692 19261
rect 553400 19261 553409 19295
rect 553409 19261 553443 19295
rect 553443 19261 553452 19295
rect 553400 19252 553452 19261
rect 560300 19252 560352 19304
rect 560760 19252 560812 19304
rect 283564 18708 283616 18760
rect 400312 18708 400364 18760
rect 269028 18640 269080 18692
rect 390652 18640 390704 18692
rect 92388 18572 92440 18624
rect 136640 18572 136692 18624
rect 139308 18572 139360 18624
rect 204260 18572 204312 18624
rect 207664 18572 207716 18624
rect 296812 18572 296864 18624
rect 380808 18572 380860 18624
rect 554872 18572 554924 18624
rect 518900 18003 518952 18012
rect 518900 17969 518909 18003
rect 518909 17969 518943 18003
rect 518943 17969 518952 18003
rect 518900 17960 518952 17969
rect 527180 18003 527232 18012
rect 527180 17969 527189 18003
rect 527189 17969 527223 18003
rect 527223 17969 527232 18003
rect 527180 17960 527232 17969
rect 568028 18003 568080 18012
rect 568028 17969 568037 18003
rect 568037 17969 568071 18003
rect 568071 17969 568080 18003
rect 568028 17960 568080 17969
rect 555424 17892 555476 17944
rect 579804 17892 579856 17944
rect 257988 17348 258040 17400
rect 376760 17348 376812 17400
rect 136548 17280 136600 17332
rect 201592 17280 201644 17332
rect 272524 17280 272576 17332
rect 396080 17280 396132 17332
rect 89628 17212 89680 17264
rect 132592 17212 132644 17264
rect 201408 17212 201460 17264
rect 293960 17212 294012 17264
rect 376668 17212 376720 17264
rect 546500 17212 546552 17264
rect 344284 15988 344336 16040
rect 451372 15988 451424 16040
rect 195888 15920 195940 15972
rect 287152 15920 287204 15972
rect 291108 15920 291160 15972
rect 425152 15920 425204 15972
rect 86868 15852 86920 15904
rect 129740 15852 129792 15904
rect 131764 15852 131816 15904
rect 193312 15852 193364 15904
rect 261484 15852 261536 15904
rect 374092 15852 374144 15904
rect 398748 15852 398800 15904
rect 578976 15852 579028 15904
rect 527180 14832 527232 14884
rect 527364 14832 527416 14884
rect 193128 14492 193180 14544
rect 282920 14492 282972 14544
rect 333796 14492 333848 14544
rect 485872 14492 485924 14544
rect 85488 14424 85540 14476
rect 126980 14424 127032 14476
rect 129648 14424 129700 14476
rect 190460 14424 190512 14476
rect 251088 14424 251140 14476
rect 365812 14424 365864 14476
rect 386328 14424 386380 14476
rect 561956 14424 562008 14476
rect 106924 13132 106976 13184
rect 128360 13132 128412 13184
rect 188988 13132 189040 13184
rect 276020 13132 276072 13184
rect 294604 13132 294656 13184
rect 382280 13132 382332 13184
rect 126888 13064 126940 13116
rect 186320 13064 186372 13116
rect 248328 13064 248380 13116
rect 362960 13064 363012 13116
rect 373908 13064 373960 13116
rect 544108 13064 544160 13116
rect 517520 12452 517572 12504
rect 518900 12452 518952 12504
rect 524420 12452 524472 12504
rect 545120 12452 545172 12504
rect 568580 12452 568632 12504
rect 133880 12384 133932 12436
rect 134800 12384 134852 12436
rect 136640 12384 136692 12436
rect 137192 12384 137244 12436
rect 143540 12384 143592 12436
rect 144460 12384 144512 12436
rect 144920 12384 144972 12436
rect 145656 12384 145708 12436
rect 195980 12384 196032 12436
rect 196808 12384 196860 12436
rect 202880 12384 202932 12436
rect 203892 12384 203944 12436
rect 204260 12384 204312 12436
rect 205088 12384 205140 12436
rect 263600 12384 263652 12436
rect 264612 12384 264664 12436
rect 266360 12384 266412 12436
rect 267004 12384 267056 12436
rect 270592 12384 270644 12436
rect 271696 12384 271748 12436
rect 487160 12384 487212 12436
rect 488172 12384 488224 12436
rect 488540 12384 488592 12436
rect 489368 12384 489420 12436
rect 505100 12384 505152 12436
rect 506020 12384 506072 12436
rect 506480 12384 506532 12436
rect 507216 12384 507268 12436
rect 513380 12384 513432 12436
rect 514392 12384 514444 12436
rect 514760 12384 514812 12436
rect 515588 12384 515640 12436
rect 517888 12316 517940 12368
rect 521660 12384 521712 12436
rect 522672 12384 522724 12436
rect 523040 12384 523092 12436
rect 523868 12384 523920 12436
rect 519084 12316 519136 12368
rect 529940 12384 529992 12436
rect 531044 12384 531096 12436
rect 531320 12384 531372 12436
rect 532240 12384 532292 12436
rect 525064 12316 525116 12368
rect 549260 12384 549312 12436
rect 550088 12384 550140 12436
rect 557540 12384 557592 12436
rect 558368 12384 558420 12436
rect 564440 12384 564492 12436
rect 565544 12384 565596 12436
rect 565820 12384 565872 12436
rect 566740 12384 566792 12436
rect 569040 12384 569092 12436
rect 545304 12316 545356 12368
rect 551192 12316 551244 12368
rect 552112 12316 552164 12368
rect 552388 12316 552440 12368
rect 186228 11840 186280 11892
rect 272892 11840 272944 11892
rect 241428 11772 241480 11824
rect 351920 11772 351972 11824
rect 363604 11772 363656 11824
rect 526260 11772 526312 11824
rect 124128 11704 124180 11756
rect 183560 11704 183612 11756
rect 259368 11704 259420 11756
rect 378140 11704 378192 11756
rect 390468 11704 390520 11756
rect 567844 11704 567896 11756
rect 266268 10412 266320 10464
rect 389180 10412 389232 10464
rect 183468 10344 183520 10396
rect 269304 10344 269356 10396
rect 351828 10344 351880 10396
rect 512092 10344 512144 10396
rect 121368 10276 121420 10328
rect 179420 10276 179472 10328
rect 246304 10276 246356 10328
rect 347872 10276 347924 10328
rect 383568 10276 383620 10328
rect 557172 10276 557224 10328
rect 199200 9664 199252 9716
rect 200396 9664 200448 9716
rect 268108 9664 268160 9716
rect 491760 9664 491812 9716
rect 492956 9664 493008 9716
rect 509608 9664 509660 9716
rect 510804 9664 510856 9716
rect 516784 9664 516836 9716
rect 533436 9664 533488 9716
rect 553584 9664 553636 9716
rect 570236 9664 570288 9716
rect 517888 9639 517940 9648
rect 517888 9605 517897 9639
rect 517897 9605 517931 9639
rect 517931 9605 517940 9639
rect 517888 9596 517940 9605
rect 519084 9639 519136 9648
rect 519084 9605 519093 9639
rect 519093 9605 519127 9639
rect 519127 9605 519136 9639
rect 519084 9596 519136 9605
rect 525064 9596 525116 9648
rect 527456 9596 527508 9648
rect 545304 9639 545356 9648
rect 545304 9605 545313 9639
rect 545313 9605 545347 9639
rect 545347 9605 545356 9639
rect 545304 9596 545356 9605
rect 548892 9639 548944 9648
rect 548892 9605 548901 9639
rect 548901 9605 548935 9639
rect 548935 9605 548944 9639
rect 548892 9596 548944 9605
rect 550088 9639 550140 9648
rect 550088 9605 550097 9639
rect 550097 9605 550131 9639
rect 550131 9605 550140 9639
rect 550088 9596 550140 9605
rect 525064 9460 525116 9512
rect 527456 9460 527508 9512
rect 171048 9052 171100 9104
rect 251456 9052 251508 9104
rect 223488 8984 223540 9036
rect 327632 8984 327684 9036
rect 349068 8984 349120 9036
rect 508412 8984 508464 9036
rect 118608 8916 118660 8968
rect 176568 8916 176620 8968
rect 244188 8916 244240 8968
rect 357348 8916 357400 8968
rect 375288 8916 375340 8968
rect 546592 8916 546644 8968
rect 135904 8644 135956 8696
rect 3424 8236 3476 8288
rect 79324 8236 79376 8288
rect 174544 7692 174596 7744
rect 244372 7692 244424 7744
rect 132592 7624 132644 7676
rect 133788 7624 133840 7676
rect 140780 7624 140832 7676
rect 142068 7624 142120 7676
rect 222108 7624 222160 7676
rect 324044 7624 324096 7676
rect 339408 7624 339460 7676
rect 494152 7692 494204 7744
rect 494060 7624 494112 7676
rect 495348 7624 495400 7676
rect 512000 7624 512052 7676
rect 513196 7624 513248 7676
rect 117228 7556 117280 7608
rect 172980 7556 173032 7608
rect 201500 7556 201552 7608
rect 202696 7556 202748 7608
rect 240048 7556 240100 7608
rect 350264 7556 350316 7608
rect 362868 7556 362920 7608
rect 485780 7488 485832 7540
rect 486976 7488 487028 7540
rect 528560 7556 528612 7608
rect 529848 7556 529900 7608
rect 546500 7556 546552 7608
rect 547696 7556 547748 7608
rect 554780 7556 554832 7608
rect 555976 7556 556028 7608
rect 563152 7556 563204 7608
rect 564348 7556 564400 7608
rect 571340 7556 571392 7608
rect 572628 7556 572680 7608
rect 528652 7488 528704 7540
rect 482192 7284 482244 7336
rect 161388 6196 161440 6248
rect 237196 6196 237248 6248
rect 336648 6196 336700 6248
rect 490564 6196 490616 6248
rect 111708 6128 111760 6180
rect 165896 6128 165948 6180
rect 233148 6128 233200 6180
rect 340696 6128 340748 6180
rect 358728 6128 358780 6180
rect 521476 6128 521528 6180
rect 84108 4836 84160 4888
rect 126612 4836 126664 4888
rect 178684 4836 178736 4888
rect 198004 4836 198056 4888
rect 198188 4836 198240 4888
rect 253848 4836 253900 4888
rect 291844 4836 291896 4888
rect 383568 4836 383620 4888
rect 420184 4836 420236 4888
rect 483480 4836 483532 4888
rect 125508 4768 125560 4820
rect 144920 4768 144972 4820
rect 145012 4768 145064 4820
rect 184848 4768 184900 4820
rect 203524 4768 203576 4820
rect 265808 4768 265860 4820
rect 267188 4768 267240 4820
rect 290740 4768 290792 4820
rect 298008 4768 298060 4820
rect 434628 4768 434680 4820
rect 493324 4768 493376 4820
rect 559564 4768 559616 4820
rect 347872 4156 347924 4208
rect 349068 4156 349120 4208
rect 400220 4156 400272 4208
rect 401324 4156 401376 4208
rect 408500 4156 408552 4208
rect 409696 4156 409748 4208
rect 306288 4088 306340 4140
rect 446588 4088 446640 4140
rect 309048 4020 309100 4072
rect 450176 4020 450228 4072
rect 88248 3952 88300 4004
rect 132592 3952 132644 4004
rect 311808 3952 311860 4004
rect 453672 3952 453724 4004
rect 91008 3884 91060 3936
rect 136088 3884 136140 3936
rect 162308 3884 162360 3936
rect 315948 3884 316000 3936
rect 460848 3884 460900 3936
rect 93768 3816 93820 3868
rect 139676 3816 139728 3868
rect 313188 3816 313240 3868
rect 457260 3816 457312 3868
rect 96528 3748 96580 3800
rect 143264 3748 143316 3800
rect 318708 3748 318760 3800
rect 464436 3748 464488 3800
rect 99288 3680 99340 3732
rect 146852 3680 146904 3732
rect 321468 3680 321520 3732
rect 467840 3680 467892 3732
rect 103428 3612 103480 3664
rect 153936 3612 153988 3664
rect 324228 3612 324280 3664
rect 471520 3612 471572 3664
rect 100668 3544 100720 3596
rect 150440 3544 150492 3596
rect 218152 3544 218204 3596
rect 219348 3544 219400 3596
rect 227720 3544 227772 3596
rect 228916 3544 228968 3596
rect 262220 3544 262272 3596
rect 263416 3544 263468 3596
rect 278872 3544 278924 3596
rect 280068 3544 280120 3596
rect 305000 3544 305052 3596
rect 306196 3544 306248 3596
rect 313372 3544 313424 3596
rect 314568 3544 314620 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 325608 3544 325660 3596
rect 475108 3544 475160 3596
rect 502432 3544 502484 3596
rect 503628 3544 503680 3596
rect 536932 3544 536984 3596
rect 538128 3544 538180 3596
rect 568212 3544 568264 3596
rect 572 3476 624 3528
rect 81440 3476 81492 3528
rect 106188 3476 106240 3528
rect 157524 3476 157576 3528
rect 158720 3476 158772 3528
rect 159916 3476 159968 3528
rect 167000 3476 167052 3528
rect 168196 3476 168248 3528
rect 209780 3476 209832 3528
rect 211068 3476 211120 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 328368 3476 328420 3528
rect 478696 3476 478748 3528
rect 1676 3408 1728 3460
rect 82912 3408 82964 3460
rect 108948 3408 109000 3460
rect 161112 3408 161164 3460
rect 331128 3408 331180 3460
rect 482284 3408 482336 3460
rect 578608 3476 578660 3528
rect 578976 3476 579028 3528
rect 579804 3476 579856 3528
rect 374000 3340 374052 3392
rect 375196 3340 375248 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 425060 3340 425112 3392
rect 426348 3340 426400 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 582196 3272 582248 3324
rect 578884 3136 578936 3188
rect 581000 3136 581052 3188
rect 287060 1368 287112 1420
rect 288348 1368 288400 1420
rect 126980 552 127032 604
rect 127808 552 127860 604
rect 128360 552 128412 604
rect 129004 552 129056 604
rect 131120 552 131172 604
rect 131396 552 131448 604
rect 200396 552 200448 604
rect 200488 552 200540 604
rect 306380 552 306432 604
rect 307392 552 307444 604
rect 307760 552 307812 604
rect 308588 552 308640 604
rect 309140 552 309192 604
rect 309784 552 309836 604
rect 310520 552 310572 604
rect 310980 552 311032 604
rect 314660 552 314712 604
rect 315764 552 315816 604
rect 517888 595 517940 604
rect 517888 561 517897 595
rect 517897 561 517931 595
rect 517931 561 517940 595
rect 517888 552 517940 561
rect 519084 595 519136 604
rect 519084 561 519093 595
rect 519093 561 519127 595
rect 519127 561 519136 595
rect 519084 552 519136 561
rect 545304 595 545356 604
rect 545304 561 545313 595
rect 545313 561 545347 595
rect 545347 561 545356 595
rect 545304 552 545356 561
rect 548892 595 548944 604
rect 548892 561 548901 595
rect 548901 561 548935 595
rect 548935 561 548944 595
rect 548892 552 548944 561
rect 550088 595 550140 604
rect 550088 561 550097 595
rect 550097 561 550131 595
rect 550131 561 550140 595
rect 550088 552 550140 561
rect 576860 552 576912 604
rect 577412 552 577464 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 8128 679046 8156 685850
rect 8944 681760 8996 681766
rect 8944 681702 8996 681708
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3238 624880 3294 624889
rect 3238 624815 3294 624824
rect 3252 623830 3280 624815
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 3054 452432 3110 452441
rect 3054 452367 3110 452376
rect 3068 451314 3096 452367
rect 3056 451308 3108 451314
rect 3056 451250 3108 451256
rect 3330 423736 3386 423745
rect 3330 423671 3332 423680
rect 3384 423671 3386 423680
rect 3332 423642 3384 423648
rect 3436 411262 3464 667927
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 3514 610464 3570 610473
rect 3514 610399 3570 610408
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3160 394738 3188 394975
rect 3148 394732 3200 394738
rect 3148 394674 3200 394680
rect 3528 389162 3556 610399
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 589286 8064 591926
rect 8024 589280 8076 589286
rect 8024 589222 8076 589228
rect 8024 579760 8076 579766
rect 7944 579708 8024 579714
rect 7944 579702 8076 579708
rect 7944 579686 8064 579702
rect 7944 579630 7972 579686
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 8116 579624 8168 579630
rect 8116 579566 8168 579572
rect 4066 567352 4122 567361
rect 4066 567287 4122 567296
rect 4080 567254 4108 567287
rect 4068 567248 4120 567254
rect 4068 567190 4120 567196
rect 8128 562970 8156 579566
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 8116 562964 8168 562970
rect 8116 562906 8168 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 3606 553072 3662 553081
rect 3606 553007 3662 553016
rect 3516 389156 3568 389162
rect 3516 389098 3568 389104
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3054 337512 3110 337521
rect 3054 337447 3110 337456
rect 3068 336802 3096 337447
rect 3056 336796 3108 336802
rect 3056 336738 3108 336744
rect 3436 296682 3464 380559
rect 3514 366208 3570 366217
rect 3514 366143 3570 366152
rect 3424 296676 3476 296682
rect 3424 296618 3476 296624
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3436 259418 3464 294335
rect 3528 289814 3556 366143
rect 3620 365702 3648 553007
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8208 541000 8260 541006
rect 8208 540942 8260 540948
rect 4066 538656 4122 538665
rect 4066 538591 4122 538600
rect 4080 538286 4108 538591
rect 4068 538280 4120 538286
rect 4068 538222 4120 538228
rect 8220 534018 8248 540942
rect 8128 533990 8248 534018
rect 8128 531321 8156 533990
rect 8114 531312 8170 531321
rect 8114 531247 8170 531256
rect 8390 531312 8446 531321
rect 8390 531247 8446 531256
rect 8404 521694 8432 531247
rect 8208 521688 8260 521694
rect 8208 521630 8260 521636
rect 8392 521688 8444 521694
rect 8392 521630 8444 521636
rect 8220 514706 8248 521630
rect 8128 514678 8248 514706
rect 8128 512009 8156 514678
rect 8114 512000 8170 512009
rect 8114 511935 8170 511944
rect 8390 512000 8446 512009
rect 8390 511935 8446 511944
rect 3882 509960 3938 509969
rect 3882 509895 3938 509904
rect 3896 509318 3924 509895
rect 3884 509312 3936 509318
rect 3884 509254 3936 509260
rect 8404 502382 8432 511935
rect 8208 502376 8260 502382
rect 8208 502318 8260 502324
rect 8392 502376 8444 502382
rect 8392 502318 8444 502324
rect 3698 495544 3754 495553
rect 3698 495479 3754 495488
rect 3608 365696 3660 365702
rect 3608 365638 3660 365644
rect 3712 343602 3740 495479
rect 8220 495394 8248 502318
rect 8128 495366 8248 495394
rect 8128 492658 8156 495366
rect 7932 492652 7984 492658
rect 7932 492594 7984 492600
rect 8116 492652 8168 492658
rect 8116 492594 8168 492600
rect 7944 483041 7972 492594
rect 7930 483032 7986 483041
rect 7930 482967 7986 482976
rect 8206 483032 8262 483041
rect 8206 482967 8262 482976
rect 8220 476082 8248 482967
rect 8036 476054 8248 476082
rect 8036 473346 8064 476054
rect 8024 473340 8076 473346
rect 8024 473282 8076 473288
rect 8116 473340 8168 473346
rect 8116 473282 8168 473288
rect 8128 463706 8156 473282
rect 8128 463678 8248 463706
rect 8220 456770 8248 463678
rect 8036 456742 8248 456770
rect 6184 451308 6236 451314
rect 6184 451250 6236 451256
rect 3790 438016 3846 438025
rect 3790 437951 3846 437960
rect 3700 343596 3752 343602
rect 3700 343538 3752 343544
rect 3606 323096 3662 323105
rect 3606 323031 3662 323040
rect 3516 289808 3568 289814
rect 3516 289750 3568 289756
rect 3514 280120 3570 280129
rect 3514 280055 3570 280064
rect 3424 259412 3476 259418
rect 3424 259354 3476 259360
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3436 235958 3464 251223
rect 3528 251190 3556 280055
rect 3620 274650 3648 323031
rect 3804 320142 3832 437951
rect 6196 327078 6224 451250
rect 8036 447166 8064 456742
rect 8024 447160 8076 447166
rect 8024 447102 8076 447108
rect 8116 447092 8168 447098
rect 8116 447034 8168 447040
rect 8128 444378 8156 447034
rect 8116 444372 8168 444378
rect 8116 444314 8168 444320
rect 8116 437436 8168 437442
rect 8116 437378 8168 437384
rect 8128 434738 8156 437378
rect 8128 434710 8248 434738
rect 8220 425134 8248 434710
rect 8024 425128 8076 425134
rect 8024 425070 8076 425076
rect 8208 425128 8260 425134
rect 8208 425070 8260 425076
rect 8036 424386 8064 425070
rect 8024 424380 8076 424386
rect 8024 424322 8076 424328
rect 7564 423700 7616 423706
rect 7564 423642 7616 423648
rect 6184 327072 6236 327078
rect 6184 327014 6236 327020
rect 3792 320136 3844 320142
rect 3792 320078 3844 320084
rect 7576 311846 7604 423642
rect 8956 419490 8984 681702
rect 14464 652792 14516 652798
rect 14464 652734 14516 652740
rect 13084 567248 13136 567254
rect 13084 567190 13136 567196
rect 10324 480276 10376 480282
rect 10324 480218 10376 480224
rect 8944 419484 8996 419490
rect 8944 419426 8996 419432
rect 10336 335306 10364 480218
rect 13096 373998 13124 567190
rect 14476 404326 14504 652734
rect 17224 538280 17276 538286
rect 17224 538222 17276 538228
rect 14464 404320 14516 404326
rect 14464 404262 14516 404268
rect 13084 373992 13136 373998
rect 13084 373934 13136 373940
rect 17236 358766 17264 538222
rect 24780 424454 24808 699654
rect 29644 623824 29696 623830
rect 29644 623766 29696 623772
rect 24768 424448 24820 424454
rect 24768 424390 24820 424396
rect 29656 396030 29684 623766
rect 39304 509312 39356 509318
rect 39304 509254 39356 509260
rect 29644 396024 29696 396030
rect 29644 395966 29696 395972
rect 21364 394732 21416 394738
rect 21364 394674 21416 394680
rect 17224 358760 17276 358766
rect 17224 358702 17276 358708
rect 10324 335300 10376 335306
rect 10324 335242 10376 335248
rect 7564 311840 7616 311846
rect 7564 311782 7616 311788
rect 3698 308816 3754 308825
rect 3698 308751 3754 308760
rect 3608 274644 3660 274650
rect 3608 274586 3660 274592
rect 3712 266354 3740 308751
rect 21376 304978 21404 394674
rect 39316 350538 39344 509254
rect 41340 424522 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 72884 637560 72936 637566
rect 72884 637502 72936 637508
rect 72896 630578 72924 637502
rect 72896 630550 73108 630578
rect 73080 626550 73108 630550
rect 73068 626544 73120 626550
rect 73068 626486 73120 626492
rect 73068 616888 73120 616894
rect 73068 616830 73120 616836
rect 73080 611454 73108 616830
rect 73068 611448 73120 611454
rect 73068 611390 73120 611396
rect 72884 611312 72936 611318
rect 72884 611254 72936 611260
rect 72896 608546 72924 611254
rect 72974 608560 73030 608569
rect 72896 608518 72974 608546
rect 72974 608495 73030 608504
rect 73158 608560 73214 608569
rect 73158 608495 73214 608504
rect 73172 601594 73200 608495
rect 72976 601588 73028 601594
rect 72976 601530 73028 601536
rect 73160 601588 73212 601594
rect 73160 601530 73212 601536
rect 72988 598942 73016 601530
rect 72976 598936 73028 598942
rect 72976 598878 73028 598884
rect 44824 594856 44876 594862
rect 44824 594798 44876 594804
rect 41328 424516 41380 424522
rect 41328 424458 41380 424464
rect 44836 380866 44864 594798
rect 72884 589348 72936 589354
rect 72884 589290 72936 589296
rect 72896 582418 72924 589290
rect 72700 582412 72752 582418
rect 72700 582354 72752 582360
rect 72884 582412 72936 582418
rect 72884 582354 72936 582360
rect 72712 579630 72740 582354
rect 72700 579624 72752 579630
rect 72700 579566 72752 579572
rect 72608 569968 72660 569974
rect 72608 569910 72660 569916
rect 72620 563106 72648 569910
rect 72608 563100 72660 563106
rect 72608 563042 72660 563048
rect 72700 562964 72752 562970
rect 72700 562906 72752 562912
rect 72712 560266 72740 562906
rect 72620 560238 72740 560266
rect 72620 553450 72648 560238
rect 72608 553444 72660 553450
rect 72608 553386 72660 553392
rect 72608 550656 72660 550662
rect 72608 550598 72660 550604
rect 72620 543794 72648 550598
rect 72608 543788 72660 543794
rect 72608 543730 72660 543736
rect 72700 543652 72752 543658
rect 72700 543594 72752 543600
rect 72712 540954 72740 543594
rect 72620 540926 72740 540954
rect 72620 534138 72648 540926
rect 72608 534132 72660 534138
rect 72608 534074 72660 534080
rect 72620 531350 72648 531381
rect 72608 531344 72660 531350
rect 72698 531312 72754 531321
rect 72660 531292 72698 531298
rect 72608 531286 72698 531292
rect 72620 531270 72698 531286
rect 72698 531247 72754 531256
rect 72882 531312 72938 531321
rect 72882 531247 72938 531256
rect 72896 524346 72924 531247
rect 72700 524340 72752 524346
rect 72700 524282 72752 524288
rect 72884 524340 72936 524346
rect 72884 524282 72936 524288
rect 72712 514706 72740 524282
rect 72712 514678 72832 514706
rect 72804 512009 72832 514678
rect 72606 512000 72662 512009
rect 72606 511935 72662 511944
rect 72790 512000 72846 512009
rect 72790 511935 72846 511944
rect 72620 502382 72648 511935
rect 72608 502376 72660 502382
rect 72608 502318 72660 502324
rect 73068 502376 73120 502382
rect 73068 502318 73120 502324
rect 73080 495394 73108 502318
rect 72988 495366 73108 495394
rect 72988 485874 73016 495366
rect 72896 485846 73016 485874
rect 72896 480282 72924 485846
rect 72884 480276 72936 480282
rect 72884 480218 72936 480224
rect 73068 480276 73120 480282
rect 73068 480218 73120 480224
rect 73080 480162 73108 480218
rect 72988 480134 73108 480162
rect 72988 470642 73016 480134
rect 72896 470614 73016 470642
rect 72896 460970 72924 470614
rect 72884 460964 72936 460970
rect 72884 460906 72936 460912
rect 73068 460964 73120 460970
rect 73068 460906 73120 460912
rect 73080 460850 73108 460906
rect 72988 460822 73108 460850
rect 72988 437510 73016 460822
rect 72792 437504 72844 437510
rect 72792 437446 72844 437452
rect 72976 437504 73028 437510
rect 72976 437446 73028 437452
rect 72804 424590 72832 437446
rect 72792 424584 72844 424590
rect 72792 424526 72844 424532
rect 89640 424386 89668 699654
rect 106200 424454 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 137756 596222 137784 605798
rect 154316 596222 154344 605798
rect 137744 596216 137796 596222
rect 137928 596216 137980 596222
rect 137744 596158 137796 596164
rect 137848 596164 137928 596170
rect 137848 596158 137980 596164
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 137848 596142 137968 596158
rect 154408 596142 154528 596158
rect 137848 591954 137876 596142
rect 154408 591954 154436 596142
rect 137756 591926 137876 591954
rect 154316 591926 154436 591954
rect 137756 589286 137784 591926
rect 154316 589286 154344 591926
rect 137744 589280 137796 589286
rect 137744 589222 137796 589228
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 137744 579760 137796 579766
rect 137664 579708 137744 579714
rect 154304 579760 154356 579766
rect 137664 579702 137796 579708
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 137664 579686 137784 579702
rect 154224 579686 154344 579702
rect 137664 579630 137692 579686
rect 154224 579630 154252 579686
rect 137652 579624 137704 579630
rect 137652 579566 137704 579572
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 137560 569968 137612 569974
rect 137560 569910 137612 569916
rect 137572 563106 137600 569910
rect 137560 563100 137612 563106
rect 137560 563042 137612 563048
rect 154408 562970 154436 579566
rect 137652 562964 137704 562970
rect 137652 562906 137704 562912
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 137664 560250 137692 562906
rect 137652 560244 137704 560250
rect 137652 560186 137704 560192
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 137836 550656 137888 550662
rect 137836 550598 137888 550604
rect 137848 543658 137876 550598
rect 154316 543810 154344 553302
rect 154316 543782 154528 543810
rect 137652 543652 137704 543658
rect 137652 543594 137704 543600
rect 137836 543652 137888 543658
rect 137836 543594 137888 543600
rect 137664 534070 137692 543594
rect 137652 534064 137704 534070
rect 137652 534006 137704 534012
rect 137836 534064 137888 534070
rect 154500 534018 154528 543782
rect 137836 534006 137888 534012
rect 137848 531321 137876 534006
rect 154408 533990 154528 534018
rect 137834 531312 137890 531321
rect 137834 531247 137890 531256
rect 138110 531312 138166 531321
rect 154408 531282 154436 533990
rect 138110 531247 138166 531256
rect 154396 531276 154448 531282
rect 138124 521694 138152 531247
rect 154396 531218 154448 531224
rect 137928 521688 137980 521694
rect 137928 521630 137980 521636
rect 138112 521688 138164 521694
rect 138112 521630 138164 521636
rect 154488 521688 154540 521694
rect 154488 521630 154540 521636
rect 137940 514706 137968 521630
rect 154500 514706 154528 521630
rect 137848 514678 137968 514706
rect 154408 514678 154528 514706
rect 137848 512009 137876 514678
rect 137834 512000 137890 512009
rect 137834 511935 137890 511944
rect 138110 512000 138166 512009
rect 154408 511970 154436 514678
rect 138110 511935 138166 511944
rect 154396 511964 154448 511970
rect 138124 502382 138152 511935
rect 154396 511906 154448 511912
rect 137928 502376 137980 502382
rect 137928 502318 137980 502324
rect 138112 502376 138164 502382
rect 138112 502318 138164 502324
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 137940 495394 137968 502318
rect 154500 495394 154528 502318
rect 137848 495366 137968 495394
rect 154408 495366 154528 495394
rect 137848 492658 137876 495366
rect 154408 492658 154436 495366
rect 137652 492652 137704 492658
rect 137652 492594 137704 492600
rect 137836 492652 137888 492658
rect 137836 492594 137888 492600
rect 154212 492652 154264 492658
rect 154212 492594 154264 492600
rect 154396 492652 154448 492658
rect 154396 492594 154448 492600
rect 137664 483041 137692 492594
rect 154224 483041 154252 492594
rect 137650 483032 137706 483041
rect 137650 482967 137706 482976
rect 137926 483032 137982 483041
rect 137926 482967 137982 482976
rect 154210 483032 154266 483041
rect 154210 482967 154266 482976
rect 154486 483032 154542 483041
rect 154486 482967 154542 482976
rect 137940 476082 137968 482967
rect 154500 476082 154528 482967
rect 137756 476054 137968 476082
rect 154316 476054 154528 476082
rect 137756 473346 137784 476054
rect 137468 473340 137520 473346
rect 137468 473282 137520 473288
rect 137744 473340 137796 473346
rect 137744 473282 137796 473288
rect 137480 463729 137508 473282
rect 154316 466478 154344 476054
rect 154304 466472 154356 466478
rect 154304 466414 154356 466420
rect 154488 466472 154540 466478
rect 154488 466414 154540 466420
rect 137466 463720 137522 463729
rect 137466 463655 137522 463664
rect 137650 463720 137706 463729
rect 137650 463655 137706 463664
rect 137664 456770 137692 463655
rect 154500 456770 154528 466414
rect 137664 456742 137784 456770
rect 137756 447166 137784 456742
rect 154316 456742 154528 456770
rect 154316 447166 154344 456742
rect 137744 447160 137796 447166
rect 137744 447102 137796 447108
rect 154304 447160 154356 447166
rect 154304 447102 154356 447108
rect 137836 447092 137888 447098
rect 137836 447034 137888 447040
rect 154396 447092 154448 447098
rect 154396 447034 154448 447040
rect 137848 444378 137876 447034
rect 154408 444378 154436 447034
rect 137836 444372 137888 444378
rect 137836 444314 137888 444320
rect 154396 444372 154448 444378
rect 154396 444314 154448 444320
rect 137836 437436 137888 437442
rect 137836 437378 137888 437384
rect 154396 437436 154448 437442
rect 154396 437378 154448 437384
rect 137848 434738 137876 437378
rect 154408 434738 154436 437378
rect 137848 434710 137968 434738
rect 154408 434710 154528 434738
rect 137940 425134 137968 434710
rect 154500 425134 154528 434710
rect 137744 425128 137796 425134
rect 137744 425070 137796 425076
rect 137928 425128 137980 425134
rect 137928 425070 137980 425076
rect 154304 425128 154356 425134
rect 154304 425070 154356 425076
rect 154488 425128 154540 425134
rect 154488 425070 154540 425076
rect 123208 424584 123260 424590
rect 123208 424526 123260 424532
rect 111432 424516 111484 424522
rect 111432 424458 111484 424464
rect 99656 424448 99708 424454
rect 99656 424390 99708 424396
rect 106188 424448 106240 424454
rect 106188 424390 106240 424396
rect 87880 424380 87932 424386
rect 87880 424322 87932 424328
rect 89628 424380 89680 424386
rect 89628 424322 89680 424328
rect 87892 422348 87920 424322
rect 99668 422348 99696 424390
rect 111444 422348 111472 424458
rect 123220 422348 123248 424526
rect 137756 424386 137784 425070
rect 154316 424454 154344 425070
rect 146760 424448 146812 424454
rect 146760 424390 146812 424396
rect 154304 424448 154356 424454
rect 154304 424390 154356 424396
rect 170404 424448 170456 424454
rect 170404 424390 170456 424396
rect 134984 424380 135036 424386
rect 134984 424322 135036 424328
rect 137744 424380 137796 424386
rect 137744 424322 137796 424328
rect 134996 422348 135024 424322
rect 146772 422348 146800 424390
rect 158536 424380 158588 424386
rect 158536 424322 158588 424328
rect 158548 422348 158576 424322
rect 170416 422348 170444 424390
rect 171060 424386 171088 700198
rect 202800 697610 202828 703520
rect 218992 703474 219020 703520
rect 235184 703474 235212 703520
rect 218992 703446 219112 703474
rect 235184 703446 235304 703474
rect 201500 697604 201552 697610
rect 201500 697546 201552 697552
rect 202788 697604 202840 697610
rect 202788 697546 202840 697552
rect 171048 424380 171100 424386
rect 171048 424322 171100 424328
rect 182180 424380 182232 424386
rect 182180 424322 182232 424328
rect 182192 422348 182220 424322
rect 201512 423706 201540 697546
rect 219084 692850 219112 703446
rect 235276 692850 235304 703446
rect 267660 697610 267688 703520
rect 283852 703474 283880 703520
rect 283852 703446 283972 703474
rect 283944 698290 283972 703446
rect 283288 698284 283340 698290
rect 283288 698226 283340 698232
rect 283932 698284 283984 698290
rect 283932 698226 283984 698232
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 218060 692844 218112 692850
rect 218060 692786 218112 692792
rect 219072 692844 219124 692850
rect 219072 692786 219124 692792
rect 234620 692844 234672 692850
rect 234620 692786 234672 692792
rect 235264 692844 235316 692850
rect 235264 692786 235316 692792
rect 218072 683074 218100 692786
rect 234632 683074 234660 692786
rect 218072 683046 218284 683074
rect 234632 683046 234844 683074
rect 218256 673538 218284 683046
rect 234816 673538 234844 683046
rect 218060 673532 218112 673538
rect 218060 673474 218112 673480
rect 218244 673532 218296 673538
rect 218244 673474 218296 673480
rect 234620 673532 234672 673538
rect 234620 673474 234672 673480
rect 234804 673532 234856 673538
rect 234804 673474 234856 673480
rect 218072 663762 218100 673474
rect 234632 663762 234660 673474
rect 218072 663734 218284 663762
rect 234632 663734 234844 663762
rect 218256 654158 218284 663734
rect 234816 654158 234844 663734
rect 218060 654152 218112 654158
rect 218060 654094 218112 654100
rect 218244 654152 218296 654158
rect 218244 654094 218296 654100
rect 234620 654152 234672 654158
rect 234620 654094 234672 654100
rect 234804 654152 234856 654158
rect 234804 654094 234856 654100
rect 218072 644450 218100 654094
rect 234632 644450 234660 654094
rect 218072 644422 218284 644450
rect 234632 644422 234844 644450
rect 218256 634846 218284 644422
rect 234816 634846 234844 644422
rect 218060 634840 218112 634846
rect 218060 634782 218112 634788
rect 218244 634840 218296 634846
rect 218244 634782 218296 634788
rect 234620 634840 234672 634846
rect 234620 634782 234672 634788
rect 234804 634840 234856 634846
rect 234804 634782 234856 634788
rect 218072 625138 218100 634782
rect 234632 625138 234660 634782
rect 218072 625110 218284 625138
rect 234632 625110 234844 625138
rect 218256 615534 218284 625110
rect 234816 615534 234844 625110
rect 218060 615528 218112 615534
rect 218060 615470 218112 615476
rect 218244 615528 218296 615534
rect 218244 615470 218296 615476
rect 234620 615528 234672 615534
rect 234620 615470 234672 615476
rect 234804 615528 234856 615534
rect 234804 615470 234856 615476
rect 218072 605826 218100 615470
rect 234632 605826 234660 615470
rect 218072 605798 218284 605826
rect 234632 605798 234844 605826
rect 218256 596222 218284 605798
rect 234816 596222 234844 605798
rect 218060 596216 218112 596222
rect 218244 596216 218296 596222
rect 218112 596164 218192 596170
rect 218060 596158 218192 596164
rect 218244 596158 218296 596164
rect 234620 596216 234672 596222
rect 234804 596216 234856 596222
rect 234672 596164 234752 596170
rect 234620 596158 234752 596164
rect 234804 596158 234856 596164
rect 218072 596142 218192 596158
rect 234632 596142 234752 596158
rect 218164 596034 218192 596142
rect 234724 596034 234752 596142
rect 218164 596006 218284 596034
rect 234724 596006 234844 596034
rect 218256 591954 218284 596006
rect 234816 591954 234844 596006
rect 218164 591926 218284 591954
rect 234724 591926 234844 591954
rect 218164 589286 218192 591926
rect 234724 589286 234752 591926
rect 218152 589280 218204 589286
rect 218152 589222 218204 589228
rect 234712 589280 234764 589286
rect 234712 589222 234764 589228
rect 218060 579692 218112 579698
rect 218060 579634 218112 579640
rect 234620 579692 234672 579698
rect 234620 579634 234672 579640
rect 218072 572642 218100 579634
rect 234632 572642 234660 579634
rect 218072 572614 218192 572642
rect 234632 572614 234752 572642
rect 218164 569906 218192 572614
rect 234724 569906 234752 572614
rect 218152 569900 218204 569906
rect 218152 569842 218204 569848
rect 234712 569900 234764 569906
rect 234712 569842 234764 569848
rect 218336 563100 218388 563106
rect 218336 563042 218388 563048
rect 234896 563100 234948 563106
rect 234896 563042 234948 563048
rect 218348 560289 218376 563042
rect 234908 560289 234936 563042
rect 218150 560280 218206 560289
rect 218150 560215 218206 560224
rect 218334 560280 218390 560289
rect 218334 560215 218390 560224
rect 234710 560280 234766 560289
rect 234710 560215 234766 560224
rect 234894 560280 234950 560289
rect 234894 560215 234950 560224
rect 218164 550662 218192 560215
rect 234724 550662 234752 560215
rect 218152 550656 218204 550662
rect 218152 550598 218204 550604
rect 218428 550656 218480 550662
rect 218428 550598 218480 550604
rect 234712 550656 234764 550662
rect 234712 550598 234764 550604
rect 234988 550656 235040 550662
rect 234988 550598 235040 550604
rect 218440 543862 218468 550598
rect 235000 543862 235028 550598
rect 218428 543856 218480 543862
rect 218428 543798 218480 543804
rect 234988 543856 235040 543862
rect 234988 543798 235040 543804
rect 218336 543720 218388 543726
rect 218336 543662 218388 543668
rect 234896 543720 234948 543726
rect 234896 543662 234948 543668
rect 218348 540977 218376 543662
rect 234908 540977 234936 543662
rect 218150 540968 218206 540977
rect 218150 540903 218206 540912
rect 218334 540968 218390 540977
rect 218334 540903 218390 540912
rect 234710 540968 234766 540977
rect 234710 540903 234766 540912
rect 234894 540968 234950 540977
rect 234894 540903 234950 540912
rect 218164 531350 218192 540903
rect 234724 531350 234752 540903
rect 218152 531344 218204 531350
rect 218152 531286 218204 531292
rect 218428 531344 218480 531350
rect 218428 531286 218480 531292
rect 234712 531344 234764 531350
rect 234712 531286 234764 531292
rect 234988 531344 235040 531350
rect 234988 531286 235040 531292
rect 218440 524550 218468 531286
rect 235000 524550 235028 531286
rect 218428 524544 218480 524550
rect 218428 524486 218480 524492
rect 234988 524544 235040 524550
rect 234988 524486 235040 524492
rect 218336 524408 218388 524414
rect 218336 524350 218388 524356
rect 234896 524408 234948 524414
rect 234896 524350 234948 524356
rect 218348 521665 218376 524350
rect 234908 521665 234936 524350
rect 218150 521656 218206 521665
rect 218150 521591 218206 521600
rect 218334 521656 218390 521665
rect 218334 521591 218390 521600
rect 234710 521656 234766 521665
rect 234710 521591 234766 521600
rect 234894 521656 234950 521665
rect 234894 521591 234950 521600
rect 218164 512038 218192 521591
rect 234724 512038 234752 521591
rect 218152 512032 218204 512038
rect 218152 511974 218204 511980
rect 218428 512032 218480 512038
rect 218428 511974 218480 511980
rect 234712 512032 234764 512038
rect 234712 511974 234764 511980
rect 234988 512032 235040 512038
rect 234988 511974 235040 511980
rect 218440 502382 218468 511974
rect 235000 502382 235028 511974
rect 218244 502376 218296 502382
rect 217966 502344 218022 502353
rect 217966 502279 218022 502288
rect 218242 502344 218244 502353
rect 218428 502376 218480 502382
rect 218296 502344 218298 502353
rect 234804 502376 234856 502382
rect 218428 502318 218480 502324
rect 234526 502344 234582 502353
rect 218242 502279 218298 502288
rect 234526 502279 234582 502288
rect 234802 502344 234804 502353
rect 234988 502376 235040 502382
rect 234856 502344 234858 502353
rect 234988 502318 235040 502324
rect 234802 502279 234858 502288
rect 217980 492697 218008 502279
rect 234540 492697 234568 502279
rect 217966 492688 218022 492697
rect 217966 492623 218022 492632
rect 218150 492688 218206 492697
rect 218150 492623 218206 492632
rect 234526 492688 234582 492697
rect 234526 492623 234582 492632
rect 234710 492688 234766 492697
rect 234710 492623 234766 492632
rect 218164 489954 218192 492623
rect 234724 489954 234752 492623
rect 218164 489926 218284 489954
rect 234724 489926 234844 489954
rect 218256 480282 218284 489926
rect 234816 480282 234844 489926
rect 218060 480276 218112 480282
rect 218060 480218 218112 480224
rect 218244 480276 218296 480282
rect 218244 480218 218296 480224
rect 234620 480276 234672 480282
rect 234620 480218 234672 480224
rect 234804 480276 234856 480282
rect 234804 480218 234856 480224
rect 218072 480162 218100 480218
rect 234632 480162 234660 480218
rect 218072 480134 218192 480162
rect 234632 480134 234752 480162
rect 218164 470642 218192 480134
rect 234724 470642 234752 480134
rect 218164 470614 218284 470642
rect 234724 470614 234844 470642
rect 218256 460970 218284 470614
rect 234816 460970 234844 470614
rect 218060 460964 218112 460970
rect 218060 460906 218112 460912
rect 218244 460964 218296 460970
rect 218244 460906 218296 460912
rect 234620 460964 234672 460970
rect 234620 460906 234672 460912
rect 234804 460964 234856 460970
rect 234804 460906 234856 460912
rect 218072 460850 218100 460906
rect 234632 460850 234660 460906
rect 218072 460822 218192 460850
rect 234632 460822 234752 460850
rect 218164 451330 218192 460822
rect 234724 451330 234752 460822
rect 218164 451302 218284 451330
rect 234724 451302 234844 451330
rect 218256 441658 218284 451302
rect 234816 441658 234844 451302
rect 218060 441652 218112 441658
rect 218060 441594 218112 441600
rect 218244 441652 218296 441658
rect 218244 441594 218296 441600
rect 234620 441652 234672 441658
rect 234620 441594 234672 441600
rect 234804 441652 234856 441658
rect 234804 441594 234856 441600
rect 218072 441538 218100 441594
rect 234632 441538 234660 441594
rect 218072 441510 218192 441538
rect 234632 441510 234752 441538
rect 218164 432018 218192 441510
rect 234724 432018 234752 441510
rect 218164 431990 218284 432018
rect 234724 431990 234844 432018
rect 218256 424454 218284 431990
rect 205732 424448 205784 424454
rect 205732 424390 205784 424396
rect 218244 424448 218296 424454
rect 218244 424390 218296 424396
rect 229284 424448 229336 424454
rect 229284 424390 229336 424396
rect 193956 423700 194008 423706
rect 193956 423642 194008 423648
rect 201500 423700 201552 423706
rect 201500 423642 201552 423648
rect 193968 422348 193996 423642
rect 205744 422348 205772 424390
rect 217508 424380 217560 424386
rect 217508 424322 217560 424328
rect 217520 422348 217548 424322
rect 229296 422348 229324 424390
rect 234816 424386 234844 431990
rect 252928 424584 252980 424590
rect 252928 424526 252980 424532
rect 234804 424380 234856 424386
rect 234804 424322 234856 424328
rect 241060 424380 241112 424386
rect 241060 424322 241112 424328
rect 241072 422348 241100 424322
rect 252940 422348 252968 424526
rect 264704 424516 264756 424522
rect 264704 424458 264756 424464
rect 264716 422348 264744 424458
rect 266372 424454 266400 697546
rect 283300 694142 283328 698226
rect 283104 694136 283156 694142
rect 283104 694078 283156 694084
rect 283288 694136 283340 694142
rect 283288 694078 283340 694084
rect 283116 692782 283144 694078
rect 283104 692776 283156 692782
rect 283104 692718 283156 692724
rect 283288 692776 283340 692782
rect 283288 692718 283340 692724
rect 283300 683233 283328 692718
rect 300136 684486 300164 703520
rect 332520 697610 332548 703520
rect 348804 703474 348832 703520
rect 364996 703474 365024 703520
rect 348804 703446 348924 703474
rect 364996 703446 365116 703474
rect 331220 697604 331272 697610
rect 331220 697546 331272 697552
rect 332508 697604 332560 697610
rect 332508 697546 332560 697552
rect 299480 684480 299532 684486
rect 299480 684422 299532 684428
rect 300124 684480 300176 684486
rect 300124 684422 300176 684428
rect 282918 683224 282974 683233
rect 282918 683159 282974 683168
rect 283286 683224 283342 683233
rect 283286 683159 283342 683168
rect 282932 683126 282960 683159
rect 299492 683126 299520 684422
rect 282920 683120 282972 683126
rect 282920 683062 282972 683068
rect 299480 683120 299532 683126
rect 299480 683062 299532 683068
rect 283380 666596 283432 666602
rect 283380 666538 283432 666544
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 283392 659682 283420 666538
rect 299952 659682 299980 666538
rect 283208 659654 283420 659682
rect 299768 659654 299980 659682
rect 283208 647290 283236 659654
rect 299768 647290 299796 659654
rect 283104 647284 283156 647290
rect 283104 647226 283156 647232
rect 283196 647284 283248 647290
rect 283196 647226 283248 647232
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 283116 640422 283144 647226
rect 299676 640422 299704 647226
rect 283104 640416 283156 640422
rect 283104 640358 283156 640364
rect 283196 640416 283248 640422
rect 283196 640358 283248 640364
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 283208 630698 283236 640358
rect 299768 630698 299796 640358
rect 283012 630692 283064 630698
rect 283012 630634 283064 630640
rect 283196 630692 283248 630698
rect 283196 630634 283248 630640
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 283024 630578 283052 630634
rect 299584 630578 299612 630634
rect 283024 630550 283144 630578
rect 299584 630550 299704 630578
rect 283116 621058 283144 630550
rect 299676 621058 299704 630550
rect 283116 621030 283236 621058
rect 299676 621030 299796 621058
rect 283208 611386 283236 621030
rect 299768 611386 299796 621030
rect 283012 611380 283064 611386
rect 283012 611322 283064 611328
rect 283196 611380 283248 611386
rect 283196 611322 283248 611328
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 283024 611266 283052 611322
rect 299584 611266 299612 611322
rect 283024 611238 283144 611266
rect 299584 611238 299704 611266
rect 283116 608598 283144 611238
rect 299676 608598 299704 611238
rect 283104 608592 283156 608598
rect 283104 608534 283156 608540
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 283288 601724 283340 601730
rect 283288 601666 283340 601672
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 283300 598942 283328 601666
rect 299860 598942 299888 601666
rect 283288 598936 283340 598942
rect 283288 598878 283340 598884
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 283380 589348 283432 589354
rect 283380 589290 283432 589296
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 283392 582486 283420 589290
rect 299952 582486 299980 589290
rect 283380 582480 283432 582486
rect 283380 582422 283432 582428
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 283288 582344 283340 582350
rect 283288 582286 283340 582292
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 283300 572642 283328 582286
rect 299860 572642 299888 582286
rect 283116 572614 283328 572642
rect 299676 572614 299888 572642
rect 283116 569922 283144 572614
rect 299676 569945 299704 572614
rect 283024 569894 283144 569922
rect 299662 569936 299718 569945
rect 283024 563174 283052 569894
rect 299662 569871 299718 569880
rect 283012 563168 283064 563174
rect 283012 563110 283064 563116
rect 283012 563032 283064 563038
rect 283012 562974 283064 562980
rect 283024 560250 283052 562974
rect 299570 560416 299626 560425
rect 299570 560351 299626 560360
rect 299584 560289 299612 560351
rect 299570 560280 299626 560289
rect 283012 560244 283064 560250
rect 299570 560215 299626 560224
rect 299754 560280 299810 560289
rect 299754 560215 299810 560224
rect 283012 560186 283064 560192
rect 299768 550662 299796 560215
rect 283196 550656 283248 550662
rect 283196 550598 283248 550604
rect 299480 550656 299532 550662
rect 299480 550598 299532 550604
rect 299756 550656 299808 550662
rect 299756 550598 299808 550604
rect 283208 543658 283236 550598
rect 299492 543794 299520 550598
rect 299480 543788 299532 543794
rect 299480 543730 299532 543736
rect 283012 543652 283064 543658
rect 283012 543594 283064 543600
rect 283196 543652 283248 543658
rect 283196 543594 283248 543600
rect 299572 543652 299624 543658
rect 299572 543594 299624 543600
rect 283024 534070 283052 543594
rect 299584 534070 299612 543594
rect 283012 534064 283064 534070
rect 283012 534006 283064 534012
rect 283196 534064 283248 534070
rect 283196 534006 283248 534012
rect 299572 534064 299624 534070
rect 299572 534006 299624 534012
rect 299756 534064 299808 534070
rect 299756 534006 299808 534012
rect 283208 524482 283236 534006
rect 299768 524482 299796 534006
rect 283196 524476 283248 524482
rect 283196 524418 283248 524424
rect 299756 524476 299808 524482
rect 299756 524418 299808 524424
rect 283288 524408 283340 524414
rect 283288 524350 283340 524356
rect 299848 524408 299900 524414
rect 299848 524350 299900 524356
rect 283300 521665 283328 524350
rect 299860 521665 299888 524350
rect 283102 521656 283158 521665
rect 283102 521591 283158 521600
rect 283286 521656 283342 521665
rect 283286 521591 283342 521600
rect 299662 521656 299718 521665
rect 299662 521591 299718 521600
rect 299846 521656 299902 521665
rect 299846 521591 299902 521600
rect 283116 512038 283144 521591
rect 299676 512038 299704 521591
rect 283104 512032 283156 512038
rect 283104 511974 283156 511980
rect 283380 512032 283432 512038
rect 283380 511974 283432 511980
rect 299664 512032 299716 512038
rect 299664 511974 299716 511980
rect 299940 512032 299992 512038
rect 299940 511974 299992 511980
rect 283392 502382 283420 511974
rect 299952 502382 299980 511974
rect 283196 502376 283248 502382
rect 282918 502344 282974 502353
rect 282918 502279 282974 502288
rect 283194 502344 283196 502353
rect 283380 502376 283432 502382
rect 283248 502344 283250 502353
rect 299756 502376 299808 502382
rect 283380 502318 283432 502324
rect 299478 502344 299534 502353
rect 283194 502279 283250 502288
rect 299478 502279 299534 502288
rect 299754 502344 299756 502353
rect 299940 502376 299992 502382
rect 299808 502344 299810 502353
rect 299940 502318 299992 502324
rect 299754 502279 299810 502288
rect 282932 492697 282960 502279
rect 299492 492697 299520 502279
rect 282918 492688 282974 492697
rect 282918 492623 282974 492632
rect 283102 492688 283158 492697
rect 283102 492623 283104 492632
rect 283156 492623 283158 492632
rect 299478 492688 299534 492697
rect 299478 492623 299534 492632
rect 299662 492688 299718 492697
rect 299662 492623 299664 492632
rect 283104 492594 283156 492600
rect 299716 492623 299718 492632
rect 299664 492594 299716 492600
rect 283104 485784 283156 485790
rect 283104 485726 283156 485732
rect 299664 485784 299716 485790
rect 299664 485726 299716 485732
rect 283116 483018 283144 485726
rect 299676 483018 299704 485726
rect 283116 482990 283236 483018
rect 299676 482990 299796 483018
rect 283208 476134 283236 482990
rect 299768 476134 299796 482990
rect 283012 476128 283064 476134
rect 283196 476128 283248 476134
rect 283064 476076 283144 476082
rect 283012 476070 283144 476076
rect 283196 476070 283248 476076
rect 299572 476128 299624 476134
rect 299756 476128 299808 476134
rect 299624 476076 299704 476082
rect 299572 476070 299704 476076
rect 299756 476070 299808 476076
rect 283024 476054 283144 476070
rect 299584 476054 299704 476070
rect 283116 473346 283144 476054
rect 299676 473346 299704 476054
rect 283104 473340 283156 473346
rect 283104 473282 283156 473288
rect 299664 473340 299716 473346
rect 299664 473282 299716 473288
rect 283104 466404 283156 466410
rect 283104 466346 283156 466352
rect 299664 466404 299716 466410
rect 299664 466346 299716 466352
rect 283116 463706 283144 466346
rect 299676 463706 299704 466346
rect 283116 463678 283236 463706
rect 299676 463678 299796 463706
rect 283208 454073 283236 463678
rect 282918 454064 282974 454073
rect 282918 453999 282974 454008
rect 283194 454064 283250 454073
rect 299768 454050 299796 463678
rect 283194 453999 283250 454008
rect 299584 454022 299796 454050
rect 282932 447166 282960 453999
rect 299584 453966 299612 454022
rect 299572 453960 299624 453966
rect 299572 453902 299624 453908
rect 282920 447160 282972 447166
rect 282920 447102 282972 447108
rect 283012 447092 283064 447098
rect 283012 447034 283064 447040
rect 299572 447092 299624 447098
rect 299572 447034 299624 447040
rect 283024 437458 283052 447034
rect 299584 437458 299612 447034
rect 283024 437430 283144 437458
rect 299584 437430 299704 437458
rect 283116 434722 283144 437430
rect 299676 434722 299704 437430
rect 283104 434716 283156 434722
rect 283104 434658 283156 434664
rect 299664 434716 299716 434722
rect 299664 434658 299716 434664
rect 283104 427780 283156 427786
rect 283104 427722 283156 427728
rect 299664 427780 299716 427786
rect 299664 427722 299716 427728
rect 283116 425082 283144 427722
rect 299676 425082 299704 427722
rect 283116 425054 283236 425082
rect 299676 425054 299796 425082
rect 266360 424448 266412 424454
rect 266360 424390 266412 424396
rect 276480 424448 276532 424454
rect 276480 424390 276532 424396
rect 276492 422348 276520 424390
rect 283208 424386 283236 425054
rect 299768 424590 299796 425054
rect 300032 424924 300084 424930
rect 300032 424866 300084 424872
rect 299756 424584 299808 424590
rect 299756 424526 299808 424532
rect 283196 424380 283248 424386
rect 283196 424322 283248 424328
rect 288256 424380 288308 424386
rect 288256 424322 288308 424328
rect 288268 422348 288296 424322
rect 300044 422348 300072 424866
rect 311808 424856 311860 424862
rect 311808 424798 311860 424804
rect 311820 422348 311848 424798
rect 323584 424788 323636 424794
rect 323584 424730 323636 424736
rect 323596 422348 323624 424730
rect 331232 424522 331260 697546
rect 348896 692850 348924 703446
rect 365088 692850 365116 703446
rect 347780 692844 347832 692850
rect 347780 692786 347832 692792
rect 348884 692844 348936 692850
rect 348884 692786 348936 692792
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 347792 683074 347820 692786
rect 364352 683074 364380 692786
rect 347792 683046 348004 683074
rect 364352 683046 364564 683074
rect 347976 673538 348004 683046
rect 364536 673538 364564 683046
rect 347780 673532 347832 673538
rect 347780 673474 347832 673480
rect 347964 673532 348016 673538
rect 347964 673474 348016 673480
rect 364340 673532 364392 673538
rect 364340 673474 364392 673480
rect 364524 673532 364576 673538
rect 364524 673474 364576 673480
rect 347792 663762 347820 673474
rect 364352 663762 364380 673474
rect 347792 663734 348004 663762
rect 364352 663734 364564 663762
rect 347976 654158 348004 663734
rect 364536 654158 364564 663734
rect 347780 654152 347832 654158
rect 347780 654094 347832 654100
rect 347964 654152 348016 654158
rect 347964 654094 348016 654100
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 347792 644450 347820 654094
rect 364352 644450 364380 654094
rect 347792 644422 348004 644450
rect 364352 644422 364564 644450
rect 347976 634846 348004 644422
rect 364536 634846 364564 644422
rect 347780 634840 347832 634846
rect 347780 634782 347832 634788
rect 347964 634840 348016 634846
rect 347964 634782 348016 634788
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 347792 625138 347820 634782
rect 364352 625138 364380 634782
rect 347792 625110 348004 625138
rect 364352 625110 364564 625138
rect 347976 615534 348004 625110
rect 364536 615534 364564 625110
rect 347780 615528 347832 615534
rect 347780 615470 347832 615476
rect 347964 615528 348016 615534
rect 347964 615470 348016 615476
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 347792 605826 347820 615470
rect 364352 605826 364380 615470
rect 347792 605798 348004 605826
rect 364352 605798 364564 605826
rect 347976 596222 348004 605798
rect 364536 596222 364564 605798
rect 347780 596216 347832 596222
rect 347964 596216 348016 596222
rect 347832 596164 347912 596170
rect 347780 596158 347912 596164
rect 347964 596158 348016 596164
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 347792 596142 347912 596158
rect 364352 596142 364472 596158
rect 347884 596034 347912 596142
rect 364444 596034 364472 596142
rect 347884 596006 348004 596034
rect 364444 596006 364564 596034
rect 347976 591954 348004 596006
rect 364536 591954 364564 596006
rect 347884 591926 348004 591954
rect 364444 591926 364564 591954
rect 347884 589286 347912 591926
rect 364444 589286 364472 591926
rect 347872 589280 347924 589286
rect 347872 589222 347924 589228
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 347780 579692 347832 579698
rect 347780 579634 347832 579640
rect 364340 579692 364392 579698
rect 364340 579634 364392 579640
rect 347792 572642 347820 579634
rect 364352 572642 364380 579634
rect 347792 572614 347912 572642
rect 364352 572614 364472 572642
rect 347884 569906 347912 572614
rect 364444 569906 364472 572614
rect 347872 569900 347924 569906
rect 347872 569842 347924 569848
rect 364432 569900 364484 569906
rect 364432 569842 364484 569848
rect 348056 563100 348108 563106
rect 348056 563042 348108 563048
rect 364616 563100 364668 563106
rect 364616 563042 364668 563048
rect 348068 560289 348096 563042
rect 364628 560289 364656 563042
rect 347870 560280 347926 560289
rect 347870 560215 347926 560224
rect 348054 560280 348110 560289
rect 348054 560215 348110 560224
rect 364430 560280 364486 560289
rect 364430 560215 364486 560224
rect 364614 560280 364670 560289
rect 364614 560215 364670 560224
rect 347884 550662 347912 560215
rect 364444 550662 364472 560215
rect 347872 550656 347924 550662
rect 347872 550598 347924 550604
rect 348148 550656 348200 550662
rect 348148 550598 348200 550604
rect 364432 550656 364484 550662
rect 364432 550598 364484 550604
rect 364708 550656 364760 550662
rect 364708 550598 364760 550604
rect 348160 543862 348188 550598
rect 364720 543862 364748 550598
rect 348148 543856 348200 543862
rect 348148 543798 348200 543804
rect 364708 543856 364760 543862
rect 364708 543798 364760 543804
rect 348056 543720 348108 543726
rect 348056 543662 348108 543668
rect 364616 543720 364668 543726
rect 364616 543662 364668 543668
rect 348068 540977 348096 543662
rect 364628 540977 364656 543662
rect 347870 540968 347926 540977
rect 347870 540903 347926 540912
rect 348054 540968 348110 540977
rect 348054 540903 348110 540912
rect 364430 540968 364486 540977
rect 364430 540903 364486 540912
rect 364614 540968 364670 540977
rect 364614 540903 364670 540912
rect 347884 531350 347912 540903
rect 364444 531350 364472 540903
rect 347872 531344 347924 531350
rect 347872 531286 347924 531292
rect 348148 531344 348200 531350
rect 348148 531286 348200 531292
rect 364432 531344 364484 531350
rect 364432 531286 364484 531292
rect 364708 531344 364760 531350
rect 364708 531286 364760 531292
rect 348160 524550 348188 531286
rect 364720 524550 364748 531286
rect 348148 524544 348200 524550
rect 348148 524486 348200 524492
rect 364708 524544 364760 524550
rect 364708 524486 364760 524492
rect 348056 524408 348108 524414
rect 348056 524350 348108 524356
rect 364616 524408 364668 524414
rect 364616 524350 364668 524356
rect 348068 521665 348096 524350
rect 364628 521665 364656 524350
rect 347870 521656 347926 521665
rect 347870 521591 347926 521600
rect 348054 521656 348110 521665
rect 348054 521591 348110 521600
rect 364430 521656 364486 521665
rect 364430 521591 364486 521600
rect 364614 521656 364670 521665
rect 364614 521591 364670 521600
rect 347884 512038 347912 521591
rect 364444 512038 364472 521591
rect 347872 512032 347924 512038
rect 347872 511974 347924 511980
rect 348148 512032 348200 512038
rect 348148 511974 348200 511980
rect 364432 512032 364484 512038
rect 364432 511974 364484 511980
rect 364708 512032 364760 512038
rect 364708 511974 364760 511980
rect 348160 502382 348188 511974
rect 364720 502382 364748 511974
rect 347964 502376 348016 502382
rect 347962 502344 347964 502353
rect 348148 502376 348200 502382
rect 348016 502344 348018 502353
rect 364524 502376 364576 502382
rect 348148 502318 348200 502324
rect 364246 502344 364302 502353
rect 347962 502279 348018 502288
rect 364246 502279 364302 502288
rect 364522 502344 364524 502353
rect 364708 502376 364760 502382
rect 364576 502344 364578 502353
rect 364708 502318 364760 502324
rect 364522 502279 364578 502288
rect 364260 492697 364288 502279
rect 347870 492688 347926 492697
rect 347870 492623 347926 492632
rect 364246 492688 364302 492697
rect 364246 492623 364302 492632
rect 364430 492688 364486 492697
rect 364430 492623 364486 492632
rect 347884 489954 347912 492623
rect 364444 489954 364472 492623
rect 347884 489926 348004 489954
rect 364444 489926 364564 489954
rect 347976 480282 348004 489926
rect 364536 480282 364564 489926
rect 347780 480276 347832 480282
rect 347780 480218 347832 480224
rect 347964 480276 348016 480282
rect 347964 480218 348016 480224
rect 364340 480276 364392 480282
rect 364340 480218 364392 480224
rect 364524 480276 364576 480282
rect 364524 480218 364576 480224
rect 347792 480162 347820 480218
rect 364352 480162 364380 480218
rect 347792 480134 347912 480162
rect 364352 480134 364472 480162
rect 347884 470642 347912 480134
rect 364444 470642 364472 480134
rect 347884 470614 348004 470642
rect 364444 470614 364564 470642
rect 347976 460970 348004 470614
rect 364536 460970 364564 470614
rect 347780 460964 347832 460970
rect 347780 460906 347832 460912
rect 347964 460964 348016 460970
rect 347964 460906 348016 460912
rect 364340 460964 364392 460970
rect 364340 460906 364392 460912
rect 364524 460964 364576 460970
rect 364524 460906 364576 460912
rect 347792 460850 347820 460906
rect 364352 460850 364380 460906
rect 347792 460822 347912 460850
rect 364352 460822 364472 460850
rect 347884 451330 347912 460822
rect 364444 451330 364472 460822
rect 347884 451302 348004 451330
rect 364444 451302 364564 451330
rect 347976 441658 348004 451302
rect 364536 441658 364564 451302
rect 347780 441652 347832 441658
rect 347780 441594 347832 441600
rect 347964 441652 348016 441658
rect 347964 441594 348016 441600
rect 364340 441652 364392 441658
rect 364340 441594 364392 441600
rect 364524 441652 364576 441658
rect 364524 441594 364576 441600
rect 347792 441538 347820 441594
rect 364352 441538 364380 441594
rect 347792 441510 347912 441538
rect 364352 441510 364472 441538
rect 347884 432018 347912 441510
rect 364444 432018 364472 441510
rect 347884 431990 348004 432018
rect 364444 431990 364564 432018
rect 335452 424720 335504 424726
rect 335452 424662 335504 424668
rect 331220 424516 331272 424522
rect 331220 424458 331272 424464
rect 335464 422348 335492 424662
rect 347228 424652 347280 424658
rect 347228 424594 347280 424600
rect 347240 422348 347268 424594
rect 347976 424454 348004 431990
rect 359004 424584 359056 424590
rect 359004 424526 359056 424532
rect 347964 424448 348016 424454
rect 347964 424390 348016 424396
rect 359016 422348 359044 424526
rect 364536 424386 364564 431990
rect 397472 424930 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 413756 698290 413784 703446
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 429856 684486 429884 703520
rect 429200 684480 429252 684486
rect 429200 684422 429252 684428
rect 429844 684480 429896 684486
rect 429844 684422 429896 684428
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 429212 683126 429240 684422
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 429200 683120 429252 683126
rect 429200 683062 429252 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 413112 659682 413140 666538
rect 429672 659682 429700 666538
rect 412928 659654 413140 659682
rect 429488 659654 429700 659682
rect 412928 647290 412956 659654
rect 429488 647290 429516 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 412836 640422 412864 647226
rect 429396 640422 429424 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 412928 630698 412956 640358
rect 429488 630698 429516 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 412744 630578 412772 630634
rect 429304 630578 429332 630634
rect 412744 630550 412864 630578
rect 429304 630550 429424 630578
rect 412836 621058 412864 630550
rect 429396 621058 429424 630550
rect 412836 621030 412956 621058
rect 429396 621030 429516 621058
rect 412928 611386 412956 621030
rect 429488 611386 429516 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 412744 611266 412772 611322
rect 429304 611266 429332 611322
rect 412744 611238 412864 611266
rect 429304 611238 429424 611266
rect 412836 608598 412864 611238
rect 429396 608598 429424 611238
rect 412824 608592 412876 608598
rect 412824 608534 412876 608540
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 413008 601724 413060 601730
rect 413008 601666 413060 601672
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 413020 598942 413048 601666
rect 429580 598942 429608 601666
rect 413008 598936 413060 598942
rect 413008 598878 413060 598884
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 413100 589348 413152 589354
rect 413100 589290 413152 589296
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 413112 582486 413140 589290
rect 429672 582486 429700 589290
rect 413100 582480 413152 582486
rect 413100 582422 413152 582428
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 413008 582344 413060 582350
rect 413008 582286 413060 582292
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 413020 572642 413048 582286
rect 429580 572642 429608 582286
rect 412836 572614 413048 572642
rect 429396 572614 429608 572642
rect 412836 569922 412864 572614
rect 429396 569922 429424 572614
rect 412744 569894 412864 569922
rect 429304 569894 429424 569922
rect 412744 563174 412772 569894
rect 429304 563174 429332 569894
rect 412732 563168 412784 563174
rect 412732 563110 412784 563116
rect 429292 563168 429344 563174
rect 429292 563110 429344 563116
rect 412732 563032 412784 563038
rect 412732 562974 412784 562980
rect 429292 563032 429344 563038
rect 429292 562974 429344 562980
rect 412744 560250 412772 562974
rect 429304 560250 429332 562974
rect 412732 560244 412784 560250
rect 412732 560186 412784 560192
rect 429292 560244 429344 560250
rect 429292 560186 429344 560192
rect 412916 550656 412968 550662
rect 412916 550598 412968 550604
rect 429476 550656 429528 550662
rect 429476 550598 429528 550604
rect 412928 543658 412956 550598
rect 429488 543658 429516 550598
rect 412732 543652 412784 543658
rect 412732 543594 412784 543600
rect 412916 543652 412968 543658
rect 412916 543594 412968 543600
rect 429292 543652 429344 543658
rect 429292 543594 429344 543600
rect 429476 543652 429528 543658
rect 429476 543594 429528 543600
rect 412744 534070 412772 543594
rect 429304 534070 429332 543594
rect 412732 534064 412784 534070
rect 412732 534006 412784 534012
rect 412916 534064 412968 534070
rect 412916 534006 412968 534012
rect 429292 534064 429344 534070
rect 429292 534006 429344 534012
rect 429476 534064 429528 534070
rect 429476 534006 429528 534012
rect 412928 524482 412956 534006
rect 429488 524482 429516 534006
rect 412916 524476 412968 524482
rect 412916 524418 412968 524424
rect 429476 524476 429528 524482
rect 429476 524418 429528 524424
rect 413008 524408 413060 524414
rect 413008 524350 413060 524356
rect 429568 524408 429620 524414
rect 429568 524350 429620 524356
rect 413020 521665 413048 524350
rect 429580 521665 429608 524350
rect 412822 521656 412878 521665
rect 412822 521591 412878 521600
rect 413006 521656 413062 521665
rect 413006 521591 413062 521600
rect 429382 521656 429438 521665
rect 429382 521591 429438 521600
rect 429566 521656 429622 521665
rect 429566 521591 429622 521600
rect 412836 512038 412864 521591
rect 429396 512038 429424 521591
rect 412824 512032 412876 512038
rect 412824 511974 412876 511980
rect 413100 512032 413152 512038
rect 413100 511974 413152 511980
rect 429384 512032 429436 512038
rect 429384 511974 429436 511980
rect 429660 512032 429712 512038
rect 429660 511974 429712 511980
rect 413112 502382 413140 511974
rect 429672 502382 429700 511974
rect 412916 502376 412968 502382
rect 412638 502344 412694 502353
rect 412638 502279 412694 502288
rect 412914 502344 412916 502353
rect 413100 502376 413152 502382
rect 412968 502344 412970 502353
rect 429476 502376 429528 502382
rect 413100 502318 413152 502324
rect 429198 502344 429254 502353
rect 412914 502279 412970 502288
rect 429198 502279 429254 502288
rect 429474 502344 429476 502353
rect 429660 502376 429712 502382
rect 429528 502344 429530 502353
rect 429660 502318 429712 502324
rect 429474 502279 429530 502288
rect 412652 492697 412680 502279
rect 429212 492697 429240 502279
rect 412638 492688 412694 492697
rect 412638 492623 412694 492632
rect 412822 492688 412878 492697
rect 412822 492623 412824 492632
rect 412876 492623 412878 492632
rect 429198 492688 429254 492697
rect 429198 492623 429254 492632
rect 429382 492688 429438 492697
rect 429382 492623 429384 492632
rect 412824 492594 412876 492600
rect 429436 492623 429438 492632
rect 429384 492594 429436 492600
rect 412824 485784 412876 485790
rect 412824 485726 412876 485732
rect 429384 485784 429436 485790
rect 429384 485726 429436 485732
rect 412836 483018 412864 485726
rect 429396 483018 429424 485726
rect 412836 482990 412956 483018
rect 429396 482990 429516 483018
rect 412928 476134 412956 482990
rect 429488 476134 429516 482990
rect 412732 476128 412784 476134
rect 412916 476128 412968 476134
rect 412784 476076 412864 476082
rect 412732 476070 412864 476076
rect 412916 476070 412968 476076
rect 429292 476128 429344 476134
rect 429476 476128 429528 476134
rect 429344 476076 429424 476082
rect 429292 476070 429424 476076
rect 429476 476070 429528 476076
rect 412744 476054 412864 476070
rect 429304 476054 429424 476070
rect 412836 473346 412864 476054
rect 429396 473346 429424 476054
rect 412824 473340 412876 473346
rect 412824 473282 412876 473288
rect 429384 473340 429436 473346
rect 429384 473282 429436 473288
rect 412824 466404 412876 466410
rect 412824 466346 412876 466352
rect 429384 466404 429436 466410
rect 429384 466346 429436 466352
rect 412836 463706 412864 466346
rect 429396 463706 429424 466346
rect 412836 463678 412956 463706
rect 429396 463678 429516 463706
rect 412928 454073 412956 463678
rect 429488 454073 429516 463678
rect 412638 454064 412694 454073
rect 412638 453999 412694 454008
rect 412914 454064 412970 454073
rect 412914 453999 412970 454008
rect 429198 454064 429254 454073
rect 429198 453999 429254 454008
rect 429474 454064 429530 454073
rect 429474 453999 429530 454008
rect 412652 447166 412680 453999
rect 429212 447166 429240 453999
rect 412640 447160 412692 447166
rect 412640 447102 412692 447108
rect 429200 447160 429252 447166
rect 429200 447102 429252 447108
rect 412732 447092 412784 447098
rect 412732 447034 412784 447040
rect 429292 447092 429344 447098
rect 429292 447034 429344 447040
rect 412744 437458 412772 447034
rect 429304 437458 429332 447034
rect 412744 437430 412864 437458
rect 429304 437430 429424 437458
rect 412836 434722 412864 437430
rect 429396 434722 429424 437430
rect 412824 434716 412876 434722
rect 412824 434658 412876 434664
rect 429384 434716 429436 434722
rect 429384 434658 429436 434664
rect 412824 427780 412876 427786
rect 412824 427722 412876 427728
rect 429384 427780 429436 427786
rect 429384 427722 429436 427728
rect 412836 425082 412864 427722
rect 429396 425082 429424 427722
rect 412836 425054 412956 425082
rect 429396 425054 429516 425082
rect 397460 424924 397512 424930
rect 397460 424866 397512 424872
rect 412928 424862 412956 425054
rect 412916 424856 412968 424862
rect 412916 424798 412968 424804
rect 429488 424794 429516 425054
rect 429476 424788 429528 424794
rect 429476 424730 429528 424736
rect 462332 424726 462360 703520
rect 478524 703474 478552 703520
rect 494808 703474 494836 703520
rect 478524 703446 478644 703474
rect 494808 703446 494928 703474
rect 478616 692850 478644 703446
rect 494900 692850 494928 703446
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 477512 683074 477540 692786
rect 494072 683074 494100 692786
rect 477512 683046 477724 683074
rect 494072 683046 494284 683074
rect 477696 673538 477724 683046
rect 494256 673538 494284 683046
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 494060 673532 494112 673538
rect 494060 673474 494112 673480
rect 494244 673532 494296 673538
rect 494244 673474 494296 673480
rect 477512 663762 477540 673474
rect 494072 663762 494100 673474
rect 477512 663734 477724 663762
rect 494072 663734 494284 663762
rect 477696 654158 477724 663734
rect 494256 654158 494284 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 477512 644450 477540 654094
rect 494072 644450 494100 654094
rect 477512 644422 477724 644450
rect 494072 644422 494284 644450
rect 477696 634846 477724 644422
rect 494256 634846 494284 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 477512 625138 477540 634782
rect 494072 625138 494100 634782
rect 477512 625110 477724 625138
rect 494072 625110 494284 625138
rect 477696 615534 477724 625110
rect 494256 615534 494284 625110
rect 477500 615528 477552 615534
rect 477500 615470 477552 615476
rect 477684 615528 477736 615534
rect 477684 615470 477736 615476
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 477512 605826 477540 615470
rect 494072 605826 494100 615470
rect 477512 605798 477724 605826
rect 494072 605798 494284 605826
rect 477696 596222 477724 605798
rect 494256 596222 494284 605798
rect 477500 596216 477552 596222
rect 477684 596216 477736 596222
rect 477552 596164 477632 596170
rect 477500 596158 477632 596164
rect 477684 596158 477736 596164
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 477512 596142 477632 596158
rect 494072 596142 494192 596158
rect 477604 596034 477632 596142
rect 494164 596034 494192 596142
rect 477604 596006 477724 596034
rect 494164 596006 494284 596034
rect 477696 591954 477724 596006
rect 494256 591954 494284 596006
rect 477604 591926 477724 591954
rect 494164 591926 494284 591954
rect 477604 589286 477632 591926
rect 494164 589286 494192 591926
rect 477592 589280 477644 589286
rect 477592 589222 477644 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 477500 579692 477552 579698
rect 477500 579634 477552 579640
rect 494060 579692 494112 579698
rect 494060 579634 494112 579640
rect 477512 572642 477540 579634
rect 494072 572642 494100 579634
rect 477512 572614 477632 572642
rect 494072 572614 494192 572642
rect 477604 569906 477632 572614
rect 494164 569906 494192 572614
rect 477592 569900 477644 569906
rect 477592 569842 477644 569848
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 477776 563100 477828 563106
rect 477776 563042 477828 563048
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 477788 560289 477816 563042
rect 494348 560289 494376 563042
rect 477590 560280 477646 560289
rect 477590 560215 477646 560224
rect 477774 560280 477830 560289
rect 477774 560215 477830 560224
rect 494150 560280 494206 560289
rect 494150 560215 494206 560224
rect 494334 560280 494390 560289
rect 494334 560215 494390 560224
rect 477604 550662 477632 560215
rect 494164 550662 494192 560215
rect 477592 550656 477644 550662
rect 477592 550598 477644 550604
rect 477868 550656 477920 550662
rect 477868 550598 477920 550604
rect 494152 550656 494204 550662
rect 494152 550598 494204 550604
rect 494428 550656 494480 550662
rect 494428 550598 494480 550604
rect 477880 543862 477908 550598
rect 494440 543862 494468 550598
rect 477868 543856 477920 543862
rect 477868 543798 477920 543804
rect 494428 543856 494480 543862
rect 494428 543798 494480 543804
rect 477776 543720 477828 543726
rect 477776 543662 477828 543668
rect 494336 543720 494388 543726
rect 494336 543662 494388 543668
rect 477788 540977 477816 543662
rect 494348 540977 494376 543662
rect 477590 540968 477646 540977
rect 477590 540903 477646 540912
rect 477774 540968 477830 540977
rect 477774 540903 477830 540912
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 477604 531350 477632 540903
rect 494164 531350 494192 540903
rect 477592 531344 477644 531350
rect 477592 531286 477644 531292
rect 477868 531344 477920 531350
rect 477868 531286 477920 531292
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 477880 524550 477908 531286
rect 494440 524550 494468 531286
rect 477868 524544 477920 524550
rect 477868 524486 477920 524492
rect 494428 524544 494480 524550
rect 494428 524486 494480 524492
rect 477776 524408 477828 524414
rect 477776 524350 477828 524356
rect 494336 524408 494388 524414
rect 494336 524350 494388 524356
rect 477788 521665 477816 524350
rect 494348 521665 494376 524350
rect 477590 521656 477646 521665
rect 477590 521591 477646 521600
rect 477774 521656 477830 521665
rect 477774 521591 477830 521600
rect 494150 521656 494206 521665
rect 494150 521591 494206 521600
rect 494334 521656 494390 521665
rect 494334 521591 494390 521600
rect 477604 512038 477632 521591
rect 494164 512038 494192 521591
rect 477592 512032 477644 512038
rect 477592 511974 477644 511980
rect 477868 512032 477920 512038
rect 477868 511974 477920 511980
rect 494152 512032 494204 512038
rect 494152 511974 494204 511980
rect 494428 512032 494480 512038
rect 494428 511974 494480 511980
rect 477880 502382 477908 511974
rect 494440 502382 494468 511974
rect 477684 502376 477736 502382
rect 477406 502344 477462 502353
rect 477406 502279 477462 502288
rect 477682 502344 477684 502353
rect 477868 502376 477920 502382
rect 477736 502344 477738 502353
rect 494244 502376 494296 502382
rect 477868 502318 477920 502324
rect 493966 502344 494022 502353
rect 477682 502279 477738 502288
rect 493966 502279 494022 502288
rect 494242 502344 494244 502353
rect 494428 502376 494480 502382
rect 494296 502344 494298 502353
rect 494428 502318 494480 502324
rect 494242 502279 494298 502288
rect 477420 492697 477448 502279
rect 493980 492697 494008 502279
rect 477406 492688 477462 492697
rect 477406 492623 477462 492632
rect 477590 492688 477646 492697
rect 477590 492623 477646 492632
rect 493966 492688 494022 492697
rect 493966 492623 494022 492632
rect 494150 492688 494206 492697
rect 494150 492623 494206 492632
rect 477604 489954 477632 492623
rect 494164 489954 494192 492623
rect 477604 489926 477724 489954
rect 494164 489926 494284 489954
rect 477696 480282 477724 489926
rect 494256 480282 494284 489926
rect 477500 480276 477552 480282
rect 477500 480218 477552 480224
rect 477684 480276 477736 480282
rect 477684 480218 477736 480224
rect 494060 480276 494112 480282
rect 494060 480218 494112 480224
rect 494244 480276 494296 480282
rect 494244 480218 494296 480224
rect 477512 480162 477540 480218
rect 494072 480162 494100 480218
rect 477512 480134 477632 480162
rect 494072 480134 494192 480162
rect 477604 470642 477632 480134
rect 494164 470642 494192 480134
rect 477604 470614 477724 470642
rect 494164 470614 494284 470642
rect 477696 460970 477724 470614
rect 494256 460970 494284 470614
rect 477500 460964 477552 460970
rect 477500 460906 477552 460912
rect 477684 460964 477736 460970
rect 477684 460906 477736 460912
rect 494060 460964 494112 460970
rect 494060 460906 494112 460912
rect 494244 460964 494296 460970
rect 494244 460906 494296 460912
rect 477512 460850 477540 460906
rect 494072 460850 494100 460906
rect 477512 460822 477632 460850
rect 494072 460822 494192 460850
rect 477604 451330 477632 460822
rect 494164 451330 494192 460822
rect 477604 451302 477724 451330
rect 494164 451302 494284 451330
rect 477696 441658 477724 451302
rect 494256 441658 494284 451302
rect 477500 441652 477552 441658
rect 477500 441594 477552 441600
rect 477684 441652 477736 441658
rect 477684 441594 477736 441600
rect 494060 441652 494112 441658
rect 494060 441594 494112 441600
rect 494244 441652 494296 441658
rect 494244 441594 494296 441600
rect 477512 441538 477540 441594
rect 494072 441538 494100 441594
rect 477512 441510 477632 441538
rect 494072 441510 494192 441538
rect 477604 432018 477632 441510
rect 494164 432018 494192 441510
rect 477604 431990 477724 432018
rect 494164 431990 494284 432018
rect 462320 424720 462372 424726
rect 462320 424662 462372 424668
rect 477696 424658 477724 431990
rect 477684 424652 477736 424658
rect 477684 424594 477736 424600
rect 494256 424590 494284 431990
rect 494244 424584 494296 424590
rect 494244 424526 494296 424532
rect 527192 424522 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 694142 542768 698226
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 692782 542584 694078
rect 542544 692776 542596 692782
rect 542544 692718 542596 692724
rect 542728 692776 542780 692782
rect 542728 692718 542780 692724
rect 542740 683233 542768 692718
rect 559668 684486 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 567844 696992 567896 696998
rect 567844 696934 567896 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 558920 684480 558972 684486
rect 558920 684422 558972 684428
rect 559656 684480 559708 684486
rect 559656 684422 559708 684428
rect 542358 683224 542414 683233
rect 542358 683159 542414 683168
rect 542726 683224 542782 683233
rect 542726 683159 542782 683168
rect 542372 683126 542400 683159
rect 558932 683126 558960 684422
rect 542360 683120 542412 683126
rect 542360 683062 542412 683068
rect 558920 683120 558972 683126
rect 558920 683062 558972 683068
rect 558184 673532 558236 673538
rect 558184 673474 558236 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 542832 659682 542860 666538
rect 542648 659654 542860 659682
rect 542648 647290 542676 659654
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 542556 640422 542584 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 542648 630698 542676 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 542464 630578 542492 630634
rect 542464 630550 542584 630578
rect 542556 621058 542584 630550
rect 556804 626612 556856 626618
rect 556804 626554 556856 626560
rect 542556 621030 542676 621058
rect 542648 611386 542676 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 542464 611266 542492 611322
rect 542464 611238 542584 611266
rect 542556 608598 542584 611238
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 542740 598942 542768 601666
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 542832 582486 542860 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 542740 572642 542768 582286
rect 555424 579692 555476 579698
rect 555424 579634 555476 579640
rect 542556 572614 542768 572642
rect 542556 569922 542584 572614
rect 542464 569894 542584 569922
rect 542464 563174 542492 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 542464 560250 542492 562974
rect 542452 560244 542504 560250
rect 542452 560186 542504 560192
rect 542636 550656 542688 550662
rect 542636 550598 542688 550604
rect 542648 543658 542676 550598
rect 552664 545148 552716 545154
rect 552664 545090 552716 545096
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542636 543652 542688 543658
rect 542636 543594 542688 543600
rect 542464 534070 542492 543594
rect 542452 534064 542504 534070
rect 542452 534006 542504 534012
rect 542636 534064 542688 534070
rect 542636 534006 542688 534012
rect 542648 524482 542676 534006
rect 542636 524476 542688 524482
rect 542636 524418 542688 524424
rect 542728 524408 542780 524414
rect 542728 524350 542780 524356
rect 542740 521665 542768 524350
rect 542542 521656 542598 521665
rect 542542 521591 542598 521600
rect 542726 521656 542782 521665
rect 542726 521591 542782 521600
rect 542556 512038 542584 521591
rect 542544 512032 542596 512038
rect 542544 511974 542596 511980
rect 542820 512032 542872 512038
rect 542820 511974 542872 511980
rect 542832 502382 542860 511974
rect 551284 509312 551336 509318
rect 551284 509254 551336 509260
rect 542636 502376 542688 502382
rect 542358 502344 542414 502353
rect 542358 502279 542414 502288
rect 542634 502344 542636 502353
rect 542820 502376 542872 502382
rect 542688 502344 542690 502353
rect 542820 502318 542872 502324
rect 542634 502279 542690 502288
rect 542372 492697 542400 502279
rect 542358 492688 542414 492697
rect 542358 492623 542414 492632
rect 542542 492688 542598 492697
rect 542542 492623 542544 492632
rect 542596 492623 542598 492632
rect 542544 492594 542596 492600
rect 542544 485784 542596 485790
rect 542544 485726 542596 485732
rect 542556 483018 542584 485726
rect 542556 482990 542676 483018
rect 542648 476134 542676 482990
rect 542452 476128 542504 476134
rect 542636 476128 542688 476134
rect 542504 476076 542584 476082
rect 542452 476070 542584 476076
rect 542636 476070 542688 476076
rect 542464 476054 542584 476070
rect 542556 473346 542584 476054
rect 542544 473340 542596 473346
rect 542544 473282 542596 473288
rect 542544 466404 542596 466410
rect 542544 466346 542596 466352
rect 542556 463706 542584 466346
rect 542556 463678 542676 463706
rect 542648 454073 542676 463678
rect 542358 454064 542414 454073
rect 542358 453999 542414 454008
rect 542634 454064 542690 454073
rect 542634 453999 542690 454008
rect 542372 447166 542400 453999
rect 542360 447160 542412 447166
rect 542360 447102 542412 447108
rect 542452 447092 542504 447098
rect 542452 447034 542504 447040
rect 542464 437458 542492 447034
rect 542464 437430 542584 437458
rect 542556 434722 542584 437430
rect 542544 434716 542596 434722
rect 542544 434658 542596 434664
rect 542544 427780 542596 427786
rect 542544 427722 542596 427728
rect 542556 425082 542584 427722
rect 542556 425054 542676 425082
rect 370780 424516 370832 424522
rect 370780 424458 370832 424464
rect 527180 424516 527232 424522
rect 527180 424458 527232 424464
rect 364524 424380 364576 424386
rect 364524 424322 364576 424328
rect 370792 422348 370820 424458
rect 542648 424454 542676 425054
rect 382556 424448 382608 424454
rect 382556 424390 382608 424396
rect 542636 424448 542688 424454
rect 542636 424390 542688 424396
rect 382568 422348 382596 424390
rect 394332 424380 394384 424386
rect 394332 424322 394384 424328
rect 394344 422348 394372 424322
rect 78680 419484 78732 419490
rect 78680 419426 78732 419432
rect 401600 419484 401652 419490
rect 401600 419426 401652 419432
rect 78692 418577 78720 419426
rect 401612 418849 401640 419426
rect 401598 418840 401654 418849
rect 401598 418775 401654 418784
rect 78678 418568 78734 418577
rect 78678 418503 78734 418512
rect 425704 415472 425756 415478
rect 425704 415414 425756 415420
rect 401600 412616 401652 412622
rect 401600 412558 401652 412564
rect 401612 411777 401640 412558
rect 401598 411768 401654 411777
rect 401598 411703 401654 411712
rect 78680 411256 78732 411262
rect 78680 411198 78732 411204
rect 78692 410961 78720 411198
rect 78678 410952 78734 410961
rect 78678 410887 78734 410896
rect 401600 405680 401652 405686
rect 401600 405622 401652 405628
rect 401612 404569 401640 405622
rect 401598 404560 401654 404569
rect 401598 404495 401654 404504
rect 78680 404320 78732 404326
rect 78680 404262 78732 404268
rect 78692 403345 78720 404262
rect 78678 403336 78734 403345
rect 78678 403271 78734 403280
rect 401600 398812 401652 398818
rect 401600 398754 401652 398760
rect 401612 397497 401640 398754
rect 401598 397488 401654 397497
rect 401598 397423 401654 397432
rect 78680 396024 78732 396030
rect 78680 395966 78732 395972
rect 78692 395729 78720 395966
rect 78678 395720 78734 395729
rect 78678 395655 78734 395664
rect 407764 392012 407816 392018
rect 407764 391954 407816 391960
rect 401600 390516 401652 390522
rect 401600 390458 401652 390464
rect 401612 390425 401640 390458
rect 401598 390416 401654 390425
rect 401598 390351 401654 390360
rect 78680 389156 78732 389162
rect 78680 389098 78732 389104
rect 78692 388113 78720 389098
rect 78678 388104 78734 388113
rect 78678 388039 78734 388048
rect 401600 383648 401652 383654
rect 401600 383590 401652 383596
rect 401612 383217 401640 383590
rect 401598 383208 401654 383217
rect 401598 383143 401654 383152
rect 44824 380860 44876 380866
rect 44824 380802 44876 380808
rect 78680 380860 78732 380866
rect 78680 380802 78732 380808
rect 78692 380497 78720 380802
rect 78678 380488 78734 380497
rect 78678 380423 78734 380432
rect 401600 376712 401652 376718
rect 401600 376654 401652 376660
rect 401612 376145 401640 376654
rect 401598 376136 401654 376145
rect 401598 376071 401654 376080
rect 78680 373992 78732 373998
rect 78680 373934 78732 373940
rect 78692 372881 78720 373934
rect 78678 372872 78734 372881
rect 78678 372807 78734 372816
rect 401600 369844 401652 369850
rect 401600 369786 401652 369792
rect 401612 369073 401640 369786
rect 401598 369064 401654 369073
rect 401598 368999 401654 369008
rect 78680 365696 78732 365702
rect 78680 365638 78732 365644
rect 78692 365265 78720 365638
rect 78678 365256 78734 365265
rect 78678 365191 78734 365200
rect 401600 362908 401652 362914
rect 401600 362850 401652 362856
rect 401612 361865 401640 362850
rect 401598 361856 401654 361865
rect 401598 361791 401654 361800
rect 78680 358760 78732 358766
rect 78680 358702 78732 358708
rect 78692 357649 78720 358702
rect 78678 357640 78734 357649
rect 78678 357575 78734 357584
rect 405004 357468 405056 357474
rect 405004 357410 405056 357416
rect 401600 356040 401652 356046
rect 401600 355982 401652 355988
rect 401612 354793 401640 355982
rect 401598 354784 401654 354793
rect 401598 354719 401654 354728
rect 39304 350532 39356 350538
rect 39304 350474 39356 350480
rect 78680 350532 78732 350538
rect 78680 350474 78732 350480
rect 78692 350033 78720 350474
rect 78678 350024 78734 350033
rect 78678 349959 78734 349968
rect 401600 347744 401652 347750
rect 401598 347712 401600 347721
rect 401652 347712 401654 347721
rect 401598 347647 401654 347656
rect 403624 345092 403676 345098
rect 403624 345034 403676 345040
rect 78680 343596 78732 343602
rect 78680 343538 78732 343544
rect 78692 342281 78720 343538
rect 78678 342272 78734 342281
rect 78678 342207 78734 342216
rect 401600 340876 401652 340882
rect 401600 340818 401652 340824
rect 401612 340513 401640 340818
rect 401598 340504 401654 340513
rect 401598 340439 401654 340448
rect 37924 336796 37976 336802
rect 37924 336738 37976 336744
rect 21364 304972 21416 304978
rect 21364 304914 21416 304920
rect 37936 281518 37964 336738
rect 78680 335300 78732 335306
rect 78680 335242 78732 335248
rect 78692 334665 78720 335242
rect 78678 334656 78734 334665
rect 78678 334591 78734 334600
rect 401600 333940 401652 333946
rect 401600 333882 401652 333888
rect 401612 333441 401640 333882
rect 401598 333432 401654 333441
rect 401598 333367 401654 333376
rect 78680 327072 78732 327078
rect 78678 327040 78680 327049
rect 401600 327072 401652 327078
rect 78732 327040 78734 327049
rect 401600 327014 401652 327020
rect 78678 326975 78734 326984
rect 401612 326369 401640 327014
rect 401598 326360 401654 326369
rect 401598 326295 401654 326304
rect 78680 320136 78732 320142
rect 78680 320078 78732 320084
rect 401600 320136 401652 320142
rect 401600 320078 401652 320084
rect 78692 319433 78720 320078
rect 78678 319424 78734 319433
rect 78678 319359 78734 319368
rect 401612 319161 401640 320078
rect 401598 319152 401654 319161
rect 401598 319087 401654 319096
rect 401600 313268 401652 313274
rect 401600 313210 401652 313216
rect 401612 312089 401640 313210
rect 401598 312080 401654 312089
rect 401598 312015 401654 312024
rect 78680 311840 78732 311846
rect 78678 311808 78680 311817
rect 78732 311808 78734 311817
rect 78678 311743 78734 311752
rect 402244 305652 402296 305658
rect 402244 305594 402296 305600
rect 78680 304972 78732 304978
rect 78680 304914 78732 304920
rect 401600 304972 401652 304978
rect 401600 304914 401652 304920
rect 78692 304201 78720 304914
rect 401612 304881 401640 304914
rect 401598 304872 401654 304881
rect 401598 304807 401654 304816
rect 78678 304192 78734 304201
rect 78678 304127 78734 304136
rect 401600 298104 401652 298110
rect 401600 298046 401652 298052
rect 401612 297809 401640 298046
rect 401598 297800 401654 297809
rect 401598 297735 401654 297744
rect 78680 296676 78732 296682
rect 78680 296618 78732 296624
rect 78692 296585 78720 296618
rect 78678 296576 78734 296585
rect 78678 296511 78734 296520
rect 401600 291168 401652 291174
rect 401600 291110 401652 291116
rect 401612 290737 401640 291110
rect 401598 290728 401654 290737
rect 401598 290663 401654 290672
rect 78680 289808 78732 289814
rect 78680 289750 78732 289756
rect 78692 288969 78720 289750
rect 78678 288960 78734 288969
rect 78678 288895 78734 288904
rect 401600 284300 401652 284306
rect 401600 284242 401652 284248
rect 401612 283529 401640 284242
rect 401598 283520 401654 283529
rect 401598 283455 401654 283464
rect 37924 281512 37976 281518
rect 37924 281454 37976 281460
rect 78680 281512 78732 281518
rect 78680 281454 78732 281460
rect 78692 281353 78720 281454
rect 78678 281344 78734 281353
rect 78678 281279 78734 281288
rect 401600 277364 401652 277370
rect 401600 277306 401652 277312
rect 401612 276457 401640 277306
rect 401598 276448 401654 276457
rect 401598 276383 401654 276392
rect 78680 274644 78732 274650
rect 78680 274586 78732 274592
rect 78692 273737 78720 274586
rect 78678 273728 78734 273737
rect 78678 273663 78734 273672
rect 401600 270496 401652 270502
rect 401600 270438 401652 270444
rect 401612 269385 401640 270438
rect 401598 269376 401654 269385
rect 401598 269311 401654 269320
rect 3700 266348 3752 266354
rect 3700 266290 3752 266296
rect 78680 266348 78732 266354
rect 78680 266290 78732 266296
rect 78692 266121 78720 266290
rect 78678 266112 78734 266121
rect 78678 266047 78734 266056
rect 3606 265704 3662 265713
rect 3606 265639 3662 265648
rect 3516 251184 3568 251190
rect 3516 251126 3568 251132
rect 3620 244254 3648 265639
rect 401600 262200 401652 262206
rect 401598 262168 401600 262177
rect 401652 262168 401654 262177
rect 401598 262103 401654 262112
rect 78680 259412 78732 259418
rect 78680 259354 78732 259360
rect 78692 258369 78720 259354
rect 78678 258360 78734 258369
rect 78678 258295 78734 258304
rect 401600 255128 401652 255134
rect 401598 255096 401600 255105
rect 401652 255096 401654 255105
rect 401598 255031 401654 255040
rect 78680 251184 78732 251190
rect 78680 251126 78732 251132
rect 78692 250753 78720 251126
rect 78678 250744 78734 250753
rect 78678 250679 78734 250688
rect 402256 248033 402284 305594
rect 403636 255134 403664 345034
rect 405016 262206 405044 357410
rect 407776 277370 407804 391954
rect 409144 310548 409196 310554
rect 409144 310490 409196 310496
rect 407764 277364 407816 277370
rect 407764 277306 407816 277312
rect 407764 263628 407816 263634
rect 407764 263570 407816 263576
rect 405004 262200 405056 262206
rect 405004 262142 405056 262148
rect 403624 255128 403676 255134
rect 403624 255070 403676 255076
rect 403624 251252 403676 251258
rect 403624 251194 403676 251200
rect 402242 248024 402298 248033
rect 402242 247959 402298 247968
rect 3608 244248 3660 244254
rect 3608 244190 3660 244196
rect 78680 244248 78732 244254
rect 78680 244190 78732 244196
rect 78692 243137 78720 244190
rect 78678 243128 78734 243137
rect 78678 243063 78734 243072
rect 401600 241460 401652 241466
rect 401600 241402 401652 241408
rect 401612 240825 401640 241402
rect 401598 240816 401654 240825
rect 401598 240751 401654 240760
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3424 235952 3476 235958
rect 3424 235894 3476 235900
rect 3528 229090 3556 236943
rect 78680 235952 78732 235958
rect 78680 235894 78732 235900
rect 78692 235521 78720 235894
rect 78678 235512 78734 235521
rect 78678 235447 78734 235456
rect 401600 234592 401652 234598
rect 401600 234534 401652 234540
rect 401612 233753 401640 234534
rect 401598 233744 401654 233753
rect 401598 233679 401654 233688
rect 3516 229084 3568 229090
rect 3516 229026 3568 229032
rect 78680 229084 78732 229090
rect 78680 229026 78732 229032
rect 78692 227905 78720 229026
rect 78678 227896 78734 227905
rect 78678 227831 78734 227840
rect 401600 227724 401652 227730
rect 401600 227666 401652 227672
rect 401612 226681 401640 227666
rect 401598 226672 401654 226681
rect 401598 226607 401654 226616
rect 2962 222592 3018 222601
rect 2962 222527 3018 222536
rect 2976 220794 3004 222527
rect 2964 220788 3016 220794
rect 2964 220730 3016 220736
rect 78680 220788 78732 220794
rect 78680 220730 78732 220736
rect 401600 220788 401652 220794
rect 401600 220730 401652 220736
rect 78692 220289 78720 220730
rect 78678 220280 78734 220289
rect 78678 220215 78734 220224
rect 401612 219473 401640 220730
rect 401598 219464 401654 219473
rect 401598 219399 401654 219408
rect 79322 212664 79378 212673
rect 79322 212599 79378 212608
rect 79336 208350 79364 212599
rect 403636 212430 403664 251194
rect 405004 227792 405056 227798
rect 405004 227734 405056 227740
rect 401600 212424 401652 212430
rect 401598 212392 401600 212401
rect 403624 212424 403676 212430
rect 401652 212392 401654 212401
rect 403624 212366 403676 212372
rect 401598 212327 401654 212336
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 79324 208344 79376 208350
rect 79324 208286 79376 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 405016 205630 405044 227734
rect 407776 220794 407804 263570
rect 409156 241466 409184 310490
rect 425716 291174 425744 415414
rect 551296 333946 551324 509254
rect 552676 347750 552704 545090
rect 554044 485852 554096 485858
rect 554044 485794 554096 485800
rect 552664 347744 552716 347750
rect 552664 347686 552716 347692
rect 551284 333940 551336 333946
rect 551284 333882 551336 333888
rect 554056 320142 554084 485794
rect 555436 362914 555464 579634
rect 556816 383654 556844 626554
rect 558196 405686 558224 673474
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 559392 659682 559420 666538
rect 559208 659654 559420 659682
rect 559208 647290 559236 659654
rect 566464 650072 566516 650078
rect 566464 650014 566516 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 559208 630698 559236 640358
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 559116 621058 559144 630550
rect 559116 621030 559236 621058
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 565084 603152 565136 603158
rect 565084 603094 565136 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 559392 582486 559420 589290
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 559300 572642 559328 582286
rect 559116 572614 559328 572642
rect 559116 569922 559144 572614
rect 559024 569894 559144 569922
rect 559024 563174 559052 569894
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 559024 560250 559052 562974
rect 559012 560244 559064 560250
rect 559012 560186 559064 560192
rect 563704 556232 563756 556238
rect 563704 556174 563756 556180
rect 559196 550656 559248 550662
rect 559196 550598 559248 550604
rect 559208 543658 559236 550598
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559196 543652 559248 543658
rect 559196 543594 559248 543600
rect 559024 534070 559052 543594
rect 559012 534064 559064 534070
rect 559012 534006 559064 534012
rect 559196 534064 559248 534070
rect 559196 534006 559248 534012
rect 559208 524482 559236 534006
rect 559196 524476 559248 524482
rect 559196 524418 559248 524424
rect 559288 524408 559340 524414
rect 559288 524350 559340 524356
rect 559300 521665 559328 524350
rect 559102 521656 559158 521665
rect 559102 521591 559158 521600
rect 559286 521656 559342 521665
rect 559286 521591 559342 521600
rect 559116 512038 559144 521591
rect 559104 512032 559156 512038
rect 559104 511974 559156 511980
rect 559380 512032 559432 512038
rect 559380 511974 559432 511980
rect 559392 502382 559420 511974
rect 559196 502376 559248 502382
rect 558918 502344 558974 502353
rect 558918 502279 558974 502288
rect 559194 502344 559196 502353
rect 559380 502376 559432 502382
rect 559248 502344 559250 502353
rect 559380 502318 559432 502324
rect 559194 502279 559250 502288
rect 558932 492697 558960 502279
rect 558918 492688 558974 492697
rect 558918 492623 558974 492632
rect 559102 492688 559158 492697
rect 559102 492623 559104 492632
rect 559156 492623 559158 492632
rect 559104 492594 559156 492600
rect 559104 485784 559156 485790
rect 559104 485726 559156 485732
rect 559116 483018 559144 485726
rect 559116 482990 559236 483018
rect 559208 476134 559236 482990
rect 559012 476128 559064 476134
rect 559196 476128 559248 476134
rect 559064 476076 559144 476082
rect 559012 476070 559144 476076
rect 559196 476070 559248 476076
rect 559024 476054 559144 476070
rect 559116 473346 559144 476054
rect 559104 473340 559156 473346
rect 559104 473282 559156 473288
rect 559104 466404 559156 466410
rect 559104 466346 559156 466352
rect 559116 463706 559144 466346
rect 559116 463678 559236 463706
rect 559208 454073 559236 463678
rect 558918 454064 558974 454073
rect 558918 453999 558974 454008
rect 559194 454064 559250 454073
rect 559194 453999 559250 454008
rect 558932 447166 558960 453999
rect 558920 447160 558972 447166
rect 558920 447102 558972 447108
rect 559012 447092 559064 447098
rect 559012 447034 559064 447040
rect 559024 437458 559052 447034
rect 560944 438932 560996 438938
rect 560944 438874 560996 438880
rect 559024 437430 559144 437458
rect 559116 434722 559144 437430
rect 559104 434716 559156 434722
rect 559104 434658 559156 434664
rect 559104 427780 559156 427786
rect 559104 427722 559156 427728
rect 559116 425082 559144 427722
rect 559116 425054 559236 425082
rect 559208 424386 559236 425054
rect 559196 424380 559248 424386
rect 559196 424322 559248 424328
rect 558184 405680 558236 405686
rect 558184 405622 558236 405628
rect 556804 383648 556856 383654
rect 556804 383590 556856 383596
rect 555424 362908 555476 362914
rect 555424 362850 555476 362856
rect 554044 320136 554096 320142
rect 554044 320078 554096 320084
rect 560956 298110 560984 438874
rect 563716 356046 563744 556174
rect 565096 376718 565124 603094
rect 566476 398818 566504 650014
rect 567856 419490 567884 696934
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 573364 638988 573416 638994
rect 573364 638930 573416 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 570604 592068 570656 592074
rect 570604 592010 570656 592016
rect 569224 498228 569276 498234
rect 569224 498170 569276 498176
rect 567844 419484 567896 419490
rect 567844 419426 567896 419432
rect 566464 398812 566516 398818
rect 566464 398754 566516 398760
rect 565084 376712 565136 376718
rect 565084 376654 565136 376660
rect 563704 356040 563756 356046
rect 563704 355982 563756 355988
rect 569236 327078 569264 498170
rect 570616 369850 570644 592010
rect 571984 462392 572036 462398
rect 571984 462334 572036 462340
rect 570604 369844 570656 369850
rect 570604 369786 570656 369792
rect 569224 327072 569276 327078
rect 569224 327014 569276 327020
rect 571996 313274 572024 462334
rect 573376 390522 573404 638930
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 578882 533896 578938 533905
rect 578882 533831 578938 533840
rect 573364 390516 573416 390522
rect 573364 390458 573416 390464
rect 576124 368552 576176 368558
rect 576124 368494 576176 368500
rect 571984 313268 572036 313274
rect 571984 313210 572036 313216
rect 560944 298104 560996 298110
rect 560944 298046 560996 298052
rect 425704 291168 425756 291174
rect 425704 291110 425756 291116
rect 425704 274712 425756 274718
rect 425704 274654 425756 274660
rect 409144 241460 409196 241466
rect 409144 241402 409196 241408
rect 425716 227730 425744 274654
rect 576136 270502 576164 368494
rect 578896 340882 578924 533831
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 579894 486840 579950 486849
rect 579894 486775 579950 486784
rect 579908 485858 579936 486775
rect 579896 485852 579948 485858
rect 579896 485794 579948 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 580276 412622 580304 686287
rect 580354 451752 580410 451761
rect 580354 451687 580410 451696
rect 580264 412616 580316 412622
rect 580264 412558 580316 412564
rect 580262 404832 580318 404841
rect 580262 404767 580318 404776
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 579894 357912 579950 357921
rect 579894 357847 579950 357856
rect 579908 357474 579936 357847
rect 579896 357468 579948 357474
rect 579896 357410 579948 357416
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 578884 340876 578936 340882
rect 578884 340818 578936 340824
rect 578882 322688 578938 322697
rect 578882 322623 578938 322632
rect 578896 305658 578924 322623
rect 579618 310856 579674 310865
rect 579618 310791 579674 310800
rect 579632 310554 579660 310791
rect 579620 310548 579672 310554
rect 579620 310490 579672 310496
rect 578884 305652 578936 305658
rect 578884 305594 578936 305600
rect 578882 299160 578938 299169
rect 578882 299095 578938 299104
rect 576124 270496 576176 270502
rect 576124 270438 576176 270444
rect 578896 234598 578924 299095
rect 580276 284306 580304 404767
rect 580368 304978 580396 451687
rect 580356 304972 580408 304978
rect 580356 304914 580408 304920
rect 580264 284300 580316 284306
rect 580264 284242 580316 284248
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580184 274718 580212 275703
rect 580172 274712 580224 274718
rect 580172 274654 580224 274660
rect 579802 263936 579858 263945
rect 579802 263871 579858 263880
rect 579816 263634 579844 263871
rect 579804 263628 579856 263634
rect 579804 263570 579856 263576
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 251258 580212 252175
rect 580172 251252 580224 251258
rect 580172 251194 580224 251200
rect 578884 234592 578936 234598
rect 578884 234534 578936 234540
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580184 227798 580212 228783
rect 580172 227792 580224 227798
rect 580172 227734 580224 227740
rect 425704 227724 425756 227730
rect 425704 227666 425756 227672
rect 407764 220788 407816 220794
rect 407764 220730 407816 220736
rect 580262 217016 580318 217025
rect 580262 216951 580318 216960
rect 401600 205624 401652 205630
rect 401600 205566 401652 205572
rect 405004 205624 405056 205630
rect 405004 205566 405056 205572
rect 401612 205193 401640 205566
rect 401598 205184 401654 205193
rect 401598 205119 401654 205128
rect 79322 205048 79378 205057
rect 79322 204983 79378 204992
rect 79336 194546 79364 204983
rect 580276 198694 580304 216951
rect 580354 205320 580410 205329
rect 580354 205255 580410 205264
rect 401600 198688 401652 198694
rect 401600 198630 401652 198636
rect 580264 198688 580316 198694
rect 580264 198630 580316 198636
rect 401612 198121 401640 198630
rect 401598 198112 401654 198121
rect 401598 198047 401654 198056
rect 79414 197432 79470 197441
rect 79414 197367 79470 197376
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 79324 194540 79376 194546
rect 79324 194482 79376 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 79322 189816 79378 189825
rect 79322 189751 79378 189760
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 78678 166832 78734 166841
rect 78678 166767 78734 166776
rect 78692 165646 78720 166767
rect 21364 165640 21416 165646
rect 21364 165582 21416 165588
rect 78680 165640 78732 165646
rect 78680 165582 78732 165588
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 8944 143608 8996 143614
rect 8944 143550 8996 143556
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 8956 79490 8984 143550
rect 21376 122806 21404 165582
rect 79336 165578 79364 189751
rect 79428 180810 79456 197367
rect 580368 191826 580396 205255
rect 401600 191820 401652 191826
rect 401600 191762 401652 191768
rect 580356 191820 580408 191826
rect 580356 191762 580408 191768
rect 401612 191049 401640 191762
rect 401598 191040 401654 191049
rect 401598 190975 401654 190984
rect 401598 183832 401654 183841
rect 401598 183767 401654 183776
rect 401612 182170 401640 183767
rect 401600 182164 401652 182170
rect 401600 182106 401652 182112
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 79506 182064 79562 182073
rect 79506 181999 79562 182008
rect 79416 180804 79468 180810
rect 79416 180746 79468 180752
rect 79414 174448 79470 174457
rect 79414 174383 79470 174392
rect 79324 165572 79376 165578
rect 79324 165514 79376 165520
rect 79322 159216 79378 159225
rect 79322 159151 79378 159160
rect 78678 143984 78734 143993
rect 78678 143919 78734 143928
rect 78692 143614 78720 143919
rect 78680 143608 78732 143614
rect 78680 143550 78732 143556
rect 21364 122800 21416 122806
rect 21364 122742 21416 122748
rect 78678 121136 78734 121145
rect 78678 121071 78734 121080
rect 78692 120154 78720 121071
rect 21364 120148 21416 120154
rect 21364 120090 21416 120096
rect 78680 120148 78732 120154
rect 78680 120090 78732 120096
rect 3516 79484 3568 79490
rect 3516 79426 3568 79432
rect 8944 79484 8996 79490
rect 8944 79426 8996 79432
rect 3528 78985 3556 79426
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 21376 35902 21404 120090
rect 79336 109002 79364 159151
rect 79428 136610 79456 174383
rect 79520 151774 79548 181999
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 402242 176760 402298 176769
rect 402242 176695 402298 176704
rect 402256 171086 402284 176695
rect 402244 171080 402296 171086
rect 402244 171022 402296 171028
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 402242 169688 402298 169697
rect 402242 169623 402298 169632
rect 402256 158710 402284 169623
rect 402334 162480 402390 162489
rect 402334 162415 402390 162424
rect 402244 158704 402296 158710
rect 402244 158646 402296 158652
rect 402242 155408 402298 155417
rect 402242 155343 402298 155352
rect 79508 151768 79560 151774
rect 79508 151710 79560 151716
rect 79690 151600 79746 151609
rect 79690 151535 79746 151544
rect 79416 136604 79468 136610
rect 79416 136546 79468 136552
rect 79598 136368 79654 136377
rect 79598 136303 79654 136312
rect 79506 128752 79562 128761
rect 79506 128687 79562 128696
rect 79414 113520 79470 113529
rect 79414 113455 79470 113464
rect 79324 108996 79376 109002
rect 79324 108938 79376 108944
rect 79322 105904 79378 105913
rect 79322 105839 79378 105848
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 21364 35896 21416 35902
rect 3476 35864 3478 35873
rect 21364 35838 21416 35844
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 79336 8294 79364 105839
rect 79428 22098 79456 113455
rect 79520 51066 79548 128687
rect 79612 64870 79640 136303
rect 79704 93838 79732 151535
rect 401598 126984 401654 126993
rect 401598 126919 401654 126928
rect 401612 125662 401640 126919
rect 401600 125656 401652 125662
rect 401600 125598 401652 125604
rect 402256 124166 402284 155343
rect 402348 135250 402376 162415
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 402610 148336 402666 148345
rect 402610 148271 402666 148280
rect 402518 141128 402574 141137
rect 402518 141063 402574 141072
rect 402336 135244 402388 135250
rect 402336 135186 402388 135192
rect 402426 134056 402482 134065
rect 402426 133991 402482 134000
rect 402244 124160 402296 124166
rect 402244 124102 402296 124108
rect 402334 119776 402390 119785
rect 402334 119711 402390 119720
rect 402242 112704 402298 112713
rect 402242 112639 402298 112648
rect 401598 105632 401654 105641
rect 401598 105567 401654 105576
rect 401612 104922 401640 105567
rect 401600 104916 401652 104922
rect 401600 104858 401652 104864
rect 370884 102190 370990 102218
rect 370884 102134 370912 102190
rect 370872 102128 370924 102134
rect 81452 102054 82386 102082
rect 82924 102054 83122 102082
rect 83950 102054 84148 102082
rect 84778 102054 85528 102082
rect 79692 93832 79744 93838
rect 79692 93774 79744 93780
rect 79600 64864 79652 64870
rect 79600 64806 79652 64812
rect 79508 51060 79560 51066
rect 79508 51002 79560 51008
rect 79416 22092 79468 22098
rect 79416 22034 79468 22040
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 79324 8288 79376 8294
rect 79324 8230 79376 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 81452 3534 81480 102054
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 81440 3528 81492 3534
rect 81440 3470 81492 3476
rect 584 480 612 3470
rect 82924 3466 82952 102054
rect 84120 4894 84148 102054
rect 85500 14482 85528 102054
rect 85592 100026 85620 102068
rect 86434 102054 86908 102082
rect 85580 100020 85632 100026
rect 85580 99962 85632 99968
rect 86880 15910 86908 102054
rect 87248 99482 87276 102068
rect 88090 102054 88288 102082
rect 87236 99476 87288 99482
rect 87236 99418 87288 99424
rect 86868 15904 86920 15910
rect 86868 15846 86920 15852
rect 85488 14476 85540 14482
rect 85488 14418 85540 14424
rect 84108 4888 84160 4894
rect 84108 4830 84160 4836
rect 88260 4010 88288 102054
rect 88904 99414 88932 102068
rect 89732 100706 89760 102068
rect 90574 102054 91048 102082
rect 89720 100700 89772 100706
rect 89720 100642 89772 100648
rect 90916 100700 90968 100706
rect 90916 100642 90968 100648
rect 88984 99476 89036 99482
rect 88984 99418 89036 99424
rect 88892 99408 88944 99414
rect 88892 99350 88944 99356
rect 88996 21418 89024 99418
rect 89628 99408 89680 99414
rect 89628 99350 89680 99356
rect 88984 21412 89036 21418
rect 88984 21354 89036 21360
rect 89640 17270 89668 99350
rect 90928 28286 90956 100642
rect 90916 28280 90968 28286
rect 90916 28222 90968 28228
rect 89628 17264 89680 17270
rect 89628 17206 89680 17212
rect 88248 4004 88300 4010
rect 88248 3946 88300 3952
rect 91020 3942 91048 102054
rect 91388 98666 91416 102068
rect 92124 102054 92230 102082
rect 93058 102054 93808 102082
rect 91376 98660 91428 98666
rect 91376 98602 91428 98608
rect 92124 95334 92152 102054
rect 92388 98660 92440 98666
rect 92388 98602 92440 98608
rect 92112 95328 92164 95334
rect 92112 95270 92164 95276
rect 92296 95260 92348 95266
rect 92296 95202 92348 95208
rect 92308 95146 92336 95202
rect 92216 95118 92336 95146
rect 92216 89758 92244 95118
rect 92204 89752 92256 89758
rect 92204 89694 92256 89700
rect 92204 85604 92256 85610
rect 92204 85546 92256 85552
rect 92216 85513 92244 85546
rect 91926 85504 91982 85513
rect 91926 85439 91982 85448
rect 92202 85504 92258 85513
rect 92202 85439 92258 85448
rect 91940 80782 91968 85439
rect 91928 80776 91980 80782
rect 91928 80718 91980 80724
rect 92296 67652 92348 67658
rect 92296 67594 92348 67600
rect 92308 60602 92336 67594
rect 92216 60574 92336 60602
rect 92216 57934 92244 60574
rect 92204 57928 92256 57934
rect 92204 57870 92256 57876
rect 92112 48340 92164 48346
rect 92112 48282 92164 48288
rect 92124 47598 92152 48282
rect 92112 47592 92164 47598
rect 92112 47534 92164 47540
rect 92400 18630 92428 98602
rect 92388 18624 92440 18630
rect 92388 18566 92440 18572
rect 91008 3936 91060 3942
rect 91008 3878 91060 3884
rect 93780 3874 93808 102054
rect 93872 100638 93900 102068
rect 94714 102054 95188 102082
rect 93860 100632 93912 100638
rect 93860 100574 93912 100580
rect 95160 49026 95188 102054
rect 95528 99754 95556 102068
rect 96264 102054 96370 102082
rect 95516 99748 95568 99754
rect 95516 99690 95568 99696
rect 96264 96665 96292 102054
rect 97184 100706 97212 102068
rect 98012 100706 98040 102068
rect 98854 102054 99236 102082
rect 97172 100700 97224 100706
rect 97172 100642 97224 100648
rect 97908 100700 97960 100706
rect 97908 100642 97960 100648
rect 98000 100700 98052 100706
rect 98000 100642 98052 100648
rect 97264 100632 97316 100638
rect 97264 100574 97316 100580
rect 96528 99748 96580 99754
rect 96528 99690 96580 99696
rect 96250 96656 96306 96665
rect 96250 96591 96306 96600
rect 96434 96656 96490 96665
rect 96434 96591 96490 96600
rect 96448 85610 96476 96591
rect 96344 85604 96396 85610
rect 96344 85546 96396 85552
rect 96436 85604 96488 85610
rect 96436 85546 96488 85552
rect 96356 80753 96384 85546
rect 96342 80744 96398 80753
rect 96342 80679 96398 80688
rect 96342 67688 96398 67697
rect 96342 67623 96398 67632
rect 96356 66230 96384 67623
rect 96344 66224 96396 66230
rect 96344 66166 96396 66172
rect 96252 56636 96304 56642
rect 96252 56578 96304 56584
rect 96264 56506 96292 56578
rect 96252 56500 96304 56506
rect 96252 56442 96304 56448
rect 95148 49020 95200 49026
rect 95148 48962 95200 48968
rect 96344 46980 96396 46986
rect 96344 46922 96396 46928
rect 96356 41478 96384 46922
rect 96344 41472 96396 41478
rect 96344 41414 96396 41420
rect 96252 41404 96304 41410
rect 96252 41346 96304 41352
rect 96264 31822 96292 41346
rect 96252 31816 96304 31822
rect 96252 31758 96304 31764
rect 96160 31748 96212 31754
rect 96160 31690 96212 31696
rect 96172 22778 96200 31690
rect 96160 22772 96212 22778
rect 96160 22714 96212 22720
rect 93768 3868 93820 3874
rect 93768 3810 93820 3816
rect 96540 3806 96568 99690
rect 97276 19990 97304 100574
rect 97920 51746 97948 100642
rect 97908 51740 97960 51746
rect 97908 51682 97960 51688
rect 99208 24138 99236 102054
rect 99668 100706 99696 102068
rect 100510 102054 100708 102082
rect 101338 102054 102088 102082
rect 99288 100700 99340 100706
rect 99288 100642 99340 100648
rect 99656 100700 99708 100706
rect 99656 100642 99708 100648
rect 100576 100700 100628 100706
rect 100576 100642 100628 100648
rect 99196 24132 99248 24138
rect 99196 24074 99248 24080
rect 97264 19984 97316 19990
rect 97264 19926 97316 19932
rect 96528 3800 96580 3806
rect 96528 3742 96580 3748
rect 99300 3738 99328 100642
rect 100588 53106 100616 100642
rect 100576 53100 100628 53106
rect 100576 53042 100628 53048
rect 99288 3732 99340 3738
rect 99288 3674 99340 3680
rect 100680 3602 100708 102054
rect 102060 25566 102088 102054
rect 102152 100706 102180 102068
rect 102994 102054 103468 102082
rect 102140 100700 102192 100706
rect 102140 100642 102192 100648
rect 103336 100700 103388 100706
rect 103336 100642 103388 100648
rect 103348 55894 103376 100642
rect 103336 55888 103388 55894
rect 103336 55830 103388 55836
rect 102048 25560 102100 25566
rect 102048 25502 102100 25508
rect 103440 3670 103468 102054
rect 103808 99618 103836 102068
rect 104544 102054 104650 102082
rect 103796 99612 103848 99618
rect 103796 99554 103848 99560
rect 104544 96665 104572 102054
rect 105372 100706 105400 102068
rect 106108 102054 106214 102082
rect 107042 102054 107608 102082
rect 105360 100700 105412 100706
rect 105360 100642 105412 100648
rect 104808 99612 104860 99618
rect 104808 99554 104860 99560
rect 104530 96656 104586 96665
rect 104530 96591 104586 96600
rect 104714 96656 104770 96665
rect 104714 96591 104770 96600
rect 104728 87038 104756 96591
rect 104624 87032 104676 87038
rect 104624 86974 104676 86980
rect 104716 87032 104768 87038
rect 104716 86974 104768 86980
rect 104636 82142 104664 86974
rect 104624 82136 104676 82142
rect 104624 82078 104676 82084
rect 104624 77376 104676 77382
rect 104544 77324 104624 77330
rect 104544 77318 104676 77324
rect 104544 77302 104664 77318
rect 104544 77246 104572 77302
rect 104532 77240 104584 77246
rect 104532 77182 104584 77188
rect 104624 67652 104676 67658
rect 104624 67594 104676 67600
rect 104636 60858 104664 67594
rect 104624 60852 104676 60858
rect 104624 60794 104676 60800
rect 104532 60716 104584 60722
rect 104532 60658 104584 60664
rect 104544 57254 104572 60658
rect 104532 57248 104584 57254
rect 104532 57190 104584 57196
rect 104820 26926 104848 99554
rect 106108 29646 106136 102054
rect 106188 100700 106240 100706
rect 106188 100642 106240 100648
rect 106096 29640 106148 29646
rect 106096 29582 106148 29588
rect 104808 26920 104860 26926
rect 104808 26862 104860 26868
rect 103428 3664 103480 3670
rect 103428 3606 103480 3612
rect 100668 3596 100720 3602
rect 100668 3538 100720 3544
rect 106200 3534 106228 100642
rect 106924 100020 106976 100026
rect 106924 99962 106976 99968
rect 106936 13190 106964 99962
rect 107580 58682 107608 102054
rect 107856 100706 107884 102068
rect 107844 100700 107896 100706
rect 107844 100642 107896 100648
rect 108684 100094 108712 102068
rect 108948 100700 109000 100706
rect 108948 100642 109000 100648
rect 108672 100088 108724 100094
rect 108672 100030 108724 100036
rect 107568 58676 107620 58682
rect 107568 58618 107620 58624
rect 106924 13184 106976 13190
rect 106924 13126 106976 13132
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 108960 3466 108988 100642
rect 109512 99414 109540 102068
rect 109500 99408 109552 99414
rect 109500 99350 109552 99356
rect 110340 61402 110368 102068
rect 111182 102054 111748 102082
rect 111064 99408 111116 99414
rect 111064 99350 111116 99356
rect 110328 61396 110380 61402
rect 110328 61338 110380 61344
rect 111076 31074 111104 99350
rect 111064 31068 111116 31074
rect 111064 31010 111116 31016
rect 111720 6186 111748 102054
rect 111996 99414 112024 102068
rect 112838 102054 113128 102082
rect 113666 102054 114416 102082
rect 111984 99408 112036 99414
rect 111984 99350 112036 99356
rect 113100 62830 113128 102054
rect 113088 62824 113140 62830
rect 113088 62766 113140 62772
rect 114388 44946 114416 102054
rect 114376 44940 114428 44946
rect 114376 44882 114428 44888
rect 114480 33794 114508 102068
rect 115322 102054 115888 102082
rect 115204 99408 115256 99414
rect 115204 99350 115256 99356
rect 114468 33788 114520 33794
rect 114468 33730 114520 33736
rect 115216 32434 115244 99350
rect 115860 64190 115888 102054
rect 116136 99414 116164 102068
rect 116978 102054 117176 102082
rect 116124 99408 116176 99414
rect 116124 99350 116176 99356
rect 115848 64184 115900 64190
rect 115848 64126 115900 64132
rect 117148 35222 117176 102054
rect 117792 99414 117820 102068
rect 117228 99408 117280 99414
rect 117228 99350 117280 99356
rect 117780 99408 117832 99414
rect 117780 99350 117832 99356
rect 118516 99408 118568 99414
rect 118516 99350 118568 99356
rect 117136 35216 117188 35222
rect 117136 35158 117188 35164
rect 115204 32428 115256 32434
rect 115204 32370 115256 32376
rect 117240 7614 117268 99350
rect 118528 66910 118556 99350
rect 118516 66904 118568 66910
rect 118516 66846 118568 66852
rect 118620 8974 118648 102068
rect 119462 102054 120028 102082
rect 120000 36582 120028 102054
rect 120276 99414 120304 102068
rect 121118 102054 121408 102082
rect 120264 99408 120316 99414
rect 120264 99350 120316 99356
rect 121276 99408 121328 99414
rect 121276 99350 121328 99356
rect 121288 68338 121316 99350
rect 121276 68332 121328 68338
rect 121276 68274 121328 68280
rect 119988 36576 120040 36582
rect 119988 36518 120040 36524
rect 121380 10334 121408 102054
rect 121932 99414 121960 102068
rect 122668 102054 122774 102082
rect 123602 102054 124168 102082
rect 121920 99408 121972 99414
rect 121920 99350 121972 99356
rect 122668 69698 122696 102054
rect 122748 99408 122800 99414
rect 122748 99350 122800 99356
rect 122656 69692 122708 69698
rect 122656 69634 122708 69640
rect 122760 37942 122788 99350
rect 122748 37936 122800 37942
rect 122748 37878 122800 37884
rect 124140 11762 124168 102054
rect 124416 99414 124444 102068
rect 125258 102054 125456 102082
rect 124404 99408 124456 99414
rect 124404 99350 124456 99356
rect 125428 71058 125456 102054
rect 126072 99414 126100 102068
rect 126808 102054 126914 102082
rect 127742 102054 128308 102082
rect 125508 99408 125560 99414
rect 125508 99350 125560 99356
rect 126060 99408 126112 99414
rect 126060 99350 126112 99356
rect 125416 71052 125468 71058
rect 125416 70994 125468 71000
rect 124128 11756 124180 11762
rect 124128 11698 124180 11704
rect 121368 10328 121420 10334
rect 121368 10270 121420 10276
rect 118608 8968 118660 8974
rect 118608 8910 118660 8916
rect 117228 7608 117280 7614
rect 117228 7550 117280 7556
rect 111708 6180 111760 6186
rect 111708 6122 111760 6128
rect 125520 4826 125548 99350
rect 126808 39370 126836 102054
rect 126888 99408 126940 99414
rect 126888 99350 126940 99356
rect 126796 39364 126848 39370
rect 126796 39306 126848 39312
rect 126900 13122 126928 99350
rect 128280 75206 128308 102054
rect 128464 99414 128492 102068
rect 129306 102054 129596 102082
rect 128452 99408 128504 99414
rect 128452 99350 128504 99356
rect 128268 75200 128320 75206
rect 128268 75142 128320 75148
rect 129568 40730 129596 102054
rect 130120 99414 130148 102068
rect 130948 99482 130976 102068
rect 131790 102054 132448 102082
rect 130936 99476 130988 99482
rect 130936 99418 130988 99424
rect 131764 99476 131816 99482
rect 131764 99418 131816 99424
rect 129648 99408 129700 99414
rect 129648 99350 129700 99356
rect 130108 99408 130160 99414
rect 130108 99350 130160 99356
rect 131028 99408 131080 99414
rect 131028 99350 131080 99356
rect 129556 40724 129608 40730
rect 129556 40666 129608 40672
rect 129660 14482 129688 99350
rect 131040 76566 131068 99350
rect 131028 76560 131080 76566
rect 131028 76502 131080 76508
rect 131120 21412 131172 21418
rect 131120 21354 131172 21360
rect 129740 15904 129792 15910
rect 129740 15846 129792 15852
rect 126980 14476 127032 14482
rect 126980 14418 127032 14424
rect 129648 14476 129700 14482
rect 129648 14418 129700 14424
rect 126888 13116 126940 13122
rect 126888 13058 126940 13064
rect 126612 4888 126664 4894
rect 126612 4830 126664 4836
rect 125508 4820 125560 4826
rect 125508 4762 125560 4768
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 82912 3460 82964 3466
rect 82912 3402 82964 3408
rect 108948 3460 109000 3466
rect 108948 3402 109000 3408
rect 1688 480 1716 3402
rect 126624 480 126652 4830
rect 126992 610 127020 14418
rect 128360 13184 128412 13190
rect 128360 13126 128412 13132
rect 128372 610 128400 13126
rect 129752 626 129780 15846
rect 126980 604 127032 610
rect 126980 546 127032 552
rect 127808 604 127860 610
rect 127808 546 127860 552
rect 128360 604 128412 610
rect 128360 546 128412 552
rect 129004 604 129056 610
rect 129752 598 130240 626
rect 131132 610 131160 21354
rect 131776 15910 131804 99418
rect 132420 42158 132448 102054
rect 132604 99414 132632 102068
rect 133432 100026 133460 102068
rect 133420 100020 133472 100026
rect 133420 99962 133472 99968
rect 134260 99414 134288 102068
rect 132592 99408 132644 99414
rect 132592 99350 132644 99356
rect 133788 99408 133840 99414
rect 133788 99350 133840 99356
rect 134248 99408 134300 99414
rect 134248 99350 134300 99356
rect 133800 77994 133828 99350
rect 135088 79354 135116 102068
rect 135930 102054 136588 102082
rect 135904 100088 135956 100094
rect 135904 100030 135956 100036
rect 135168 99408 135220 99414
rect 135168 99350 135220 99356
rect 135076 79348 135128 79354
rect 135076 79290 135128 79296
rect 133788 77988 133840 77994
rect 133788 77930 133840 77936
rect 135180 43450 135208 99350
rect 135168 43444 135220 43450
rect 135168 43386 135220 43392
rect 132408 42152 132460 42158
rect 132408 42094 132460 42100
rect 133880 28280 133932 28286
rect 133880 28222 133932 28228
rect 132592 17264 132644 17270
rect 132592 17206 132644 17212
rect 131764 15904 131816 15910
rect 131764 15846 131816 15852
rect 132604 7682 132632 17206
rect 133892 12442 133920 28222
rect 133880 12436 133932 12442
rect 133880 12378 133932 12384
rect 134800 12436 134852 12442
rect 134800 12378 134852 12384
rect 134812 12322 134840 12378
rect 134812 12294 134932 12322
rect 132592 7676 132644 7682
rect 132592 7618 132644 7624
rect 133788 7676 133840 7682
rect 133788 7618 133840 7624
rect 132592 4004 132644 4010
rect 132592 3946 132644 3952
rect 129004 546 129056 552
rect 127820 480 127848 546
rect 129016 480 129044 546
rect 130212 480 130240 598
rect 131120 604 131172 610
rect 131120 546 131172 552
rect 131396 604 131448 610
rect 131396 546 131448 552
rect 131408 480 131436 546
rect 132604 480 132632 3946
rect 133800 480 133828 7618
rect 134904 480 134932 12294
rect 135916 8702 135944 100030
rect 136560 17338 136588 102054
rect 136744 99414 136772 102068
rect 137586 102054 137876 102082
rect 136732 99408 136784 99414
rect 136732 99350 136784 99356
rect 137848 80714 137876 102054
rect 138400 99414 138428 102068
rect 137928 99408 137980 99414
rect 137928 99350 137980 99356
rect 138388 99408 138440 99414
rect 138388 99350 138440 99356
rect 137836 80708 137888 80714
rect 137836 80650 137888 80656
rect 137940 46306 137968 99350
rect 139228 47598 139256 102068
rect 140070 102054 140728 102082
rect 139308 99408 139360 99414
rect 139308 99350 139360 99356
rect 138020 47592 138072 47598
rect 138020 47534 138072 47540
rect 139216 47592 139268 47598
rect 139216 47534 139268 47540
rect 138032 46918 138060 47534
rect 138020 46912 138072 46918
rect 138020 46854 138072 46860
rect 137928 46300 137980 46306
rect 137928 46242 137980 46248
rect 138020 37324 138072 37330
rect 138020 37266 138072 37272
rect 138032 27606 138060 37266
rect 138020 27600 138072 27606
rect 138020 27542 138072 27548
rect 138480 27600 138532 27606
rect 138480 27542 138532 27548
rect 136640 18624 136692 18630
rect 136640 18566 136692 18572
rect 136548 17332 136600 17338
rect 136548 17274 136600 17280
rect 136652 12442 136680 18566
rect 136640 12436 136692 12442
rect 136640 12378 136692 12384
rect 137192 12436 137244 12442
rect 137192 12378 137244 12384
rect 137204 12322 137232 12378
rect 137204 12294 137324 12322
rect 135904 8696 135956 8702
rect 135904 8638 135956 8644
rect 136088 3936 136140 3942
rect 136088 3878 136140 3884
rect 136100 480 136128 3878
rect 137296 480 137324 12294
rect 138492 480 138520 27542
rect 139320 18630 139348 99350
rect 140700 82210 140728 102054
rect 140884 99414 140912 102068
rect 141726 102054 142016 102082
rect 140872 99408 140924 99414
rect 140872 99350 140924 99356
rect 140688 82204 140740 82210
rect 140688 82146 140740 82152
rect 141988 49026 142016 102054
rect 142540 99414 142568 102068
rect 143368 99498 143396 102068
rect 144210 102054 144868 102082
rect 143368 99470 143488 99498
rect 142068 99408 142120 99414
rect 142068 99350 142120 99356
rect 142528 99408 142580 99414
rect 142528 99350 142580 99356
rect 143356 99408 143408 99414
rect 143356 99350 143408 99356
rect 140780 49020 140832 49026
rect 140780 48962 140832 48968
rect 141976 49020 142028 49026
rect 141976 48962 142028 48968
rect 139308 18624 139360 18630
rect 139308 18566 139360 18572
rect 140792 7682 140820 48962
rect 142080 20058 142108 99350
rect 143368 86290 143396 99350
rect 143356 86284 143408 86290
rect 143356 86226 143408 86232
rect 143460 21418 143488 99470
rect 144840 50454 144868 102054
rect 145024 99414 145052 102068
rect 145012 99408 145064 99414
rect 145012 99350 145064 99356
rect 145852 98666 145880 102068
rect 146680 99414 146708 102068
rect 146116 99408 146168 99414
rect 146116 99350 146168 99356
rect 146668 99408 146720 99414
rect 146668 99350 146720 99356
rect 145840 98660 145892 98666
rect 145840 98602 145892 98608
rect 146128 87718 146156 99350
rect 147508 93158 147536 102068
rect 148350 102054 149008 102082
rect 147588 99408 147640 99414
rect 147588 99350 147640 99356
rect 147496 93152 147548 93158
rect 147496 93094 147548 93100
rect 146116 87712 146168 87718
rect 146116 87654 146168 87660
rect 147600 51746 147628 99350
rect 144920 51740 144972 51746
rect 144920 51682 144972 51688
rect 147588 51740 147640 51746
rect 147588 51682 147640 51688
rect 144828 50448 144880 50454
rect 144828 50390 144880 50396
rect 143540 22772 143592 22778
rect 143540 22714 143592 22720
rect 143448 21412 143500 21418
rect 143448 21354 143500 21360
rect 142068 20052 142120 20058
rect 142068 19994 142120 20000
rect 140872 19984 140924 19990
rect 140872 19926 140924 19932
rect 140780 7676 140832 7682
rect 140780 7618 140832 7624
rect 139676 3868 139728 3874
rect 139676 3810 139728 3816
rect 139688 480 139716 3810
rect 140884 480 140912 19926
rect 143552 12442 143580 22714
rect 144932 12442 144960 51682
rect 147680 24132 147732 24138
rect 147680 24074 147732 24080
rect 143540 12436 143592 12442
rect 143540 12378 143592 12384
rect 144460 12436 144512 12442
rect 144460 12378 144512 12384
rect 144920 12436 144972 12442
rect 144920 12378 144972 12384
rect 145656 12436 145708 12442
rect 145656 12378 145708 12384
rect 142068 7676 142120 7682
rect 142068 7618 142120 7624
rect 142080 480 142108 7618
rect 143264 3800 143316 3806
rect 143264 3742 143316 3748
rect 143276 480 143304 3742
rect 144472 480 144500 12378
rect 144920 4820 144972 4826
rect 144920 4762 144972 4768
rect 145012 4820 145064 4826
rect 145012 4762 145064 4768
rect 144932 4706 144960 4762
rect 145024 4706 145052 4762
rect 144932 4678 145052 4706
rect 145668 480 145696 12378
rect 146852 3732 146904 3738
rect 146852 3674 146904 3680
rect 146864 480 146892 3674
rect 147692 3380 147720 24074
rect 148980 22778 149008 102054
rect 149164 99754 149192 102068
rect 149152 99748 149204 99754
rect 149152 99690 149204 99696
rect 149992 95946 150020 102068
rect 150728 99754 150756 102068
rect 151464 102054 151570 102082
rect 150348 99748 150400 99754
rect 150348 99690 150400 99696
rect 150716 99748 150768 99754
rect 150716 99690 150768 99696
rect 149980 95940 150032 95946
rect 149980 95882 150032 95888
rect 150360 53106 150388 99690
rect 151464 96665 151492 102054
rect 152384 100162 152412 102068
rect 153212 100706 153240 102068
rect 154054 102054 154436 102082
rect 153200 100700 153252 100706
rect 153200 100642 153252 100648
rect 152372 100156 152424 100162
rect 152372 100098 152424 100104
rect 153108 100156 153160 100162
rect 153108 100098 153160 100104
rect 151728 99748 151780 99754
rect 151728 99690 151780 99696
rect 151450 96656 151506 96665
rect 151450 96591 151506 96600
rect 151634 96656 151690 96665
rect 151634 96591 151690 96600
rect 151648 89758 151676 96591
rect 151452 89752 151504 89758
rect 151636 89752 151688 89758
rect 151504 89700 151636 89706
rect 151452 89694 151688 89700
rect 151464 89678 151676 89694
rect 151648 80209 151676 89678
rect 151634 80200 151690 80209
rect 151634 80135 151690 80144
rect 151542 77344 151598 77353
rect 151542 77279 151598 77288
rect 151556 77246 151584 77279
rect 151544 77240 151596 77246
rect 151544 77182 151596 77188
rect 151636 67652 151688 67658
rect 151636 67594 151688 67600
rect 151648 67522 151676 67594
rect 151452 67516 151504 67522
rect 151452 67458 151504 67464
rect 151636 67516 151688 67522
rect 151636 67458 151688 67464
rect 151464 54602 151492 67458
rect 151452 54596 151504 54602
rect 151452 54538 151504 54544
rect 149060 53100 149112 53106
rect 149060 53042 149112 53048
rect 150348 53100 150400 53106
rect 150348 53042 150400 53048
rect 148968 22772 149020 22778
rect 148968 22714 149020 22720
rect 149072 3380 149100 53042
rect 150532 25560 150584 25566
rect 150532 25502 150584 25508
rect 150440 3596 150492 3602
rect 150440 3538 150492 3544
rect 147692 3352 148088 3380
rect 149072 3352 149284 3380
rect 148060 480 148088 3352
rect 149256 480 149284 3352
rect 150452 480 150480 3538
rect 150544 3380 150572 25502
rect 151740 24138 151768 99690
rect 153120 91866 153148 100098
rect 153108 91860 153160 91866
rect 153108 91802 153160 91808
rect 154408 55894 154436 102054
rect 154868 100706 154896 102068
rect 155710 102054 155908 102082
rect 156538 102054 157288 102082
rect 154488 100700 154540 100706
rect 154488 100642 154540 100648
rect 154856 100700 154908 100706
rect 154856 100642 154908 100648
rect 155776 100700 155828 100706
rect 155776 100642 155828 100648
rect 151820 55888 151872 55894
rect 151820 55830 151872 55836
rect 154396 55888 154448 55894
rect 154396 55830 154448 55836
rect 151728 24132 151780 24138
rect 151728 24074 151780 24080
rect 151832 3482 151860 55830
rect 154500 25566 154528 100642
rect 155788 90438 155816 100642
rect 155776 90432 155828 90438
rect 155776 90374 155828 90380
rect 155880 26926 155908 102054
rect 157260 57254 157288 102054
rect 157352 99414 157380 102068
rect 158194 102054 158668 102082
rect 157340 99408 157392 99414
rect 157340 99350 157392 99356
rect 158536 99408 158588 99414
rect 158536 99350 158588 99356
rect 158548 89078 158576 99350
rect 158536 89072 158588 89078
rect 158536 89014 158588 89020
rect 155960 57248 156012 57254
rect 155960 57190 156012 57196
rect 157248 57248 157300 57254
rect 157248 57190 157300 57196
rect 154580 26920 154632 26926
rect 154580 26862 154632 26868
rect 155868 26920 155920 26926
rect 155868 26862 155920 26868
rect 154488 25560 154540 25566
rect 154488 25502 154540 25508
rect 153936 3664 153988 3670
rect 153936 3606 153988 3612
rect 151832 3454 152780 3482
rect 150544 3352 151584 3380
rect 151556 480 151584 3352
rect 152752 480 152780 3454
rect 153948 480 153976 3606
rect 154592 3482 154620 26862
rect 155972 3482 156000 57190
rect 158640 28286 158668 102054
rect 159008 99414 159036 102068
rect 159850 102054 160048 102082
rect 158996 99408 159048 99414
rect 158996 99350 159048 99356
rect 159916 99408 159968 99414
rect 159916 99350 159968 99356
rect 159928 58682 159956 99350
rect 158720 58676 158772 58682
rect 158720 58618 158772 58624
rect 159916 58676 159968 58682
rect 159916 58618 159968 58624
rect 158628 28280 158680 28286
rect 158628 28222 158680 28228
rect 158732 3534 158760 58618
rect 160020 42090 160048 102054
rect 160664 99414 160692 102068
rect 161492 99414 161520 102068
rect 162334 102054 162808 102082
rect 160652 99408 160704 99414
rect 160652 99350 160704 99356
rect 161388 99408 161440 99414
rect 161388 99350 161440 99356
rect 161480 99408 161532 99414
rect 161480 99350 161532 99356
rect 162676 99408 162728 99414
rect 162676 99350 162728 99356
rect 160008 42084 160060 42090
rect 160008 42026 160060 42032
rect 158812 29640 158864 29646
rect 158812 29582 158864 29588
rect 157524 3528 157576 3534
rect 154592 3454 155172 3482
rect 155972 3454 156368 3482
rect 157524 3470 157576 3476
rect 158720 3528 158772 3534
rect 158720 3470 158772 3476
rect 155144 480 155172 3454
rect 156340 480 156368 3454
rect 157536 480 157564 3470
rect 158824 1442 158852 29582
rect 161400 6254 161428 99350
rect 162688 60042 162716 99350
rect 162676 60036 162728 60042
rect 162676 59978 162728 59984
rect 162780 38078 162808 102054
rect 163148 97374 163176 102068
rect 163976 99414 164004 102068
rect 164804 99482 164832 102068
rect 165632 100162 165660 102068
rect 166474 102054 166948 102082
rect 165620 100156 165672 100162
rect 165620 100098 165672 100104
rect 164792 99476 164844 99482
rect 164792 99418 164844 99424
rect 163964 99408 164016 99414
rect 163964 99350 164016 99356
rect 164884 99408 164936 99414
rect 164884 99350 164936 99356
rect 163136 97368 163188 97374
rect 163136 97310 163188 97316
rect 164240 61396 164292 61402
rect 164240 61338 164292 61344
rect 162768 38072 162820 38078
rect 162768 38014 162820 38020
rect 162860 31068 162912 31074
rect 162860 31010 162912 31016
rect 161388 6248 161440 6254
rect 161388 6190 161440 6196
rect 162308 3936 162360 3942
rect 162308 3878 162360 3884
rect 159916 3528 159968 3534
rect 159916 3470 159968 3476
rect 158732 1414 158852 1442
rect 158732 480 158760 1414
rect 159928 480 159956 3470
rect 161112 3460 161164 3466
rect 161112 3402 161164 3408
rect 161124 480 161152 3402
rect 162320 480 162348 3878
rect 162872 3482 162900 31010
rect 164252 3482 164280 61338
rect 164896 44878 164924 99350
rect 166920 61470 166948 102054
rect 167288 99414 167316 102068
rect 168130 102054 168328 102082
rect 167276 99408 167328 99414
rect 167276 99350 167328 99356
rect 168196 99408 168248 99414
rect 168196 99350 168248 99356
rect 167000 62824 167052 62830
rect 167000 62766 167052 62772
rect 166908 61464 166960 61470
rect 166908 61406 166960 61412
rect 164884 44872 164936 44878
rect 164884 44814 164936 44820
rect 165896 6180 165948 6186
rect 165896 6122 165948 6128
rect 162872 3454 163544 3482
rect 164252 3454 164740 3482
rect 163516 480 163544 3454
rect 164712 480 164740 3454
rect 165908 480 165936 6122
rect 167012 3534 167040 62766
rect 168208 43518 168236 99350
rect 168196 43512 168248 43518
rect 168196 43454 168248 43460
rect 167092 32428 167144 32434
rect 167092 32370 167144 32376
rect 167000 3528 167052 3534
rect 167000 3470 167052 3476
rect 167104 480 167132 32370
rect 168300 29646 168328 102054
rect 168944 99414 168972 102068
rect 169024 99476 169076 99482
rect 169024 99418 169076 99424
rect 168932 99408 168984 99414
rect 168932 99350 168984 99356
rect 169036 46238 169064 99418
rect 169772 99414 169800 102068
rect 170614 102054 171088 102082
rect 169668 99408 169720 99414
rect 169668 99350 169720 99356
rect 169760 99408 169812 99414
rect 169760 99350 169812 99356
rect 170956 99408 171008 99414
rect 170956 99350 171008 99356
rect 169680 62830 169708 99350
rect 169668 62824 169720 62830
rect 169668 62766 169720 62772
rect 170968 47666 170996 99350
rect 170956 47660 171008 47666
rect 170956 47602 171008 47608
rect 169024 46232 169076 46238
rect 169024 46174 169076 46180
rect 168380 44940 168432 44946
rect 168380 44882 168432 44888
rect 168288 29640 168340 29646
rect 168288 29582 168340 29588
rect 168196 3528 168248 3534
rect 168196 3470 168248 3476
rect 168392 3482 168420 44882
rect 169760 33788 169812 33794
rect 169760 33730 169812 33736
rect 169772 3482 169800 33730
rect 171060 9110 171088 102054
rect 171428 99414 171456 102068
rect 172256 100094 172284 102068
rect 172244 100088 172296 100094
rect 172244 100030 172296 100036
rect 173084 99414 173112 102068
rect 173728 102054 173834 102082
rect 174662 102054 175228 102082
rect 171416 99408 171468 99414
rect 171416 99350 171468 99356
rect 172428 99408 172480 99414
rect 172428 99350 172480 99356
rect 173072 99408 173124 99414
rect 173072 99350 173124 99356
rect 172440 64190 172468 99350
rect 173728 65618 173756 102054
rect 174544 100156 174596 100162
rect 174544 100098 174596 100104
rect 173808 99408 173860 99414
rect 173808 99350 173860 99356
rect 173716 65612 173768 65618
rect 173716 65554 173768 65560
rect 171140 64184 171192 64190
rect 171140 64126 171192 64132
rect 172428 64184 172480 64190
rect 172428 64126 172480 64132
rect 171048 9104 171100 9110
rect 171048 9046 171100 9052
rect 171152 3482 171180 64126
rect 173820 31074 173848 99350
rect 173900 35216 173952 35222
rect 173900 35158 173952 35164
rect 173808 31068 173860 31074
rect 173808 31010 173860 31016
rect 172980 7608 173032 7614
rect 172980 7550 173032 7556
rect 168208 480 168236 3470
rect 168392 3454 169432 3482
rect 169772 3454 170628 3482
rect 171152 3454 171824 3482
rect 169404 480 169432 3454
rect 170600 480 170628 3454
rect 171796 480 171824 3454
rect 172992 480 173020 7550
rect 173912 3482 173940 35158
rect 174556 7750 174584 100098
rect 175200 82142 175228 102054
rect 175476 99414 175504 102068
rect 176318 102054 176516 102082
rect 177146 102054 177896 102082
rect 175464 99408 175516 99414
rect 175464 99350 175516 99356
rect 175188 82136 175240 82142
rect 175188 82078 175240 82084
rect 176488 66978 176516 102054
rect 176568 99408 176620 99414
rect 176568 99350 176620 99356
rect 176476 66972 176528 66978
rect 176476 66914 176528 66920
rect 175280 66904 175332 66910
rect 175280 66846 175332 66852
rect 174544 7744 174596 7750
rect 174544 7686 174596 7692
rect 175292 3482 175320 66846
rect 176580 32434 176608 99350
rect 177868 50386 177896 102054
rect 177856 50380 177908 50386
rect 177856 50322 177908 50328
rect 176660 36576 176712 36582
rect 176660 36518 176712 36524
rect 176568 32428 176620 32434
rect 176568 32370 176620 32376
rect 176568 8968 176620 8974
rect 176568 8910 176620 8916
rect 173912 3454 174216 3482
rect 175292 3454 175412 3482
rect 174188 480 174216 3454
rect 175384 480 175412 3454
rect 176580 480 176608 8910
rect 176672 3482 176700 36518
rect 177960 33794 177988 102068
rect 178802 102054 179368 102082
rect 178684 100020 178736 100026
rect 178684 99962 178736 99968
rect 178040 68332 178092 68338
rect 178040 68274 178092 68280
rect 177948 33788 178000 33794
rect 177948 33730 178000 33736
rect 178052 3618 178080 68274
rect 178696 4894 178724 99962
rect 179340 68406 179368 102054
rect 179616 99414 179644 102068
rect 180444 100162 180472 102068
rect 180432 100156 180484 100162
rect 180432 100098 180484 100104
rect 181272 99414 181300 102068
rect 179604 99408 179656 99414
rect 179604 99350 179656 99356
rect 180708 99408 180760 99414
rect 180708 99350 180760 99356
rect 181260 99408 181312 99414
rect 181260 99350 181312 99356
rect 179328 68400 179380 68406
rect 179328 68342 179380 68348
rect 180720 51814 180748 99350
rect 182100 53174 182128 102068
rect 182942 102054 183508 102082
rect 182824 99408 182876 99414
rect 182824 99350 182876 99356
rect 182836 69834 182864 99350
rect 182824 69828 182876 69834
rect 182824 69770 182876 69776
rect 182180 69692 182232 69698
rect 182180 69634 182232 69640
rect 182088 53168 182140 53174
rect 182088 53110 182140 53116
rect 180708 51808 180760 51814
rect 180708 51750 180760 51756
rect 180800 37936 180852 37942
rect 180800 37878 180852 37884
rect 179420 10328 179472 10334
rect 179420 10270 179472 10276
rect 178684 4888 178736 4894
rect 178684 4830 178736 4836
rect 178052 3590 179000 3618
rect 176672 3454 177804 3482
rect 177776 480 177804 3454
rect 178972 480 179000 3590
rect 179432 3482 179460 10270
rect 180812 3482 180840 37878
rect 182192 3482 182220 69634
rect 183480 10402 183508 102054
rect 183756 99482 183784 102068
rect 184598 102054 184888 102082
rect 183744 99476 183796 99482
rect 183744 99418 183796 99424
rect 184860 39438 184888 102054
rect 185412 99414 185440 102068
rect 186148 102054 186254 102082
rect 187082 102054 187648 102082
rect 185400 99408 185452 99414
rect 185400 99350 185452 99356
rect 186148 72554 186176 102054
rect 186964 99476 187016 99482
rect 186964 99418 187016 99424
rect 186228 99408 186280 99414
rect 186228 99350 186280 99356
rect 186136 72548 186188 72554
rect 186136 72490 186188 72496
rect 184940 71052 184992 71058
rect 184940 70994 184992 71000
rect 184848 39432 184900 39438
rect 184848 39374 184900 39380
rect 183560 11756 183612 11762
rect 183560 11698 183612 11704
rect 183468 10396 183520 10402
rect 183468 10338 183520 10344
rect 183572 3482 183600 11698
rect 184848 4820 184900 4826
rect 184848 4762 184900 4768
rect 179432 3454 180196 3482
rect 180812 3454 181392 3482
rect 182192 3454 182588 3482
rect 183572 3454 183784 3482
rect 180168 480 180196 3454
rect 181364 480 181392 3454
rect 182560 480 182588 3454
rect 183756 480 183784 3454
rect 184860 480 184888 4762
rect 184952 3482 184980 70994
rect 186240 11898 186268 99350
rect 186976 71126 187004 99418
rect 187620 87650 187648 102054
rect 187896 99414 187924 102068
rect 188738 102054 188936 102082
rect 187884 99408 187936 99414
rect 187884 99350 187936 99356
rect 187608 87644 187660 87650
rect 187608 87586 187660 87592
rect 188908 73914 188936 102054
rect 189552 99414 189580 102068
rect 188988 99408 189040 99414
rect 188988 99350 189040 99356
rect 189540 99408 189592 99414
rect 189540 99350 189592 99356
rect 188896 73908 188948 73914
rect 188896 73850 188948 73856
rect 186964 71120 187016 71126
rect 186964 71062 187016 71068
rect 187700 39364 187752 39370
rect 187700 39306 187752 39312
rect 186320 13116 186372 13122
rect 186320 13058 186372 13064
rect 186228 11892 186280 11898
rect 186228 11834 186280 11840
rect 186332 3482 186360 13058
rect 187712 3482 187740 39306
rect 189000 13190 189028 99350
rect 189080 75200 189132 75206
rect 189080 75142 189132 75148
rect 188988 13184 189040 13190
rect 188988 13126 189040 13132
rect 189092 3482 189120 75142
rect 190380 35290 190408 102068
rect 191222 102054 191788 102082
rect 191104 99408 191156 99414
rect 191104 99350 191156 99356
rect 191116 55962 191144 99350
rect 191760 75274 191788 102054
rect 192036 99414 192064 102068
rect 192878 102054 193168 102082
rect 193706 102054 194456 102082
rect 192024 99408 192076 99414
rect 192024 99350 192076 99356
rect 193036 99408 193088 99414
rect 193036 99350 193088 99356
rect 191748 75268 191800 75274
rect 191748 75210 191800 75216
rect 193048 57322 193076 99350
rect 193036 57316 193088 57322
rect 193036 57258 193088 57264
rect 191104 55956 191156 55962
rect 191104 55898 191156 55904
rect 191840 40724 191892 40730
rect 191840 40666 191892 40672
rect 190368 35284 190420 35290
rect 190368 35226 190420 35232
rect 190460 14476 190512 14482
rect 190460 14418 190512 14424
rect 190472 3482 190500 14418
rect 191852 3482 191880 40666
rect 193140 14550 193168 102054
rect 194428 76566 194456 102054
rect 193220 76560 193272 76566
rect 193220 76502 193272 76508
rect 194416 76560 194468 76566
rect 194416 76502 194468 76508
rect 193128 14544 193180 14550
rect 193128 14486 193180 14492
rect 184952 3454 186084 3482
rect 186332 3454 187280 3482
rect 187712 3454 188476 3482
rect 189092 3454 189672 3482
rect 190472 3454 190868 3482
rect 191852 3454 192064 3482
rect 186056 480 186084 3454
rect 187252 480 187280 3454
rect 188448 480 188476 3454
rect 189644 480 189672 3454
rect 190840 480 190868 3454
rect 192036 480 192064 3454
rect 193232 480 193260 76502
rect 194520 54534 194548 102068
rect 195362 102054 195928 102082
rect 194508 54528 194560 54534
rect 194508 54470 194560 54476
rect 194600 42152 194652 42158
rect 194600 42094 194652 42100
rect 193312 15904 193364 15910
rect 193312 15846 193364 15852
rect 193324 3482 193352 15846
rect 194612 3482 194640 42094
rect 195900 15978 195928 102054
rect 196084 94518 196112 102068
rect 196926 102054 197308 102082
rect 196072 94512 196124 94518
rect 196072 94454 196124 94460
rect 195980 77988 196032 77994
rect 195980 77930 196032 77936
rect 195888 15972 195940 15978
rect 195888 15914 195940 15920
rect 195992 12442 196020 77930
rect 197280 49094 197308 102054
rect 197740 100026 197768 102068
rect 197728 100020 197780 100026
rect 197728 99962 197780 99968
rect 198004 95260 198056 95266
rect 198004 95202 198056 95208
rect 198016 95130 198044 95202
rect 198004 95124 198056 95130
rect 198004 95066 198056 95072
rect 198568 89758 198596 102068
rect 199410 102054 200068 102082
rect 198556 89752 198608 89758
rect 198556 89694 198608 89700
rect 198096 85604 198148 85610
rect 198096 85546 198148 85552
rect 198556 85604 198608 85610
rect 198556 85546 198608 85552
rect 198108 80238 198136 85546
rect 198096 80232 198148 80238
rect 198096 80174 198148 80180
rect 198568 78062 198596 85546
rect 198556 78056 198608 78062
rect 198556 77998 198608 78004
rect 198004 75948 198056 75954
rect 198004 75890 198056 75896
rect 198016 67561 198044 75890
rect 197726 67552 197782 67561
rect 197726 67487 197782 67496
rect 198002 67552 198058 67561
rect 198002 67487 198058 67496
rect 197740 58002 197768 67487
rect 200040 61402 200068 102054
rect 200224 99754 200252 102068
rect 201066 102054 201356 102082
rect 200212 99748 200264 99754
rect 200212 99690 200264 99696
rect 201328 79422 201356 102054
rect 201880 100706 201908 102068
rect 201868 100700 201920 100706
rect 201868 100642 201920 100648
rect 201408 99748 201460 99754
rect 201408 99690 201460 99696
rect 201316 79416 201368 79422
rect 201316 79358 201368 79364
rect 200120 79348 200172 79354
rect 200120 79290 200172 79296
rect 200132 66230 200160 79290
rect 200120 66224 200172 66230
rect 200120 66166 200172 66172
rect 200028 61396 200080 61402
rect 200028 61338 200080 61344
rect 197728 57996 197780 58002
rect 197728 57938 197780 57944
rect 198004 57996 198056 58002
rect 198004 57938 198056 57944
rect 197268 49088 197320 49094
rect 197268 49030 197320 49036
rect 198016 31754 198044 57938
rect 200120 56636 200172 56642
rect 200120 56578 200172 56584
rect 200132 46918 200160 56578
rect 200120 46912 200172 46918
rect 200120 46854 200172 46860
rect 198740 43444 198792 43450
rect 198740 43386 198792 43392
rect 198752 38622 198780 43386
rect 198556 38616 198608 38622
rect 198556 38558 198608 38564
rect 198740 38616 198792 38622
rect 198740 38558 198792 38564
rect 198004 31748 198056 31754
rect 198004 31690 198056 31696
rect 198188 31748 198240 31754
rect 198188 31690 198240 31696
rect 198200 28966 198228 31690
rect 198568 29073 198596 38558
rect 200120 37324 200172 37330
rect 200120 37266 200172 37272
rect 198554 29064 198610 29073
rect 198554 28999 198610 29008
rect 198738 29064 198794 29073
rect 198738 28999 198794 29008
rect 198188 28960 198240 28966
rect 198188 28902 198240 28908
rect 198752 27606 198780 28999
rect 198740 27600 198792 27606
rect 198740 27542 198792 27548
rect 200132 22846 200160 37266
rect 200120 22840 200172 22846
rect 200120 22782 200172 22788
rect 198096 19372 198148 19378
rect 198096 19314 198148 19320
rect 198108 12458 198136 19314
rect 201420 17270 201448 99690
rect 202708 99482 202736 102068
rect 203550 102054 204208 102082
rect 202788 100700 202840 100706
rect 202788 100642 202840 100648
rect 202696 99476 202748 99482
rect 202696 99418 202748 99424
rect 202800 62898 202828 100642
rect 203524 100156 203576 100162
rect 203524 100098 203576 100104
rect 202880 80708 202932 80714
rect 202880 80650 202932 80656
rect 202788 62892 202840 62898
rect 202788 62834 202840 62840
rect 201500 46300 201552 46306
rect 201500 46242 201552 46248
rect 201408 17264 201460 17270
rect 201408 17206 201460 17212
rect 195980 12436 196032 12442
rect 195980 12378 196032 12384
rect 196808 12436 196860 12442
rect 198108 12430 198228 12458
rect 196808 12378 196860 12384
rect 193324 3454 194456 3482
rect 194612 3454 195652 3482
rect 194428 480 194456 3454
rect 195624 480 195652 3454
rect 196820 480 196848 12378
rect 198200 4894 198228 12430
rect 199200 9716 199252 9722
rect 199200 9658 199252 9664
rect 200396 9716 200448 9722
rect 200396 9658 200448 9664
rect 198004 4888 198056 4894
rect 198004 4830 198056 4836
rect 198188 4888 198240 4894
rect 198188 4830 198240 4836
rect 198016 480 198044 4830
rect 199212 480 199240 9658
rect 200408 9602 200436 9658
rect 200408 9574 200528 9602
rect 200500 610 200528 9574
rect 201512 7614 201540 46242
rect 201592 17332 201644 17338
rect 201592 17274 201644 17280
rect 201500 7608 201552 7614
rect 201500 7550 201552 7556
rect 201604 7426 201632 17274
rect 202892 12442 202920 80650
rect 202880 12436 202932 12442
rect 202880 12378 202932 12384
rect 202696 7608 202748 7614
rect 202696 7550 202748 7556
rect 201512 7398 201632 7426
rect 200396 604 200448 610
rect 200396 546 200448 552
rect 200488 604 200540 610
rect 200488 546 200540 552
rect 200408 480 200436 546
rect 201512 480 201540 7398
rect 202708 480 202736 7550
rect 203536 4826 203564 100098
rect 204180 80714 204208 102054
rect 204364 100706 204392 102068
rect 205206 102054 205588 102082
rect 204352 100700 204404 100706
rect 204352 100642 204404 100648
rect 205456 100700 205508 100706
rect 205456 100642 205508 100648
rect 204168 80708 204220 80714
rect 204168 80650 204220 80656
rect 205468 64258 205496 100642
rect 205456 64252 205508 64258
rect 205456 64194 205508 64200
rect 205560 19990 205588 102054
rect 206020 99414 206048 102068
rect 206848 99498 206876 102068
rect 207690 102054 208348 102082
rect 206848 99470 206968 99498
rect 206008 99408 206060 99414
rect 206008 99350 206060 99356
rect 206836 99408 206888 99414
rect 206836 99350 206888 99356
rect 206848 83502 206876 99350
rect 206836 83496 206888 83502
rect 206836 83438 206888 83444
rect 206940 65550 206968 99470
rect 207664 99476 207716 99482
rect 207664 99418 207716 99424
rect 207020 82204 207072 82210
rect 207020 82146 207072 82152
rect 206928 65544 206980 65550
rect 206928 65486 206980 65492
rect 205640 47592 205692 47598
rect 205640 47534 205692 47540
rect 205548 19984 205600 19990
rect 205548 19926 205600 19932
rect 204260 18624 204312 18630
rect 204260 18566 204312 18572
rect 204272 12442 204300 18566
rect 203892 12436 203944 12442
rect 203892 12378 203944 12384
rect 204260 12436 204312 12442
rect 204260 12378 204312 12384
rect 205088 12436 205140 12442
rect 205088 12378 205140 12384
rect 203524 4820 203576 4826
rect 203524 4762 203576 4768
rect 203904 480 203932 12378
rect 205100 480 205128 12378
rect 205652 3346 205680 47534
rect 207032 3346 207060 82146
rect 207676 18630 207704 99418
rect 208320 21486 208348 102054
rect 208504 99414 208532 102068
rect 209346 102054 209728 102082
rect 208492 99408 208544 99414
rect 208492 99350 208544 99356
rect 209596 99408 209648 99414
rect 209596 99350 209648 99356
rect 209608 84862 209636 99350
rect 209596 84856 209648 84862
rect 209596 84798 209648 84804
rect 209700 69766 209728 102054
rect 210160 99414 210188 102068
rect 210988 99498 211016 102068
rect 211830 102054 212488 102082
rect 210988 99470 211108 99498
rect 210148 99408 210200 99414
rect 210148 99350 210200 99356
rect 210976 99408 211028 99414
rect 210976 99350 211028 99356
rect 210988 89010 211016 99350
rect 210976 89004 211028 89010
rect 210976 88946 211028 88952
rect 211080 86290 211108 99470
rect 209780 86284 209832 86290
rect 209780 86226 209832 86232
rect 211068 86284 211120 86290
rect 211068 86226 211120 86232
rect 209688 69760 209740 69766
rect 209688 69702 209740 69708
rect 208308 21480 208360 21486
rect 208308 21422 208360 21428
rect 208400 20052 208452 20058
rect 208400 19994 208452 20000
rect 207664 18624 207716 18630
rect 207664 18566 207716 18572
rect 208412 3346 208440 19994
rect 209792 3534 209820 86226
rect 212460 66910 212488 102054
rect 212644 99414 212672 102068
rect 213486 102054 213776 102082
rect 212632 99408 212684 99414
rect 212632 99350 212684 99356
rect 213748 90370 213776 102054
rect 214300 99414 214328 102068
rect 213828 99408 213880 99414
rect 213828 99350 213880 99356
rect 214288 99408 214340 99414
rect 214288 99350 214340 99356
rect 213736 90364 213788 90370
rect 213736 90306 213788 90312
rect 212448 66904 212500 66910
rect 212448 66846 212500 66852
rect 212540 50448 212592 50454
rect 212540 50390 212592 50396
rect 209872 49020 209924 49026
rect 209872 48962 209924 48968
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 205652 3318 206324 3346
rect 207032 3318 207520 3346
rect 208412 3318 208716 3346
rect 206296 480 206324 3318
rect 207492 480 207520 3318
rect 208688 480 208716 3318
rect 209884 480 209912 48962
rect 211160 21412 211212 21418
rect 211160 21354 211212 21360
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 211172 3482 211200 21354
rect 212552 3482 212580 50390
rect 213840 36582 213868 99350
rect 215128 93786 215156 102068
rect 215970 102054 216628 102082
rect 215944 99408 215996 99414
rect 215944 99350 215996 99356
rect 215300 98660 215352 98666
rect 215300 98602 215352 98608
rect 215128 93758 215248 93786
rect 213920 87712 213972 87718
rect 213920 87654 213972 87660
rect 213828 36576 213880 36582
rect 213828 36518 213880 36524
rect 213932 3482 213960 87654
rect 215220 80050 215248 93758
rect 215036 80022 215248 80050
rect 215036 74526 215064 80022
rect 215024 74520 215076 74526
rect 215024 74462 215076 74468
rect 215208 74520 215260 74526
rect 215208 74462 215260 74468
rect 215220 64977 215248 74462
rect 215022 64968 215078 64977
rect 214944 64926 215022 64954
rect 214944 63510 214972 64926
rect 215022 64903 215078 64912
rect 215206 64968 215262 64977
rect 215206 64903 215262 64912
rect 214932 63504 214984 63510
rect 214932 63446 214984 63452
rect 215024 63504 215076 63510
rect 215024 63446 215076 63452
rect 215036 60761 215064 63446
rect 215022 60752 215078 60761
rect 215022 60687 215078 60696
rect 215022 48376 215078 48385
rect 214944 48334 215022 48362
rect 214944 41478 214972 48334
rect 215022 48311 215078 48320
rect 214932 41472 214984 41478
rect 214932 41414 214984 41420
rect 215024 41336 215076 41342
rect 215024 41278 215076 41284
rect 215036 37262 215064 41278
rect 215024 37256 215076 37262
rect 215024 37198 215076 37204
rect 215116 27668 215168 27674
rect 215116 27610 215168 27616
rect 215128 22846 215156 27610
rect 215116 22840 215168 22846
rect 215116 22782 215168 22788
rect 215312 3482 215340 98602
rect 215956 68338 215984 99350
rect 216600 91798 216628 102054
rect 216784 99414 216812 102068
rect 217612 100162 217640 102068
rect 217600 100156 217652 100162
rect 217600 100098 217652 100104
rect 218440 99414 218468 102068
rect 219190 102054 219388 102082
rect 220018 102054 220768 102082
rect 216772 99408 216824 99414
rect 216772 99350 216824 99356
rect 217968 99408 218020 99414
rect 217968 99350 218020 99356
rect 218428 99408 218480 99414
rect 218428 99350 218480 99356
rect 219256 99408 219308 99414
rect 219256 99350 219308 99356
rect 216588 91792 216640 91798
rect 216588 91734 216640 91740
rect 215944 68332 215996 68338
rect 215944 68274 215996 68280
rect 216680 51740 216732 51746
rect 216680 51682 216732 51688
rect 216692 3482 216720 51682
rect 217980 21418 218008 99350
rect 219268 93158 219296 99350
rect 218060 93152 218112 93158
rect 218060 93094 218112 93100
rect 219256 93152 219308 93158
rect 219256 93094 219308 93100
rect 217968 21412 218020 21418
rect 217968 21354 218020 21360
rect 218072 3482 218100 93094
rect 219360 71058 219388 102054
rect 219348 71052 219400 71058
rect 219348 70994 219400 71000
rect 219440 53100 219492 53106
rect 219440 53042 219492 53048
rect 218152 22772 218204 22778
rect 218152 22714 218204 22720
rect 218164 3602 218192 22714
rect 218152 3596 218204 3602
rect 218152 3538 218204 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 211080 480 211108 3470
rect 211172 3454 212304 3482
rect 212552 3454 213500 3482
rect 213932 3454 214696 3482
rect 215312 3454 215892 3482
rect 216692 3454 217088 3482
rect 218072 3454 218192 3482
rect 212276 480 212304 3454
rect 213472 480 213500 3454
rect 214668 480 214696 3454
rect 215864 480 215892 3454
rect 217060 480 217088 3454
rect 218164 480 218192 3454
rect 219360 480 219388 3538
rect 219452 3482 219480 53042
rect 220740 38010 220768 102054
rect 220832 99414 220860 102068
rect 221660 100094 221688 102068
rect 221648 100088 221700 100094
rect 221648 100030 221700 100036
rect 222488 99414 222516 102068
rect 223330 102054 223528 102082
rect 220820 99408 220872 99414
rect 220820 99350 220872 99356
rect 222108 99408 222160 99414
rect 222108 99350 222160 99356
rect 222476 99408 222528 99414
rect 222476 99350 222528 99356
rect 223396 99408 223448 99414
rect 223396 99350 223448 99356
rect 220820 95940 220872 95946
rect 220820 95882 220872 95888
rect 220728 38004 220780 38010
rect 220728 37946 220780 37952
rect 220832 3482 220860 95882
rect 222120 7682 222148 99350
rect 223408 39370 223436 99350
rect 223396 39364 223448 39370
rect 223396 39306 223448 39312
rect 222200 24132 222252 24138
rect 222200 24074 222252 24080
rect 222108 7676 222160 7682
rect 222108 7618 222160 7624
rect 222212 3482 222240 24074
rect 223500 9042 223528 102054
rect 224144 99414 224172 102068
rect 224224 100156 224276 100162
rect 224224 100098 224276 100104
rect 224132 99408 224184 99414
rect 224132 99350 224184 99356
rect 223580 54596 223632 54602
rect 223580 54538 223632 54544
rect 223488 9036 223540 9042
rect 223488 8978 223540 8984
rect 223592 3482 223620 54538
rect 224236 24206 224264 100098
rect 224972 99414 225000 102068
rect 224868 99408 224920 99414
rect 224868 99350 224920 99356
rect 224960 99408 225012 99414
rect 224960 99350 225012 99356
rect 224880 72486 224908 99350
rect 225800 95946 225828 102068
rect 226628 99414 226656 102068
rect 226248 99408 226300 99414
rect 226248 99350 226300 99356
rect 226616 99408 226668 99414
rect 226616 99350 226668 99356
rect 225788 95940 225840 95946
rect 225788 95882 225840 95888
rect 224960 91860 225012 91866
rect 224960 91802 225012 91808
rect 224868 72480 224920 72486
rect 224868 72422 224920 72428
rect 224224 24200 224276 24206
rect 224224 24142 224276 24148
rect 224972 3482 225000 91802
rect 226260 40866 226288 99350
rect 227456 89758 227484 102068
rect 227628 99408 227680 99414
rect 227628 99350 227680 99356
rect 227444 89752 227496 89758
rect 227444 89694 227496 89700
rect 227444 87032 227496 87038
rect 227444 86974 227496 86980
rect 227456 82074 227484 86974
rect 227076 82068 227128 82074
rect 227076 82010 227128 82016
rect 227444 82068 227496 82074
rect 227444 82010 227496 82016
rect 227088 77353 227116 82010
rect 227074 77344 227130 77353
rect 227074 77279 227130 77288
rect 227258 77344 227314 77353
rect 227314 77302 227392 77330
rect 227258 77279 227314 77288
rect 227364 70514 227392 77302
rect 227352 70508 227404 70514
rect 227352 70450 227404 70456
rect 227260 70372 227312 70378
rect 227260 70314 227312 70320
rect 227272 67833 227300 70314
rect 227258 67824 227314 67833
rect 227258 67759 227314 67768
rect 227258 67688 227314 67697
rect 227258 67623 227314 67632
rect 227272 66230 227300 67623
rect 227260 66224 227312 66230
rect 227260 66166 227312 66172
rect 227444 66224 227496 66230
rect 227444 66166 227496 66172
rect 227456 61441 227484 66166
rect 227442 61432 227498 61441
rect 227442 61367 227498 61376
rect 227350 48376 227406 48385
rect 227272 48334 227350 48362
rect 227272 41478 227300 48334
rect 227350 48311 227406 48320
rect 227260 41472 227312 41478
rect 227260 41414 227312 41420
rect 227352 41336 227404 41342
rect 227352 41278 227404 41284
rect 226248 40860 226300 40866
rect 226248 40802 226300 40808
rect 227364 37262 227392 41278
rect 227352 37256 227404 37262
rect 227352 37198 227404 37204
rect 227444 27668 227496 27674
rect 227444 27610 227496 27616
rect 227456 25566 227484 27610
rect 226340 25560 226392 25566
rect 226340 25502 226392 25508
rect 227444 25560 227496 25566
rect 227444 25502 227496 25508
rect 226352 3482 226380 25502
rect 227640 22778 227668 99350
rect 228284 98802 228312 102068
rect 229112 99414 229140 102068
rect 229954 102054 230428 102082
rect 229100 99408 229152 99414
rect 229100 99350 229152 99356
rect 230296 99408 230348 99414
rect 230296 99350 230348 99356
rect 228272 98796 228324 98802
rect 228272 98738 228324 98744
rect 227720 90432 227772 90438
rect 227720 90374 227772 90380
rect 227628 22772 227680 22778
rect 227628 22714 227680 22720
rect 227732 3602 227760 90374
rect 230308 55894 230336 99350
rect 227812 55888 227864 55894
rect 227812 55830 227864 55836
rect 230296 55888 230348 55894
rect 230296 55830 230348 55836
rect 227720 3596 227772 3602
rect 227720 3538 227772 3544
rect 227824 3482 227852 55830
rect 230400 26926 230428 102054
rect 230768 97306 230796 102068
rect 231610 102054 231808 102082
rect 231124 100088 231176 100094
rect 231124 100030 231176 100036
rect 230756 97300 230808 97306
rect 230756 97242 230808 97248
rect 231136 57254 231164 100030
rect 230480 57248 230532 57254
rect 230480 57190 230532 57196
rect 231124 57248 231176 57254
rect 231124 57190 231176 57196
rect 229100 26920 229152 26926
rect 229100 26862 229152 26868
rect 230388 26920 230440 26926
rect 230388 26862 230440 26868
rect 228916 3596 228968 3602
rect 228916 3538 228968 3544
rect 219452 3454 220584 3482
rect 220832 3454 221780 3482
rect 222212 3454 222976 3482
rect 223592 3454 224172 3482
rect 224972 3454 225368 3482
rect 226352 3454 226564 3482
rect 220556 480 220584 3454
rect 221752 480 221780 3454
rect 222948 480 222976 3454
rect 224144 480 224172 3454
rect 225340 480 225368 3454
rect 226536 480 226564 3454
rect 227732 3454 227852 3482
rect 227732 480 227760 3454
rect 228928 480 228956 3538
rect 229112 3482 229140 26862
rect 230492 3482 230520 57190
rect 231780 50454 231808 102054
rect 232424 99414 232452 102068
rect 233252 99414 233280 102068
rect 234094 102054 234568 102082
rect 232412 99408 232464 99414
rect 232412 99350 232464 99356
rect 233148 99408 233200 99414
rect 233148 99350 233200 99356
rect 233240 99408 233292 99414
rect 233240 99350 233292 99356
rect 234436 99408 234488 99414
rect 234436 99350 234488 99356
rect 231860 89072 231912 89078
rect 231860 89014 231912 89020
rect 231768 50448 231820 50454
rect 231768 50390 231820 50396
rect 231872 3482 231900 89014
rect 233160 6186 233188 99350
rect 234448 58818 234476 99350
rect 234436 58812 234488 58818
rect 234436 58754 234488 58760
rect 233240 28280 233292 28286
rect 233240 28222 233292 28228
rect 233148 6180 233200 6186
rect 233148 6122 233200 6128
rect 233252 3482 233280 28222
rect 234540 24138 234568 102054
rect 234908 100706 234936 102068
rect 235750 102054 235948 102082
rect 236578 102054 237328 102082
rect 234896 100700 234948 100706
rect 234896 100642 234948 100648
rect 235920 60110 235948 102054
rect 236644 100700 236696 100706
rect 236644 100642 236696 100648
rect 235908 60104 235960 60110
rect 235908 60046 235960 60052
rect 234620 58676 234672 58682
rect 234620 58618 234672 58624
rect 234528 24132 234580 24138
rect 234528 24074 234580 24080
rect 234632 3482 234660 58618
rect 236000 42084 236052 42090
rect 236000 42026 236052 42032
rect 229112 3454 230152 3482
rect 230492 3454 231348 3482
rect 231872 3454 232544 3482
rect 233252 3454 233740 3482
rect 234632 3454 234844 3482
rect 230124 480 230152 3454
rect 231320 480 231348 3454
rect 232516 480 232544 3454
rect 233712 480 233740 3454
rect 234816 480 234844 3454
rect 236012 480 236040 42026
rect 236656 28286 236684 100642
rect 237300 37942 237328 102054
rect 237392 100706 237420 102068
rect 237380 100700 237432 100706
rect 237380 100642 237432 100648
rect 238220 100094 238248 102068
rect 238668 100700 238720 100706
rect 238668 100642 238720 100648
rect 238208 100088 238260 100094
rect 238208 100030 238260 100036
rect 237380 60036 237432 60042
rect 237380 59978 237432 59984
rect 237288 37936 237340 37942
rect 237288 37878 237340 37884
rect 236644 28280 236696 28286
rect 236644 28222 236696 28228
rect 237196 6248 237248 6254
rect 237196 6190 237248 6196
rect 237208 480 237236 6190
rect 237392 3482 237420 59978
rect 238680 42090 238708 100642
rect 239048 99754 239076 102068
rect 239784 102054 239890 102082
rect 239036 99748 239088 99754
rect 239036 99690 239088 99696
rect 239784 96665 239812 102054
rect 240704 100162 240732 102068
rect 240692 100156 240744 100162
rect 240692 100098 240744 100104
rect 241428 100156 241480 100162
rect 241428 100098 241480 100104
rect 240048 99748 240100 99754
rect 240048 99690 240100 99696
rect 239770 96656 239826 96665
rect 239770 96591 239826 96600
rect 239954 96656 240010 96665
rect 239954 96591 240010 96600
rect 239968 87038 239996 96591
rect 239864 87032 239916 87038
rect 239864 86974 239916 86980
rect 239956 87032 240008 87038
rect 239956 86974 240008 86980
rect 239876 81870 239904 86974
rect 239864 81864 239916 81870
rect 239864 81806 239916 81812
rect 239864 77376 239916 77382
rect 239784 77324 239864 77330
rect 239784 77318 239916 77324
rect 239784 77302 239904 77318
rect 239784 77246 239812 77302
rect 239772 77240 239824 77246
rect 239772 77182 239824 77188
rect 239864 67652 239916 67658
rect 239864 67594 239916 67600
rect 239876 62966 239904 67594
rect 239864 62960 239916 62966
rect 239864 62902 239916 62908
rect 239680 57996 239732 58002
rect 239680 57938 239732 57944
rect 239692 51134 239720 57938
rect 239680 51128 239732 51134
rect 239680 51070 239732 51076
rect 239680 48340 239732 48346
rect 239680 48282 239732 48288
rect 239692 43450 239720 48282
rect 239680 43444 239732 43450
rect 239680 43386 239732 43392
rect 238668 42084 238720 42090
rect 238668 42026 238720 42032
rect 238760 38072 238812 38078
rect 238760 38014 238812 38020
rect 238772 3482 238800 38014
rect 240060 7614 240088 99690
rect 240140 97368 240192 97374
rect 240140 97310 240192 97316
rect 240048 7608 240100 7614
rect 240048 7550 240100 7556
rect 240152 3482 240180 97310
rect 241440 11830 241468 100098
rect 241532 99482 241560 102068
rect 242282 102054 242848 102082
rect 241520 99476 241572 99482
rect 241520 99418 241572 99424
rect 242820 44878 242848 102054
rect 243096 100706 243124 102068
rect 243938 102054 244228 102082
rect 243084 100700 243136 100706
rect 243084 100642 243136 100648
rect 244096 100700 244148 100706
rect 244096 100642 244148 100648
rect 244108 73846 244136 100642
rect 244096 73840 244148 73846
rect 244096 73782 244148 73788
rect 242900 46232 242952 46238
rect 242900 46174 242952 46180
rect 241520 44872 241572 44878
rect 241520 44814 241572 44820
rect 242808 44872 242860 44878
rect 242808 44814 242860 44820
rect 241428 11824 241480 11830
rect 241428 11766 241480 11772
rect 241532 3482 241560 44814
rect 242912 3482 242940 46174
rect 244200 8974 244228 102054
rect 244752 99414 244780 102068
rect 245488 102054 245594 102082
rect 246422 102054 246988 102082
rect 244740 99408 244792 99414
rect 244740 99350 244792 99356
rect 245488 75206 245516 102054
rect 246304 100156 246356 100162
rect 246304 100098 246356 100104
rect 245568 99408 245620 99414
rect 245568 99350 245620 99356
rect 245476 75200 245528 75206
rect 245476 75142 245528 75148
rect 244280 61464 244332 61470
rect 244280 61406 244332 61412
rect 244188 8968 244240 8974
rect 244188 8910 244240 8916
rect 244292 3534 244320 61406
rect 245580 46238 245608 99350
rect 245568 46232 245620 46238
rect 245568 46174 245620 46180
rect 245660 43512 245712 43518
rect 245660 43454 245712 43460
rect 244372 7744 244424 7750
rect 244372 7686 244424 7692
rect 244280 3528 244332 3534
rect 237392 3454 238432 3482
rect 238772 3454 239628 3482
rect 240152 3454 240824 3482
rect 241532 3454 242020 3482
rect 242912 3454 243216 3482
rect 244280 3470 244332 3476
rect 238404 480 238432 3454
rect 239600 480 239628 3454
rect 240796 480 240824 3454
rect 241992 480 242020 3454
rect 243188 480 243216 3454
rect 244384 480 244412 7686
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245672 3482 245700 43454
rect 246316 10334 246344 100098
rect 246960 51746 246988 102054
rect 247236 99414 247264 102068
rect 248078 102054 248368 102082
rect 248906 102054 249656 102082
rect 247224 99408 247276 99414
rect 247224 99350 247276 99356
rect 248236 99408 248288 99414
rect 248236 99350 248288 99356
rect 246948 51740 247000 51746
rect 246948 51682 247000 51688
rect 248248 29714 248276 99350
rect 248236 29708 248288 29714
rect 248236 29650 248288 29656
rect 247040 29640 247092 29646
rect 247040 29582 247092 29588
rect 246304 10328 246356 10334
rect 246304 10270 246356 10276
rect 247052 3482 247080 29582
rect 248340 13122 248368 102054
rect 248420 62824 248472 62830
rect 248420 62766 248472 62772
rect 248328 13116 248380 13122
rect 248328 13058 248380 13064
rect 248432 3482 248460 62766
rect 249628 53106 249656 102054
rect 249616 53100 249668 53106
rect 249616 53042 249668 53048
rect 249720 47598 249748 102068
rect 250562 102054 251128 102082
rect 250444 99476 250496 99482
rect 250444 99418 250496 99424
rect 250456 62830 250484 99418
rect 250444 62824 250496 62830
rect 250444 62766 250496 62772
rect 249800 47660 249852 47666
rect 249800 47602 249852 47608
rect 249708 47592 249760 47598
rect 249708 47534 249760 47540
rect 249812 3482 249840 47602
rect 251100 14482 251128 102054
rect 251376 99414 251404 102068
rect 252218 102054 252416 102082
rect 251364 99408 251416 99414
rect 251364 99350 251416 99356
rect 252388 49026 252416 102054
rect 253032 99414 253060 102068
rect 252468 99408 252520 99414
rect 252468 99350 252520 99356
rect 253020 99408 253072 99414
rect 253020 99350 253072 99356
rect 252376 49020 252428 49026
rect 252376 48962 252428 48968
rect 252480 35222 252508 99350
rect 253860 64190 253888 102068
rect 254702 102054 255268 102082
rect 254584 99408 254636 99414
rect 254584 99350 254636 99356
rect 254596 76634 254624 99350
rect 254584 76628 254636 76634
rect 254584 76570 254636 76576
rect 252560 64184 252612 64190
rect 252560 64126 252612 64132
rect 253848 64184 253900 64190
rect 253848 64126 253900 64132
rect 252468 35216 252520 35222
rect 252468 35158 252520 35164
rect 251088 14476 251140 14482
rect 251088 14418 251140 14424
rect 251456 9104 251508 9110
rect 251456 9046 251508 9052
rect 245580 480 245608 3470
rect 245672 3454 246804 3482
rect 247052 3454 248000 3482
rect 248432 3454 249196 3482
rect 249812 3454 250392 3482
rect 246776 480 246804 3454
rect 247972 480 248000 3454
rect 249168 480 249196 3454
rect 250364 480 250392 3454
rect 251468 480 251496 9046
rect 252572 3482 252600 64126
rect 255240 31074 255268 102054
rect 255516 100162 255544 102068
rect 256358 102054 256648 102082
rect 257186 102054 257936 102082
rect 255504 100156 255556 100162
rect 255504 100098 255556 100104
rect 256620 69698 256648 102054
rect 257908 82142 257936 102054
rect 256700 82136 256752 82142
rect 256700 82078 256752 82084
rect 257896 82136 257948 82142
rect 257896 82078 257948 82084
rect 256608 69692 256660 69698
rect 256608 69634 256660 69640
rect 255320 65612 255372 65618
rect 255320 65554 255372 65560
rect 253940 31068 253992 31074
rect 253940 31010 253992 31016
rect 255228 31068 255280 31074
rect 255228 31010 255280 31016
rect 253848 4888 253900 4894
rect 253848 4830 253900 4836
rect 252572 3454 252692 3482
rect 252664 480 252692 3454
rect 253860 480 253888 4830
rect 253952 3482 253980 31010
rect 255332 3482 255360 65554
rect 256712 3482 256740 82078
rect 258000 17406 258028 102068
rect 258842 102054 259408 102082
rect 258080 32428 258132 32434
rect 258080 32370 258132 32376
rect 257988 17400 258040 17406
rect 257988 17342 258040 17348
rect 258092 3482 258120 32370
rect 259380 11762 259408 102054
rect 259656 99414 259684 102068
rect 260498 102054 260696 102082
rect 259644 99408 259696 99414
rect 259644 99350 259696 99356
rect 260668 77994 260696 102054
rect 261312 100094 261340 102068
rect 262140 100230 262168 102068
rect 262982 102054 263548 102082
rect 262128 100224 262180 100230
rect 262128 100166 262180 100172
rect 261484 100156 261536 100162
rect 261484 100098 261536 100104
rect 261300 100088 261352 100094
rect 261300 100030 261352 100036
rect 260748 99408 260800 99414
rect 260748 99350 260800 99356
rect 260656 77988 260708 77994
rect 260656 77930 260708 77936
rect 259460 66972 259512 66978
rect 259460 66914 259512 66920
rect 259368 11756 259420 11762
rect 259368 11698 259420 11704
rect 259472 3482 259500 66914
rect 260760 32434 260788 99350
rect 260840 50380 260892 50386
rect 260840 50322 260892 50328
rect 260748 32428 260800 32434
rect 260748 32370 260800 32376
rect 260852 3482 260880 50322
rect 261496 15910 261524 100098
rect 263520 79354 263548 102054
rect 263796 100706 263824 102068
rect 264546 102054 264928 102082
rect 263784 100700 263836 100706
rect 263784 100642 263836 100648
rect 264796 100700 264848 100706
rect 264796 100642 264848 100648
rect 264808 87718 264836 100642
rect 264796 87712 264848 87718
rect 264796 87654 264848 87660
rect 263508 79348 263560 79354
rect 263508 79290 263560 79296
rect 262220 68400 262272 68406
rect 262220 68342 262272 68348
rect 261484 15904 261536 15910
rect 261484 15846 261536 15852
rect 262232 3602 262260 68342
rect 263600 51808 263652 51814
rect 263600 51750 263652 51756
rect 262312 33788 262364 33794
rect 262312 33730 262364 33736
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 262324 3482 262352 33730
rect 263612 12442 263640 51750
rect 264900 33794 264928 102054
rect 265360 100434 265388 102068
rect 266188 100722 266216 102068
rect 267030 102054 267688 102082
rect 266188 100694 266308 100722
rect 265348 100428 265400 100434
rect 265348 100370 265400 100376
rect 266176 100428 266228 100434
rect 266176 100370 266228 100376
rect 266188 80850 266216 100370
rect 266176 80844 266228 80850
rect 266176 80786 266228 80792
rect 264888 33788 264940 33794
rect 264888 33730 264940 33736
rect 263600 12436 263652 12442
rect 263600 12378 263652 12384
rect 264612 12436 264664 12442
rect 264612 12378 264664 12384
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 253952 3454 255084 3482
rect 255332 3454 256280 3482
rect 256712 3454 257476 3482
rect 258092 3454 258672 3482
rect 259472 3454 259868 3482
rect 260852 3454 261064 3482
rect 255056 480 255084 3454
rect 256252 480 256280 3454
rect 257448 480 257476 3454
rect 258644 480 258672 3454
rect 259840 480 259868 3454
rect 261036 480 261064 3454
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3538
rect 264624 480 264652 12378
rect 266280 10470 266308 100694
rect 267004 100020 267056 100026
rect 267004 99962 267056 99968
rect 267016 96626 267044 99962
rect 267004 96620 267056 96626
rect 267004 96562 267056 96568
rect 267004 89684 267056 89690
rect 267004 89626 267056 89632
rect 267016 86986 267044 89626
rect 267016 86958 267136 86986
rect 267108 80170 267136 86958
rect 267096 80164 267148 80170
rect 267096 80106 267148 80112
rect 267096 77308 267148 77314
rect 267096 77250 267148 77256
rect 267108 70446 267136 77250
rect 267096 70440 267148 70446
rect 267096 70382 267148 70388
rect 266360 69828 266412 69834
rect 266360 69770 266412 69776
rect 266372 12442 266400 69770
rect 267096 67652 267148 67658
rect 267096 67594 267148 67600
rect 267108 62762 267136 67594
rect 267096 62756 267148 62762
rect 267096 62698 267148 62704
rect 267096 57996 267148 58002
rect 267096 57938 267148 57944
rect 267108 51134 267136 57938
rect 267096 51128 267148 51134
rect 267096 51070 267148 51076
rect 267660 50386 267688 102054
rect 267844 100706 267872 102068
rect 268686 102054 268976 102082
rect 267832 100700 267884 100706
rect 267832 100642 267884 100648
rect 268948 65686 268976 102054
rect 269028 100700 269080 100706
rect 269028 100642 269080 100648
rect 268936 65680 268988 65686
rect 268936 65622 268988 65628
rect 267648 50380 267700 50386
rect 267648 50322 267700 50328
rect 267096 48340 267148 48346
rect 267096 48282 267148 48288
rect 267108 41546 267136 48282
rect 267740 46980 267792 46986
rect 267740 46922 267792 46928
rect 267096 41540 267148 41546
rect 267096 41482 267148 41488
rect 267004 38684 267056 38690
rect 267004 38626 267056 38632
rect 267016 31754 267044 38626
rect 267004 31748 267056 31754
rect 267004 31690 267056 31696
rect 267188 31748 267240 31754
rect 267188 31690 267240 31696
rect 267200 28966 267228 31690
rect 267188 28960 267240 28966
rect 267188 28902 267240 28908
rect 267752 22710 267780 46922
rect 267740 22704 267792 22710
rect 267740 22646 267792 22652
rect 267096 19372 267148 19378
rect 267096 19314 267148 19320
rect 267108 12458 267136 19314
rect 269040 18698 269068 100642
rect 269500 99958 269528 102068
rect 270328 100722 270356 102068
rect 270328 100694 270448 100722
rect 269488 99952 269540 99958
rect 269488 99894 269540 99900
rect 270316 99952 270368 99958
rect 270316 99894 270368 99900
rect 270328 51814 270356 99894
rect 270316 51808 270368 51814
rect 270316 51750 270368 51756
rect 270420 40798 270448 100694
rect 271156 100026 271184 102068
rect 271984 100706 272012 102068
rect 272826 102054 273116 102082
rect 271972 100700 272024 100706
rect 271972 100642 272024 100648
rect 271144 100020 271196 100026
rect 271144 99962 271196 99968
rect 272524 100020 272576 100026
rect 272524 99962 272576 99968
rect 270500 71120 270552 71126
rect 270500 71062 270552 71068
rect 270408 40792 270460 40798
rect 270408 40734 270460 40740
rect 269028 18692 269080 18698
rect 269028 18634 269080 18640
rect 266360 12436 266412 12442
rect 266360 12378 266412 12384
rect 267004 12436 267056 12442
rect 267108 12430 267228 12458
rect 267004 12378 267056 12384
rect 266268 10464 266320 10470
rect 266268 10406 266320 10412
rect 265808 4820 265860 4826
rect 265808 4762 265860 4768
rect 265820 480 265848 4762
rect 267016 480 267044 12378
rect 267200 4826 267228 12430
rect 269304 10396 269356 10402
rect 269304 10338 269356 10344
rect 268108 9716 268160 9722
rect 268108 9658 268160 9664
rect 267188 4820 267240 4826
rect 267188 4762 267240 4768
rect 268120 480 268148 9658
rect 269316 480 269344 10338
rect 270512 480 270540 71062
rect 270592 39432 270644 39438
rect 270592 39374 270644 39380
rect 270604 12442 270632 39374
rect 272536 17338 272564 99962
rect 273088 83570 273116 102054
rect 273168 100700 273220 100706
rect 273168 100642 273220 100648
rect 273076 83564 273128 83570
rect 273076 83506 273128 83512
rect 273180 53174 273208 100642
rect 273640 100026 273668 102068
rect 274376 102054 274482 102082
rect 275310 102054 275968 102082
rect 273628 100020 273680 100026
rect 273628 99962 273680 99968
rect 274376 96665 274404 102054
rect 274362 96656 274418 96665
rect 274362 96591 274418 96600
rect 274546 96656 274602 96665
rect 274546 96591 274602 96600
rect 274560 89758 274588 96591
rect 274364 89752 274416 89758
rect 274548 89752 274600 89758
rect 274416 89700 274496 89706
rect 274364 89694 274496 89700
rect 274548 89694 274600 89700
rect 274376 89678 274496 89694
rect 274468 89570 274496 89678
rect 274468 89542 274588 89570
rect 273260 72548 273312 72554
rect 273260 72490 273312 72496
rect 273168 53168 273220 53174
rect 273168 53110 273220 53116
rect 272524 17332 272576 17338
rect 272524 17274 272576 17280
rect 270592 12436 270644 12442
rect 270592 12378 270644 12384
rect 271696 12436 271748 12442
rect 271696 12378 271748 12384
rect 271708 480 271736 12378
rect 272892 11892 272944 11898
rect 272892 11834 272944 11840
rect 272904 480 272932 11834
rect 273272 3482 273300 72490
rect 274560 71194 274588 89542
rect 274640 87644 274692 87650
rect 274640 87586 274692 87592
rect 274548 71188 274600 71194
rect 274548 71130 274600 71136
rect 274548 67652 274600 67658
rect 274548 67594 274600 67600
rect 274560 67522 274588 67594
rect 274364 67516 274416 67522
rect 274364 67458 274416 67464
rect 274548 67516 274600 67522
rect 274548 67458 274600 67464
rect 274376 54670 274404 67458
rect 274364 54664 274416 54670
rect 274364 54606 274416 54612
rect 274652 3482 274680 87586
rect 275940 84998 275968 102054
rect 276124 100706 276152 102068
rect 276966 102054 277256 102082
rect 276112 100700 276164 100706
rect 276112 100642 276164 100648
rect 277228 87650 277256 102054
rect 277308 100700 277360 100706
rect 277308 100642 277360 100648
rect 277216 87644 277268 87650
rect 277216 87586 277268 87592
rect 275928 84992 275980 84998
rect 275928 84934 275980 84940
rect 277320 80782 277348 100642
rect 277780 94654 277808 102068
rect 278516 102054 278622 102082
rect 279450 102054 280108 102082
rect 278516 96762 278544 102054
rect 278504 96756 278556 96762
rect 278504 96698 278556 96704
rect 278688 96756 278740 96762
rect 278688 96698 278740 96704
rect 278700 96626 278728 96698
rect 278688 96620 278740 96626
rect 278688 96562 278740 96568
rect 277768 94648 277820 94654
rect 277768 94590 277820 94596
rect 278596 87032 278648 87038
rect 278596 86974 278648 86980
rect 277308 80776 277360 80782
rect 277308 80718 277360 80724
rect 278608 80102 278636 86974
rect 278596 80096 278648 80102
rect 278596 80038 278648 80044
rect 278688 79960 278740 79966
rect 278688 79902 278740 79908
rect 277400 73908 277452 73914
rect 277400 73850 277452 73856
rect 276020 13184 276072 13190
rect 276020 13126 276072 13132
rect 276032 3482 276060 13126
rect 277412 3482 277440 73850
rect 278700 70530 278728 79902
rect 278608 70502 278728 70530
rect 278608 67046 278636 70502
rect 278596 67040 278648 67046
rect 278596 66982 278648 66988
rect 278780 55956 278832 55962
rect 278780 55898 278832 55904
rect 278792 3482 278820 55898
rect 280080 35290 280108 102054
rect 280264 100162 280292 102068
rect 281106 102054 281488 102082
rect 280252 100156 280304 100162
rect 280252 100098 280304 100104
rect 281356 100156 281408 100162
rect 281356 100098 281408 100104
rect 281368 86358 281396 100098
rect 281356 86352 281408 86358
rect 281356 86294 281408 86300
rect 280160 75268 280212 75274
rect 280160 75210 280212 75216
rect 278872 35284 278924 35290
rect 278872 35226 278924 35232
rect 280068 35284 280120 35290
rect 280068 35226 280120 35232
rect 278884 3602 278912 35226
rect 278872 3596 278924 3602
rect 278872 3538 278924 3544
rect 280068 3596 280120 3602
rect 280068 3538 280120 3544
rect 273272 3454 274128 3482
rect 274652 3454 275324 3482
rect 276032 3454 276520 3482
rect 277412 3454 277716 3482
rect 278792 3454 278912 3482
rect 274100 480 274128 3454
rect 275296 480 275324 3454
rect 276492 480 276520 3454
rect 277688 480 277716 3454
rect 278884 480 278912 3454
rect 280080 480 280108 3538
rect 280172 3482 280200 75210
rect 281460 54602 281488 102054
rect 281920 99754 281948 102068
rect 281908 99748 281960 99754
rect 281908 99690 281960 99696
rect 282748 89146 282776 102068
rect 283590 102054 284248 102082
rect 283564 100020 283616 100026
rect 283564 99962 283616 99968
rect 282828 99748 282880 99754
rect 282828 99690 282880 99696
rect 282736 89140 282788 89146
rect 282736 89082 282788 89088
rect 282840 72554 282868 99690
rect 282828 72548 282880 72554
rect 282828 72490 282880 72496
rect 281540 57316 281592 57322
rect 281540 57258 281592 57264
rect 281448 54596 281500 54602
rect 281448 54538 281500 54544
rect 281552 3482 281580 57258
rect 283576 18766 283604 99962
rect 284220 40730 284248 102054
rect 284404 99414 284432 102068
rect 285246 102054 285536 102082
rect 284392 99408 284444 99414
rect 284392 99350 284444 99356
rect 285508 90438 285536 102054
rect 286060 99414 286088 102068
rect 286888 99498 286916 102068
rect 286888 99470 287008 99498
rect 285588 99408 285640 99414
rect 285588 99350 285640 99356
rect 286048 99408 286100 99414
rect 286048 99350 286100 99356
rect 286876 99408 286928 99414
rect 286876 99350 286928 99356
rect 285496 90432 285548 90438
rect 285496 90374 285548 90380
rect 284300 76560 284352 76566
rect 284300 76502 284352 76508
rect 284208 40724 284260 40730
rect 284208 40666 284260 40672
rect 283564 18760 283616 18766
rect 283564 18702 283616 18708
rect 282920 14544 282972 14550
rect 282920 14486 282972 14492
rect 282932 3482 282960 14486
rect 284312 3482 284340 76502
rect 285600 71194 285628 99350
rect 285588 71188 285640 71194
rect 285588 71130 285640 71136
rect 286888 57390 286916 99350
rect 286876 57384 286928 57390
rect 286876 57326 286928 57332
rect 286980 56030 287008 99470
rect 287624 99414 287652 102068
rect 288452 99414 288480 102068
rect 289280 100162 289308 102068
rect 289268 100156 289320 100162
rect 289268 100098 289320 100104
rect 290108 99414 290136 102068
rect 290950 102054 291148 102082
rect 291778 102054 292528 102082
rect 287612 99408 287664 99414
rect 287612 99350 287664 99356
rect 288348 99408 288400 99414
rect 288348 99350 288400 99356
rect 288440 99408 288492 99414
rect 288440 99350 288492 99356
rect 289728 99408 289780 99414
rect 289728 99350 289780 99356
rect 290096 99408 290148 99414
rect 290096 99350 290148 99356
rect 291016 99408 291068 99414
rect 291016 99350 291068 99356
rect 287060 94512 287112 94518
rect 287060 94454 287112 94460
rect 286968 56024 287020 56030
rect 286968 55966 287020 55972
rect 285680 54528 285732 54534
rect 285680 54470 285732 54476
rect 285692 3482 285720 54470
rect 280172 3454 281304 3482
rect 281552 3454 282500 3482
rect 282932 3454 283696 3482
rect 284312 3454 284800 3482
rect 285692 3454 285996 3482
rect 281276 480 281304 3454
rect 282472 480 282500 3454
rect 283668 480 283696 3454
rect 284772 480 284800 3454
rect 285968 480 285996 3454
rect 287072 1426 287100 94454
rect 288360 29646 288388 99350
rect 289740 84930 289768 99350
rect 291028 91866 291056 99350
rect 291016 91860 291068 91866
rect 291016 91802 291068 91808
rect 289728 84924 289780 84930
rect 289728 84866 289780 84872
rect 288440 49088 288492 49094
rect 288440 49030 288492 49036
rect 288348 29640 288400 29646
rect 288348 29582 288400 29588
rect 287152 15972 287204 15978
rect 287152 15914 287204 15920
rect 287060 1420 287112 1426
rect 287060 1362 287112 1368
rect 287164 480 287192 15914
rect 288452 3482 288480 49030
rect 291120 15978 291148 102054
rect 291844 100224 291896 100230
rect 291844 100166 291896 100172
rect 291200 78056 291252 78062
rect 291200 77998 291252 78004
rect 291108 15972 291160 15978
rect 291108 15914 291160 15920
rect 290740 4820 290792 4826
rect 290740 4762 290792 4768
rect 288452 3454 289584 3482
rect 288348 1420 288400 1426
rect 288348 1362 288400 1368
rect 288360 480 288388 1362
rect 289556 480 289584 3454
rect 290752 480 290780 4762
rect 291212 3618 291240 77998
rect 291856 4894 291884 100166
rect 292500 68474 292528 102054
rect 292592 100026 292620 102068
rect 293420 100230 293448 102068
rect 293408 100224 293460 100230
rect 293408 100166 293460 100172
rect 292580 100020 292632 100026
rect 292580 99962 292632 99968
rect 294248 99414 294276 102068
rect 294604 100088 294656 100094
rect 294604 100030 294656 100036
rect 294236 99408 294288 99414
rect 294236 99350 294288 99356
rect 292488 68468 292540 68474
rect 292488 68410 292540 68416
rect 292580 61396 292632 61402
rect 292580 61338 292632 61344
rect 291844 4888 291896 4894
rect 291844 4830 291896 4836
rect 291212 3590 291976 3618
rect 291948 480 291976 3590
rect 292592 3482 292620 61338
rect 293960 17264 294012 17270
rect 293960 17206 294012 17212
rect 293972 3482 294000 17206
rect 294616 13190 294644 100030
rect 295076 93226 295104 102068
rect 295904 99414 295932 102068
rect 296732 99414 296760 102068
rect 297574 102054 298048 102082
rect 295248 99408 295300 99414
rect 295248 99350 295300 99356
rect 295892 99408 295944 99414
rect 295892 99350 295944 99356
rect 296628 99408 296680 99414
rect 296628 99350 296680 99356
rect 296720 99408 296772 99414
rect 296720 99350 296772 99356
rect 297916 99408 297968 99414
rect 297916 99350 297968 99356
rect 295064 93220 295116 93226
rect 295064 93162 295116 93168
rect 295260 66978 295288 99350
rect 295340 79416 295392 79422
rect 295340 79358 295392 79364
rect 295248 66972 295300 66978
rect 295248 66914 295300 66920
rect 294604 13184 294656 13190
rect 294604 13126 294656 13132
rect 295352 3482 295380 79358
rect 296640 55962 296668 99350
rect 297928 65618 297956 99350
rect 297916 65612 297968 65618
rect 297916 65554 297968 65560
rect 296720 62892 296772 62898
rect 296720 62834 296772 62840
rect 296628 55956 296680 55962
rect 296628 55898 296680 55904
rect 292592 3454 293172 3482
rect 293972 3454 294368 3482
rect 295352 3454 295564 3482
rect 293144 480 293172 3454
rect 294340 480 294368 3454
rect 295536 480 295564 3454
rect 296732 480 296760 62834
rect 296812 18624 296864 18630
rect 296812 18566 296864 18572
rect 296824 3346 296852 18566
rect 298020 4826 298048 102054
rect 298388 99414 298416 102068
rect 299230 102054 299428 102082
rect 300058 102054 300808 102082
rect 298376 99408 298428 99414
rect 298376 99350 298428 99356
rect 299296 99408 299348 99414
rect 299296 99350 299348 99356
rect 299308 89078 299336 99350
rect 299296 89072 299348 89078
rect 299296 89014 299348 89020
rect 298100 80708 298152 80714
rect 298100 80650 298152 80656
rect 298008 4820 298060 4826
rect 298008 4762 298060 4768
rect 298112 3346 298140 80650
rect 299400 57322 299428 102054
rect 300124 100020 300176 100026
rect 300124 99962 300176 99968
rect 300136 73914 300164 99962
rect 300780 75274 300808 102054
rect 300872 99414 300900 102068
rect 301714 102054 302188 102082
rect 300860 99408 300912 99414
rect 300860 99350 300912 99356
rect 302056 99408 302108 99414
rect 302056 99350 302108 99356
rect 300768 75268 300820 75274
rect 300768 75210 300820 75216
rect 300124 73908 300176 73914
rect 300124 73850 300176 73856
rect 302068 68406 302096 99350
rect 302056 68400 302108 68406
rect 302056 68342 302108 68348
rect 302160 64258 302188 102054
rect 302528 99482 302556 102068
rect 303370 102054 303568 102082
rect 302516 99476 302568 99482
rect 302516 99418 302568 99424
rect 302240 83496 302292 83502
rect 302240 83438 302292 83444
rect 299480 64252 299532 64258
rect 299480 64194 299532 64200
rect 302148 64252 302200 64258
rect 302148 64194 302200 64200
rect 299388 57316 299440 57322
rect 299388 57258 299440 57264
rect 299492 3346 299520 64194
rect 300860 19984 300912 19990
rect 300860 19926 300912 19932
rect 300872 3346 300900 19926
rect 302252 3346 302280 83438
rect 303540 71126 303568 102054
rect 304184 99414 304212 102068
rect 304264 99476 304316 99482
rect 304264 99418 304316 99424
rect 304172 99408 304224 99414
rect 304172 99350 304224 99356
rect 304276 76566 304304 99418
rect 304908 99408 304960 99414
rect 304908 99350 304960 99356
rect 304264 76560 304316 76566
rect 304264 76502 304316 76508
rect 303528 71120 303580 71126
rect 303528 71062 303580 71068
rect 303620 65544 303672 65550
rect 303620 65486 303672 65492
rect 303632 3346 303660 65486
rect 304920 20058 304948 99350
rect 305012 96014 305040 102068
rect 305854 102054 306328 102082
rect 305000 96008 305052 96014
rect 305000 95950 305052 95956
rect 305000 84856 305052 84862
rect 305000 84798 305052 84804
rect 304908 20052 304960 20058
rect 304908 19994 304960 20000
rect 305012 3602 305040 84798
rect 305092 21480 305144 21486
rect 305092 21422 305144 21428
rect 305000 3596 305052 3602
rect 305000 3538 305052 3544
rect 305104 3482 305132 21422
rect 306300 4146 306328 102054
rect 306668 99550 306696 102068
rect 307510 102054 307708 102082
rect 308338 102054 309088 102082
rect 306656 99544 306708 99550
rect 306656 99486 306708 99492
rect 307680 78062 307708 102054
rect 307760 89004 307812 89010
rect 307760 88946 307812 88952
rect 307668 78056 307720 78062
rect 307668 77998 307720 78004
rect 306380 69760 306432 69766
rect 306380 69702 306432 69708
rect 306288 4140 306340 4146
rect 306288 4082 306340 4088
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 305012 3454 305132 3482
rect 296824 3318 297956 3346
rect 298112 3318 299152 3346
rect 299492 3318 300348 3346
rect 300872 3318 301452 3346
rect 302252 3318 302648 3346
rect 303632 3318 303844 3346
rect 297928 480 297956 3318
rect 299124 480 299152 3318
rect 300320 480 300348 3318
rect 301424 480 301452 3318
rect 302620 480 302648 3318
rect 303816 480 303844 3318
rect 305012 480 305040 3454
rect 306208 480 306236 3538
rect 306392 610 306420 69702
rect 307772 610 307800 88946
rect 309060 4078 309088 102054
rect 309152 99414 309180 102068
rect 309784 100224 309836 100230
rect 309784 100166 309836 100172
rect 309140 99408 309192 99414
rect 309140 99350 309192 99356
rect 309796 86426 309824 100166
rect 309888 100026 309916 102068
rect 309876 100020 309928 100026
rect 309876 99962 309928 99968
rect 310716 99414 310744 102068
rect 311544 99482 311572 102068
rect 311532 99476 311584 99482
rect 311532 99418 311584 99424
rect 310428 99408 310480 99414
rect 310428 99350 310480 99356
rect 310704 99408 310756 99414
rect 310704 99350 310756 99356
rect 311808 99408 311860 99414
rect 311808 99350 311860 99356
rect 309784 86420 309836 86426
rect 309784 86362 309836 86368
rect 309140 86284 309192 86290
rect 309140 86226 309192 86232
rect 309048 4072 309100 4078
rect 309048 4014 309100 4020
rect 309152 610 309180 86226
rect 310440 61470 310468 99350
rect 310520 66904 310572 66910
rect 310520 66846 310572 66852
rect 310428 61464 310480 61470
rect 310428 61406 310480 61412
rect 310532 610 310560 66846
rect 311820 4010 311848 99350
rect 312372 97374 312400 102068
rect 312360 97368 312412 97374
rect 312360 97310 312412 97316
rect 311900 36576 311952 36582
rect 311900 36518 311952 36524
rect 311808 4004 311860 4010
rect 311808 3946 311860 3952
rect 311912 626 311940 36518
rect 313200 3874 313228 102068
rect 314042 102054 314608 102082
rect 313924 99544 313976 99550
rect 313924 99486 313976 99492
rect 313280 90364 313332 90370
rect 313280 90306 313332 90312
rect 313188 3868 313240 3874
rect 313188 3810 313240 3816
rect 313292 3482 313320 90306
rect 313372 68332 313424 68338
rect 313372 68274 313424 68280
rect 313384 3602 313412 68274
rect 313936 62898 313964 99486
rect 313924 62892 313976 62898
rect 313924 62834 313976 62840
rect 314580 36650 314608 102054
rect 314856 99414 314884 102068
rect 315698 102054 315988 102082
rect 314844 99408 314896 99414
rect 314844 99350 314896 99356
rect 315856 99408 315908 99414
rect 315856 99350 315908 99356
rect 315868 82210 315896 99350
rect 315856 82204 315908 82210
rect 315856 82146 315908 82152
rect 314568 36644 314620 36650
rect 314568 36586 314620 36592
rect 314660 22840 314712 22846
rect 314660 22782 314712 22788
rect 313372 3596 313424 3602
rect 313372 3538 313424 3544
rect 314568 3596 314620 3602
rect 314568 3538 314620 3544
rect 313292 3454 313412 3482
rect 306380 604 306432 610
rect 306380 546 306432 552
rect 307392 604 307444 610
rect 307392 546 307444 552
rect 307760 604 307812 610
rect 307760 546 307812 552
rect 308588 604 308640 610
rect 308588 546 308640 552
rect 309140 604 309192 610
rect 309140 546 309192 552
rect 309784 604 309836 610
rect 309784 546 309836 552
rect 310520 604 310572 610
rect 310520 546 310572 552
rect 310980 604 311032 610
rect 311912 598 312216 626
rect 310980 546 311032 552
rect 307404 480 307432 546
rect 308600 480 308628 546
rect 309796 480 309824 546
rect 310992 480 311020 546
rect 312188 480 312216 598
rect 313384 480 313412 3454
rect 314580 480 314608 3538
rect 314672 610 314700 22782
rect 315960 3942 315988 102054
rect 316512 99414 316540 102068
rect 316500 99408 316552 99414
rect 316500 99350 316552 99356
rect 317236 99408 317288 99414
rect 317236 99350 317288 99356
rect 316040 91792 316092 91798
rect 316040 91734 316092 91740
rect 315948 3936 316000 3942
rect 315948 3878 316000 3884
rect 316052 3346 316080 91734
rect 317248 60042 317276 99350
rect 317340 98734 317368 102068
rect 318182 102054 318748 102082
rect 318064 99476 318116 99482
rect 318064 99418 318116 99424
rect 317328 98728 317380 98734
rect 317328 98670 317380 98676
rect 317236 60036 317288 60042
rect 317236 59978 317288 59984
rect 318076 21486 318104 99418
rect 318064 21480 318116 21486
rect 318064 21422 318116 21428
rect 317420 21412 317472 21418
rect 317420 21354 317472 21360
rect 317432 3346 317460 21354
rect 318720 3806 318748 102054
rect 318996 99414 319024 102068
rect 319838 102054 320128 102082
rect 318984 99408 319036 99414
rect 318984 99350 319036 99356
rect 319996 99408 320048 99414
rect 319996 99350 320048 99356
rect 320008 58750 320036 99350
rect 319996 58744 320048 58750
rect 319996 58686 320048 58692
rect 318800 24200 318852 24206
rect 318800 24142 318852 24148
rect 318708 3800 318760 3806
rect 318708 3742 318760 3748
rect 318812 3346 318840 24142
rect 320100 19990 320128 102054
rect 320652 99414 320680 102068
rect 321388 102054 321494 102082
rect 322322 102054 322888 102082
rect 320640 99408 320692 99414
rect 320640 99350 320692 99356
rect 320180 93152 320232 93158
rect 320180 93094 320232 93100
rect 320088 19984 320140 19990
rect 320088 19926 320140 19932
rect 320192 3346 320220 93094
rect 321388 22846 321416 102054
rect 322204 100156 322256 100162
rect 322204 100098 322256 100104
rect 321468 99408 321520 99414
rect 321468 99350 321520 99356
rect 321376 22840 321428 22846
rect 321376 22782 321428 22788
rect 321480 3738 321508 99350
rect 321560 71052 321612 71058
rect 321560 70994 321612 71000
rect 321468 3732 321520 3738
rect 321468 3674 321520 3680
rect 321572 3482 321600 70994
rect 322216 69766 322244 100098
rect 322204 69760 322256 69766
rect 322204 69702 322256 69708
rect 322860 61402 322888 102054
rect 323136 99414 323164 102068
rect 323978 102054 324176 102082
rect 323124 99408 323176 99414
rect 323124 99350 323176 99356
rect 322848 61396 322900 61402
rect 322848 61338 322900 61344
rect 321652 38004 321704 38010
rect 321652 37946 321704 37952
rect 321664 3602 321692 37946
rect 324148 24206 324176 102054
rect 324792 99414 324820 102068
rect 324228 99408 324280 99414
rect 324228 99350 324280 99356
rect 324780 99408 324832 99414
rect 324780 99350 324832 99356
rect 324136 24200 324188 24206
rect 324136 24142 324188 24148
rect 324044 7676 324096 7682
rect 324044 7618 324096 7624
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 321572 3454 321692 3482
rect 316052 3318 317000 3346
rect 317432 3318 318104 3346
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 314660 604 314712 610
rect 314660 546 314712 552
rect 315764 604 315816 610
rect 315764 546 315816 552
rect 315776 480 315804 546
rect 316972 480 317000 3318
rect 318076 480 318104 3318
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 3454
rect 322860 480 322888 3538
rect 324056 480 324084 7618
rect 324240 3670 324268 99350
rect 324320 57248 324372 57254
rect 324320 57190 324372 57196
rect 324228 3664 324280 3670
rect 324228 3606 324280 3612
rect 324332 3346 324360 57190
rect 325620 3602 325648 102068
rect 326462 102054 327028 102082
rect 326344 99408 326396 99414
rect 326344 99350 326396 99356
rect 325700 39364 325752 39370
rect 325700 39306 325752 39312
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 325712 3482 325740 39306
rect 326356 21418 326384 99350
rect 327000 39438 327028 102054
rect 327276 99414 327304 102068
rect 328118 102054 328408 102082
rect 327264 99408 327316 99414
rect 327264 99350 327316 99356
rect 328276 99408 328328 99414
rect 328276 99350 328328 99356
rect 326988 39432 327040 39438
rect 326988 39374 327040 39380
rect 328288 36582 328316 99350
rect 328276 36576 328328 36582
rect 328276 36518 328328 36524
rect 326344 21412 326396 21418
rect 326344 21354 326396 21360
rect 327632 9036 327684 9042
rect 327632 8978 327684 8984
rect 325712 3454 326476 3482
rect 324332 3318 325280 3346
rect 325252 480 325280 3318
rect 326448 480 326476 3454
rect 327644 480 327672 8978
rect 328380 3534 328408 102054
rect 328932 99414 328960 102068
rect 328920 99408 328972 99414
rect 328920 99350 328972 99356
rect 329760 79422 329788 102068
rect 330602 102054 331168 102082
rect 329748 79416 329800 79422
rect 329748 79358 329800 79364
rect 328460 72480 328512 72486
rect 328460 72422 328512 72428
rect 328368 3528 328420 3534
rect 328368 3470 328420 3476
rect 328472 3482 328500 72422
rect 329840 40860 329892 40866
rect 329840 40802 329892 40808
rect 329852 3482 329880 40802
rect 328472 3454 328868 3482
rect 329852 3454 330064 3482
rect 331140 3466 331168 102054
rect 331416 100094 331444 102068
rect 332258 102054 332548 102082
rect 331404 100088 331456 100094
rect 331404 100030 331456 100036
rect 331864 99408 331916 99414
rect 331864 99350 331916 99356
rect 331220 95940 331272 95946
rect 331220 95882 331272 95888
rect 328840 480 328868 3454
rect 330036 480 330064 3454
rect 331128 3460 331180 3466
rect 331128 3402 331180 3408
rect 331232 480 331260 95882
rect 331876 38010 331904 99350
rect 331864 38004 331916 38010
rect 331864 37946 331916 37952
rect 332520 25634 332548 102054
rect 332980 99414 333008 102068
rect 333716 102054 333822 102082
rect 334650 102054 335308 102082
rect 332968 99408 333020 99414
rect 332968 99350 333020 99356
rect 333716 98666 333744 102054
rect 333796 99408 333848 99414
rect 333796 99350 333848 99356
rect 333704 98660 333756 98666
rect 333704 98602 333756 98608
rect 332508 25628 332560 25634
rect 332508 25570 332560 25576
rect 332600 25560 332652 25566
rect 332600 25502 332652 25508
rect 331312 22772 331364 22778
rect 331312 22714 331364 22720
rect 331324 3482 331352 22714
rect 332612 3482 332640 25502
rect 333808 14550 333836 99350
rect 333980 98796 334032 98802
rect 333980 98738 334032 98744
rect 333796 14544 333848 14550
rect 333796 14486 333848 14492
rect 333992 3482 334020 98738
rect 335280 26994 335308 102054
rect 335464 100162 335492 102068
rect 336306 102054 336688 102082
rect 335452 100156 335504 100162
rect 335452 100098 335504 100104
rect 335360 55888 335412 55894
rect 335360 55830 335412 55836
rect 335268 26988 335320 26994
rect 335268 26930 335320 26936
rect 335372 3482 335400 55830
rect 336660 6254 336688 102054
rect 337120 99414 337148 102068
rect 337948 99498 337976 102068
rect 338790 102054 339448 102082
rect 337948 99470 338068 99498
rect 337108 99408 337160 99414
rect 337108 99350 337160 99356
rect 337936 99408 337988 99414
rect 337936 99350 337988 99356
rect 337948 28354 337976 99350
rect 337936 28348 337988 28354
rect 337936 28290 337988 28296
rect 336740 26920 336792 26926
rect 336740 26862 336792 26868
rect 336648 6248 336700 6254
rect 336648 6190 336700 6196
rect 336752 3482 336780 26862
rect 338040 22778 338068 99470
rect 338120 97300 338172 97306
rect 338120 97242 338172 97248
rect 338028 22772 338080 22778
rect 338028 22714 338080 22720
rect 338132 3482 338160 97242
rect 339420 7682 339448 102054
rect 339604 99414 339632 102068
rect 340446 102054 340736 102082
rect 339592 99408 339644 99414
rect 339592 99350 339644 99356
rect 340708 58682 340736 102054
rect 340788 99408 340840 99414
rect 340788 99350 340840 99356
rect 340696 58676 340748 58682
rect 340696 58618 340748 58624
rect 339500 50448 339552 50454
rect 339500 50390 339552 50396
rect 339408 7676 339460 7682
rect 339408 7618 339460 7624
rect 331324 3454 332456 3482
rect 332612 3454 333652 3482
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 332428 480 332456 3454
rect 333624 480 333652 3454
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339512 480 339540 50390
rect 340800 42158 340828 99350
rect 341260 97306 341288 102068
rect 342088 98598 342116 102068
rect 342930 102054 343588 102082
rect 342076 98592 342128 98598
rect 342076 98534 342128 98540
rect 341248 97300 341300 97306
rect 341248 97242 341300 97248
rect 342076 87032 342128 87038
rect 342076 86974 342128 86980
rect 342088 82074 342116 86974
rect 341708 82068 341760 82074
rect 341708 82010 341760 82016
rect 342076 82068 342128 82074
rect 342076 82010 342128 82016
rect 341720 77353 341748 82010
rect 341706 77344 341762 77353
rect 341706 77279 341762 77288
rect 341890 77344 341946 77353
rect 341946 77302 342024 77330
rect 341890 77279 341946 77288
rect 341996 70514 342024 77302
rect 341984 70508 342036 70514
rect 341984 70450 342036 70456
rect 341892 70372 341944 70378
rect 341892 70314 341944 70320
rect 341904 67833 341932 70314
rect 341890 67824 341946 67833
rect 341890 67759 341946 67768
rect 341890 67688 341946 67697
rect 341890 67623 341946 67632
rect 341904 66230 341932 67623
rect 341892 66224 341944 66230
rect 341892 66166 341944 66172
rect 340880 58812 340932 58818
rect 340880 58754 340932 58760
rect 340788 42152 340840 42158
rect 340788 42094 340840 42100
rect 340696 6180 340748 6186
rect 340696 6122 340748 6128
rect 340708 480 340736 6122
rect 340892 3482 340920 58754
rect 342076 56636 342128 56642
rect 342076 56578 342128 56584
rect 342088 51134 342116 56578
rect 342076 51128 342128 51134
rect 342076 51070 342128 51076
rect 342076 50992 342128 50998
rect 342076 50934 342128 50940
rect 342088 43518 342116 50934
rect 342076 43512 342128 43518
rect 342076 43454 342128 43460
rect 343560 24138 343588 102054
rect 343744 95946 343772 102068
rect 344586 102054 344968 102082
rect 344284 100020 344336 100026
rect 344284 99962 344336 99968
rect 343732 95940 343784 95946
rect 343732 95882 343784 95888
rect 343640 28280 343692 28286
rect 343640 28222 343692 28228
rect 342260 24132 342312 24138
rect 342260 24074 342312 24080
rect 343548 24132 343600 24138
rect 343548 24074 343600 24080
rect 342272 3482 342300 24074
rect 343652 3482 343680 28222
rect 344296 16046 344324 99962
rect 344940 44946 344968 102054
rect 345400 100706 345428 102068
rect 345388 100700 345440 100706
rect 345388 100642 345440 100648
rect 346228 94586 346256 102068
rect 347070 102054 347728 102082
rect 346308 100700 346360 100706
rect 346308 100642 346360 100648
rect 346216 94580 346268 94586
rect 346216 94522 346268 94528
rect 345020 60104 345072 60110
rect 345020 60046 345072 60052
rect 344928 44940 344980 44946
rect 344928 44882 344980 44888
rect 344284 16040 344336 16046
rect 344284 15982 344336 15988
rect 345032 3482 345060 60046
rect 346320 39370 346348 100642
rect 347700 46306 347728 102054
rect 347884 100706 347912 102068
rect 348726 102054 349108 102082
rect 347872 100700 347924 100706
rect 347872 100642 347924 100648
rect 348976 100700 349028 100706
rect 348976 100642 349028 100648
rect 347688 46300 347740 46306
rect 347688 46242 347740 46248
rect 347780 42084 347832 42090
rect 347780 42026 347832 42032
rect 346308 39364 346360 39370
rect 346308 39306 346360 39312
rect 346400 37936 346452 37942
rect 346400 37878 346452 37884
rect 346412 3482 346440 37878
rect 347792 3482 347820 42026
rect 348988 37942 349016 100642
rect 348976 37936 349028 37942
rect 348976 37878 349028 37884
rect 347872 10328 347924 10334
rect 347872 10270 347924 10276
rect 347884 4214 347912 10270
rect 349080 9042 349108 102054
rect 349540 100706 349568 102068
rect 350368 100858 350396 102068
rect 351210 102054 351868 102082
rect 350368 100830 350488 100858
rect 349528 100700 349580 100706
rect 349528 100642 349580 100648
rect 350356 100700 350408 100706
rect 350356 100642 350408 100648
rect 350368 47666 350396 100642
rect 350356 47660 350408 47666
rect 350356 47602 350408 47608
rect 350460 25566 350488 100830
rect 350540 43444 350592 43450
rect 350540 43386 350592 43392
rect 350448 25560 350500 25566
rect 350448 25502 350500 25508
rect 349068 9036 349120 9042
rect 349068 8978 349120 8984
rect 350264 7608 350316 7614
rect 350264 7550 350316 7556
rect 347872 4208 347924 4214
rect 347872 4150 347924 4156
rect 349068 4208 349120 4214
rect 349068 4150 349120 4156
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 343652 3454 344324 3482
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 347792 3454 347912 3482
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 3454
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 3454
rect 349080 480 349108 4150
rect 350276 480 350304 7550
rect 350552 3482 350580 43386
rect 351840 10402 351868 102054
rect 352024 99414 352052 102068
rect 352866 102054 353248 102082
rect 352012 99408 352064 99414
rect 352012 99350 352064 99356
rect 353116 99408 353168 99414
rect 353116 99350 353168 99356
rect 353128 49094 353156 99350
rect 353116 49088 353168 49094
rect 353116 49030 353168 49036
rect 353220 26926 353248 102054
rect 353680 99414 353708 102068
rect 354508 99498 354536 102068
rect 355258 102054 356008 102082
rect 355324 100156 355376 100162
rect 355324 100098 355376 100104
rect 354508 99470 354628 99498
rect 353668 99408 353720 99414
rect 353668 99350 353720 99356
rect 354496 99408 354548 99414
rect 354496 99350 354548 99356
rect 354508 93158 354536 99350
rect 354496 93152 354548 93158
rect 354496 93094 354548 93100
rect 353300 62824 353352 62830
rect 353300 62766 353352 62772
rect 353208 26920 353260 26926
rect 353208 26862 353260 26868
rect 351920 11824 351972 11830
rect 351920 11766 351972 11772
rect 351828 10396 351880 10402
rect 351828 10338 351880 10344
rect 351932 3482 351960 11766
rect 353312 3482 353340 62766
rect 354600 31142 354628 99470
rect 355336 60110 355364 100098
rect 355324 60104 355376 60110
rect 355324 60046 355376 60052
rect 354680 44872 354732 44878
rect 354680 44814 354732 44820
rect 354588 31136 354640 31142
rect 354588 31078 354640 31084
rect 354692 3482 354720 44814
rect 355980 42090 356008 102054
rect 356072 99414 356100 102068
rect 356914 102054 357388 102082
rect 356060 99408 356112 99414
rect 356060 99350 356112 99356
rect 357256 99408 357308 99414
rect 357256 99350 357308 99356
rect 357268 91798 357296 99350
rect 357256 91792 357308 91798
rect 357256 91734 357308 91740
rect 356060 73840 356112 73846
rect 356060 73782 356112 73788
rect 355968 42084 356020 42090
rect 355968 42026 356020 42032
rect 356072 3482 356100 73782
rect 357360 32502 357388 102054
rect 357728 99414 357756 102068
rect 357716 99408 357768 99414
rect 357716 99350 357768 99356
rect 358556 90370 358584 102068
rect 359384 99414 359412 102068
rect 360212 99414 360240 102068
rect 361040 99482 361068 102068
rect 361028 99476 361080 99482
rect 361028 99418 361080 99424
rect 361868 99414 361896 102068
rect 362710 102054 362908 102082
rect 363538 102054 364288 102082
rect 358728 99408 358780 99414
rect 358728 99350 358780 99356
rect 359372 99408 359424 99414
rect 359372 99350 359424 99356
rect 360108 99408 360160 99414
rect 360108 99350 360160 99356
rect 360200 99408 360252 99414
rect 360200 99350 360252 99356
rect 361488 99408 361540 99414
rect 361488 99350 361540 99356
rect 361856 99408 361908 99414
rect 361856 99350 361908 99356
rect 362776 99408 362828 99414
rect 362776 99350 362828 99356
rect 358544 90364 358596 90370
rect 358544 90306 358596 90312
rect 357440 46232 357492 46238
rect 357440 46174 357492 46180
rect 357348 32496 357400 32502
rect 357348 32438 357400 32444
rect 357348 8968 357400 8974
rect 357348 8910 357400 8916
rect 350552 3454 351408 3482
rect 351932 3454 352604 3482
rect 353312 3454 353800 3482
rect 354692 3454 354996 3482
rect 356072 3454 356192 3482
rect 351380 480 351408 3454
rect 352576 480 352604 3454
rect 353772 480 353800 3454
rect 354968 480 354996 3454
rect 356164 480 356192 3454
rect 357360 480 357388 8910
rect 357452 3482 357480 46174
rect 358740 6186 358768 99350
rect 358820 75200 358872 75206
rect 358820 75142 358872 75148
rect 358728 6180 358780 6186
rect 358728 6122 358780 6128
rect 358832 3482 358860 75142
rect 360120 33862 360148 99350
rect 360200 51740 360252 51746
rect 360200 51682 360252 51688
rect 360108 33856 360160 33862
rect 360108 33798 360160 33804
rect 360212 3482 360240 51682
rect 361500 28286 361528 99350
rect 362788 50454 362816 99350
rect 362776 50448 362828 50454
rect 362776 50390 362828 50396
rect 361580 29708 361632 29714
rect 361580 29650 361632 29656
rect 361488 28280 361540 28286
rect 361488 28222 361540 28228
rect 361592 3482 361620 29650
rect 362880 7614 362908 102054
rect 363604 99476 363656 99482
rect 363604 99418 363656 99424
rect 362960 13116 363012 13122
rect 362960 13058 363012 13064
rect 362868 7608 362920 7614
rect 362868 7550 362920 7556
rect 362972 3482 363000 13058
rect 363616 11830 363644 99418
rect 364260 89010 364288 102054
rect 364352 99482 364380 102068
rect 365194 102054 365668 102082
rect 364340 99476 364392 99482
rect 364340 99418 364392 99424
rect 364248 89004 364300 89010
rect 364248 88946 364300 88952
rect 364340 53100 364392 53106
rect 364340 53042 364392 53048
rect 363604 11824 363656 11830
rect 363604 11766 363656 11772
rect 364352 3482 364380 53042
rect 365640 43450 365668 102054
rect 366008 99414 366036 102068
rect 366850 102054 367048 102082
rect 365996 99408 366048 99414
rect 365996 99350 366048 99356
rect 366916 99408 366968 99414
rect 366916 99350 366968 99356
rect 366928 86290 366956 99350
rect 366916 86284 366968 86290
rect 366916 86226 366968 86232
rect 367020 53106 367048 102054
rect 367664 99414 367692 102068
rect 367744 99476 367796 99482
rect 367744 99418 367796 99424
rect 367652 99408 367704 99414
rect 367652 99350 367704 99356
rect 367008 53100 367060 53106
rect 367008 53042 367060 53048
rect 367756 51746 367784 99418
rect 368492 99414 368520 102068
rect 369334 102054 369808 102082
rect 370872 102070 370924 102076
rect 368388 99408 368440 99414
rect 368388 99350 368440 99356
rect 368480 99408 368532 99414
rect 368480 99350 368532 99356
rect 369676 99408 369728 99414
rect 369676 99350 369728 99356
rect 367744 51740 367796 51746
rect 367744 51682 367796 51688
rect 365720 47592 365772 47598
rect 365720 47534 365772 47540
rect 365628 43444 365680 43450
rect 365628 43386 365680 43392
rect 357452 3454 358584 3482
rect 358832 3454 359780 3482
rect 360212 3454 360976 3482
rect 361592 3454 362172 3482
rect 362972 3454 363368 3482
rect 364352 3454 364564 3482
rect 358556 480 358584 3454
rect 359752 480 359780 3454
rect 360948 480 360976 3454
rect 362144 480 362172 3454
rect 363340 480 363368 3454
rect 364536 480 364564 3454
rect 365732 480 365760 47534
rect 368400 44878 368428 99350
rect 369688 84862 369716 99350
rect 369676 84856 369728 84862
rect 369676 84798 369728 84804
rect 369780 54534 369808 102054
rect 370148 100706 370176 102068
rect 371818 102054 372568 102082
rect 370136 100700 370188 100706
rect 370136 100642 370188 100648
rect 371148 100700 371200 100706
rect 371148 100642 371200 100648
rect 370872 99340 370924 99346
rect 370872 99282 370924 99288
rect 370884 87009 370912 99282
rect 370686 87000 370742 87009
rect 370686 86935 370742 86944
rect 370870 87000 370926 87009
rect 370870 86935 370926 86944
rect 370700 83502 370728 86935
rect 370688 83496 370740 83502
rect 370688 83438 370740 83444
rect 369860 76628 369912 76634
rect 369860 76570 369912 76576
rect 369768 54528 369820 54534
rect 369768 54470 369820 54476
rect 368480 49020 368532 49026
rect 368480 48962 368532 48968
rect 368388 44872 368440 44878
rect 368388 44814 368440 44820
rect 367100 35216 367152 35222
rect 367100 35158 367152 35164
rect 365812 14476 365864 14482
rect 365812 14418 365864 14424
rect 365824 3482 365852 14418
rect 367112 3482 367140 35158
rect 368492 3482 368520 48962
rect 369872 3482 369900 76570
rect 371160 46238 371188 100642
rect 371240 64184 371292 64190
rect 371240 64126 371292 64132
rect 371148 46232 371200 46238
rect 371148 46174 371200 46180
rect 371252 3482 371280 64126
rect 372540 35222 372568 102054
rect 372632 100162 372660 102068
rect 373474 102054 373948 102082
rect 372620 100156 372672 100162
rect 372620 100098 372672 100104
rect 373816 100156 373868 100162
rect 373816 100098 373868 100104
rect 373828 47598 373856 100098
rect 373816 47592 373868 47598
rect 373816 47534 373868 47540
rect 372528 35216 372580 35222
rect 372528 35158 372580 35164
rect 372620 31068 372672 31074
rect 372620 31010 372672 31016
rect 372632 3482 372660 31010
rect 373920 13122 373948 102054
rect 374288 100706 374316 102068
rect 375130 102054 375328 102082
rect 374276 100700 374328 100706
rect 374276 100642 374328 100648
rect 375196 100700 375248 100706
rect 375196 100642 375248 100648
rect 375208 72486 375236 100642
rect 375196 72480 375248 72486
rect 375196 72422 375248 72428
rect 374000 69692 374052 69698
rect 374000 69634 374052 69640
rect 373908 13116 373960 13122
rect 373908 13058 373960 13064
rect 365824 3454 366956 3482
rect 367112 3454 368060 3482
rect 368492 3454 369256 3482
rect 369872 3454 370452 3482
rect 371252 3454 371648 3482
rect 372632 3454 372844 3482
rect 366928 480 366956 3454
rect 368032 480 368060 3454
rect 369228 480 369256 3454
rect 370424 480 370452 3454
rect 371620 480 371648 3454
rect 372816 480 372844 3454
rect 374012 3398 374040 69634
rect 374092 15904 374144 15910
rect 374092 15846 374144 15852
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 1442 374132 15846
rect 375300 8974 375328 102054
rect 375944 100706 375972 102068
rect 375932 100700 375984 100706
rect 375932 100642 375984 100648
rect 376668 100700 376720 100706
rect 376668 100642 376720 100648
rect 375380 82136 375432 82142
rect 375380 82078 375432 82084
rect 375288 8968 375340 8974
rect 375288 8910 375340 8916
rect 375392 3482 375420 82078
rect 376680 17270 376708 100642
rect 376772 99890 376800 102068
rect 377614 102054 378088 102082
rect 376760 99884 376812 99890
rect 376760 99826 376812 99832
rect 377956 99884 378008 99890
rect 377956 99826 378008 99832
rect 377968 71058 377996 99826
rect 377956 71052 378008 71058
rect 377956 70994 378008 71000
rect 378060 49026 378088 102054
rect 378336 99482 378364 102068
rect 379164 100230 379192 102068
rect 379152 100224 379204 100230
rect 379152 100166 379204 100172
rect 378324 99476 378376 99482
rect 378324 99418 378376 99424
rect 379992 99414 380020 102068
rect 379980 99408 380032 99414
rect 379980 99350 380032 99356
rect 380716 99408 380768 99414
rect 380716 99350 380768 99356
rect 378048 49020 378100 49026
rect 378048 48962 378100 48968
rect 379520 32428 379572 32434
rect 379520 32370 379572 32376
rect 376760 17400 376812 17406
rect 376760 17342 376812 17348
rect 376668 17264 376720 17270
rect 376668 17206 376720 17212
rect 376772 3482 376800 17342
rect 378140 11756 378192 11762
rect 378140 11698 378192 11704
rect 378152 3482 378180 11698
rect 379532 3482 379560 32370
rect 380728 31074 380756 99350
rect 380716 31068 380768 31074
rect 380716 31010 380768 31016
rect 380820 18630 380848 102068
rect 381662 102054 382228 102082
rect 381544 99476 381596 99482
rect 381544 99418 381596 99424
rect 381556 82142 381584 99418
rect 381544 82136 381596 82142
rect 381544 82078 381596 82084
rect 380900 77988 380952 77994
rect 380900 77930 380952 77936
rect 380808 18624 380860 18630
rect 380808 18566 380860 18572
rect 380912 3482 380940 77930
rect 382200 69698 382228 102054
rect 382476 99414 382504 102068
rect 383304 99482 383332 102068
rect 384132 100026 384160 102068
rect 384120 100020 384172 100026
rect 384120 99962 384172 99968
rect 383292 99476 383344 99482
rect 383292 99418 383344 99424
rect 382464 99408 382516 99414
rect 382464 99350 382516 99356
rect 383568 99408 383620 99414
rect 383568 99350 383620 99356
rect 382188 69692 382240 69698
rect 382188 69634 382240 69640
rect 382280 13184 382332 13190
rect 382280 13126 382332 13132
rect 382292 3482 382320 13126
rect 383580 10334 383608 99350
rect 383660 79348 383712 79354
rect 383660 79290 383712 79296
rect 383568 10328 383620 10334
rect 383568 10270 383620 10276
rect 383568 4888 383620 4894
rect 383568 4830 383620 4836
rect 375392 3454 376432 3482
rect 376772 3454 377628 3482
rect 378152 3454 378824 3482
rect 379532 3454 380020 3482
rect 380912 3454 381216 3482
rect 382292 3454 382412 3482
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3334
rect 376404 480 376432 3454
rect 377600 480 377628 3454
rect 378796 480 378824 3454
rect 379992 480 380020 3454
rect 381188 480 381216 3454
rect 382384 480 382412 3454
rect 383580 480 383608 4830
rect 383672 3482 383700 79290
rect 384960 32434 384988 102068
rect 385802 102054 386368 102082
rect 385684 99476 385736 99482
rect 385684 99418 385736 99424
rect 385040 87712 385092 87718
rect 385040 87654 385092 87660
rect 384948 32428 385000 32434
rect 384948 32370 385000 32376
rect 385052 3482 385080 87654
rect 385696 80714 385724 99418
rect 385684 80708 385736 80714
rect 385684 80650 385736 80656
rect 386340 14482 386368 102054
rect 386616 99414 386644 102068
rect 387458 102054 387748 102082
rect 386604 99408 386656 99414
rect 386604 99350 386656 99356
rect 387616 99408 387668 99414
rect 387616 99350 387668 99356
rect 387628 68338 387656 99350
rect 387616 68332 387668 68338
rect 387616 68274 387668 68280
rect 387720 33794 387748 102054
rect 388272 99414 388300 102068
rect 388260 99408 388312 99414
rect 388260 99350 388312 99356
rect 388996 99408 389048 99414
rect 388996 99350 389048 99356
rect 387800 80844 387852 80850
rect 387800 80786 387852 80792
rect 386420 33788 386472 33794
rect 386420 33730 386472 33736
rect 387708 33788 387760 33794
rect 387708 33730 387760 33736
rect 386328 14476 386380 14482
rect 386328 14418 386380 14424
rect 386432 3482 386460 33730
rect 387812 3482 387840 80786
rect 389008 79354 389036 99350
rect 388996 79348 389048 79354
rect 388996 79290 389048 79296
rect 389100 66910 389128 102068
rect 389942 102054 390508 102082
rect 389088 66904 389140 66910
rect 389088 66846 389140 66852
rect 390480 11762 390508 102054
rect 390756 99414 390784 102068
rect 391598 102054 391888 102082
rect 390744 99408 390796 99414
rect 390744 99350 390796 99356
rect 391756 99408 391808 99414
rect 391756 99350 391808 99356
rect 391768 77994 391796 99350
rect 391756 77988 391808 77994
rect 391756 77930 391808 77936
rect 391860 65550 391888 102054
rect 392412 100162 392440 102068
rect 392400 100156 392452 100162
rect 392400 100098 392452 100104
rect 393240 75206 393268 102068
rect 394082 102054 394648 102082
rect 393228 75200 393280 75206
rect 393228 75142 393280 75148
rect 391940 65680 391992 65686
rect 391940 65622 391992 65628
rect 391848 65544 391900 65550
rect 391848 65486 391900 65492
rect 390560 50380 390612 50386
rect 390560 50322 390612 50328
rect 390468 11756 390520 11762
rect 390468 11698 390520 11704
rect 389180 10464 389232 10470
rect 389180 10406 389232 10412
rect 389192 3482 389220 10406
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 386432 3454 387104 3482
rect 387812 3454 388300 3482
rect 389192 3454 389496 3482
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 3454
rect 388272 480 388300 3454
rect 389468 480 389496 3454
rect 390572 1578 390600 50322
rect 390652 18692 390704 18698
rect 390652 18634 390704 18640
rect 390664 3398 390692 18634
rect 391952 3482 391980 65622
rect 394620 57254 394648 102054
rect 394896 94518 394924 102068
rect 395738 102054 396028 102082
rect 394884 94512 394936 94518
rect 394884 94454 394936 94460
rect 396000 73846 396028 102054
rect 396552 99414 396580 102068
rect 396540 99408 396592 99414
rect 396540 99350 396592 99356
rect 395988 73840 396040 73846
rect 395988 73782 396040 73788
rect 394608 57248 394660 57254
rect 394608 57190 394660 57196
rect 393320 51808 393372 51814
rect 393320 51750 393372 51756
rect 393332 3482 393360 51750
rect 397380 50386 397408 102068
rect 398222 102054 398788 102082
rect 398104 99408 398156 99414
rect 398104 99350 398156 99356
rect 398116 64190 398144 99350
rect 398104 64184 398156 64190
rect 398104 64126 398156 64132
rect 397460 53168 397512 53174
rect 397460 53110 397512 53116
rect 397368 50380 397420 50386
rect 397368 50322 397420 50328
rect 394700 40792 394752 40798
rect 394700 40734 394752 40740
rect 394712 3482 394740 40734
rect 396080 17332 396132 17338
rect 396080 17274 396132 17280
rect 396092 3482 396120 17274
rect 397472 3482 397500 53110
rect 398760 15910 398788 102054
rect 399036 99414 399064 102068
rect 399878 102054 400076 102082
rect 399024 99408 399076 99414
rect 399024 99350 399076 99356
rect 400048 83570 400076 102054
rect 400128 99408 400180 99414
rect 400128 99350 400180 99356
rect 398840 83564 398892 83570
rect 398840 83506 398892 83512
rect 400036 83564 400088 83570
rect 400036 83506 400088 83512
rect 398748 15904 398800 15910
rect 398748 15846 398800 15852
rect 398852 3482 398880 83506
rect 400140 62830 400168 99350
rect 401600 84992 401652 84998
rect 401600 84934 401652 84940
rect 400128 62824 400180 62830
rect 400128 62766 400180 62772
rect 400220 54664 400272 54670
rect 400220 54606 400272 54612
rect 400232 4214 400260 54606
rect 400312 18760 400364 18766
rect 400312 18702 400364 18708
rect 400220 4208 400272 4214
rect 400220 4150 400272 4156
rect 400324 3482 400352 18702
rect 401324 4208 401376 4214
rect 401324 4150 401376 4156
rect 391952 3454 393084 3482
rect 393332 3454 394280 3482
rect 394712 3454 395476 3482
rect 396092 3454 396672 3482
rect 397472 3454 397868 3482
rect 398852 3454 399064 3482
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 1550 390692 1578
rect 390664 480 390692 1550
rect 391860 480 391888 3334
rect 393056 480 393084 3454
rect 394252 480 394280 3454
rect 395448 480 395476 3454
rect 396644 480 396672 3454
rect 397840 480 397868 3454
rect 399036 480 399064 3454
rect 400232 3454 400352 3482
rect 400232 480 400260 3454
rect 401336 480 401364 4150
rect 401612 3482 401640 84934
rect 402256 30326 402284 112639
rect 402348 41410 402376 119711
rect 402440 77246 402468 133991
rect 402532 88330 402560 141063
rect 402624 111790 402652 148271
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 578884 125656 578936 125662
rect 578884 125598 578936 125604
rect 402612 111784 402664 111790
rect 402612 111726 402664 111732
rect 555424 104916 555476 104922
rect 555424 104858 555476 104864
rect 403624 100224 403676 100230
rect 403624 100166 403676 100172
rect 402520 88324 402572 88330
rect 402520 88266 402572 88272
rect 402980 80776 403032 80782
rect 402980 80718 403032 80724
rect 402428 77240 402480 77246
rect 402428 77182 402480 77188
rect 402336 41404 402388 41410
rect 402336 41346 402388 41352
rect 402244 30320 402296 30326
rect 402244 30262 402296 30268
rect 402992 3482 403020 80718
rect 403636 55894 403664 100166
rect 446404 100156 446456 100162
rect 446404 100098 446456 100104
rect 420184 100088 420236 100094
rect 420184 100030 420236 100036
rect 405740 94648 405792 94654
rect 405740 94590 405792 94596
rect 404360 87644 404412 87650
rect 404360 87586 404412 87592
rect 403624 55888 403676 55894
rect 403624 55830 403676 55836
rect 404372 3482 404400 87586
rect 405752 3482 405780 94590
rect 416780 90432 416832 90438
rect 416780 90374 416832 90380
rect 412640 89140 412692 89146
rect 412640 89082 412692 89088
rect 408500 86352 408552 86358
rect 408500 86294 408552 86300
rect 407120 67040 407172 67046
rect 407120 66982 407172 66988
rect 407132 3482 407160 66982
rect 408512 4214 408540 86294
rect 411260 72548 411312 72554
rect 411260 72490 411312 72496
rect 409880 54596 409932 54602
rect 409880 54538 409932 54544
rect 408592 35284 408644 35290
rect 408592 35226 408644 35232
rect 408500 4208 408552 4214
rect 408500 4150 408552 4156
rect 408604 3482 408632 35226
rect 409696 4208 409748 4214
rect 409696 4150 409748 4156
rect 401612 3454 402560 3482
rect 402992 3454 403756 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 407132 3454 407344 3482
rect 402532 480 402560 3454
rect 403728 480 403756 3454
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407316 480 407344 3454
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 4150
rect 409892 3482 409920 54538
rect 411272 3482 411300 72490
rect 412652 3482 412680 89082
rect 415400 71188 415452 71194
rect 415400 71130 415452 71136
rect 414020 40724 414072 40730
rect 414020 40666 414072 40672
rect 414032 3482 414060 40666
rect 415412 3482 415440 71130
rect 416792 3482 416820 90374
rect 416872 57384 416924 57390
rect 416872 57326 416924 57332
rect 416884 3618 416912 57326
rect 418160 56024 418212 56030
rect 418160 55966 418212 55972
rect 416884 3590 418016 3618
rect 409892 3454 410932 3482
rect 411272 3454 412128 3482
rect 412652 3454 413324 3482
rect 414032 3454 414520 3482
rect 415412 3454 415716 3482
rect 416792 3454 416912 3482
rect 410904 480 410932 3454
rect 412100 480 412128 3454
rect 413296 480 413324 3454
rect 414492 480 414520 3454
rect 415688 480 415716 3454
rect 416884 480 416912 3454
rect 417988 480 418016 3590
rect 418172 3482 418200 55966
rect 419540 29640 419592 29646
rect 419540 29582 419592 29588
rect 419552 3618 419580 29582
rect 420196 4894 420224 100030
rect 444380 96008 444432 96014
rect 444380 95950 444432 95956
rect 430580 93220 430632 93226
rect 430580 93162 430632 93168
rect 423680 91860 423732 91866
rect 423680 91802 423732 91808
rect 420920 84924 420972 84930
rect 420920 84866 420972 84872
rect 420184 4888 420236 4894
rect 420184 4830 420236 4836
rect 419552 3590 420408 3618
rect 418172 3454 419212 3482
rect 419184 480 419212 3454
rect 420380 480 420408 3590
rect 420932 3482 420960 84866
rect 422300 69760 422352 69766
rect 422300 69702 422352 69708
rect 422312 3482 422340 69702
rect 423692 3482 423720 91802
rect 427820 86420 427872 86426
rect 427820 86362 427872 86368
rect 426440 73908 426492 73914
rect 426440 73850 426492 73856
rect 425060 68468 425112 68474
rect 425060 68410 425112 68416
rect 420932 3454 421604 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 421576 480 421604 3454
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425072 3398 425100 68410
rect 425152 15972 425204 15978
rect 425152 15914 425204 15920
rect 425060 3392 425112 3398
rect 425060 3334 425112 3340
rect 425164 480 425192 15914
rect 426452 3482 426480 73850
rect 427832 3482 427860 86362
rect 429200 66972 429252 66978
rect 429200 66914 429252 66920
rect 429212 3482 429240 66914
rect 430592 3482 430620 93162
rect 434720 89072 434772 89078
rect 434720 89014 434772 89020
rect 433340 65612 433392 65618
rect 433340 65554 433392 65560
rect 431960 55956 432012 55962
rect 431960 55898 432012 55904
rect 431972 3482 432000 55898
rect 433352 3482 433380 65554
rect 434628 4820 434680 4826
rect 434628 4762 434680 4768
rect 426452 3454 427584 3482
rect 427832 3454 428780 3482
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 431972 3454 432368 3482
rect 433352 3454 433564 3482
rect 426348 3392 426400 3398
rect 426348 3334 426400 3340
rect 426360 480 426388 3334
rect 427556 480 427584 3454
rect 428752 480 428780 3454
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3454
rect 433536 480 433564 3454
rect 434640 480 434668 4762
rect 434732 3482 434760 89014
rect 441620 76560 441672 76566
rect 441620 76502 441672 76508
rect 437480 75268 437532 75274
rect 437480 75210 437532 75216
rect 436100 57316 436152 57322
rect 436100 57258 436152 57264
rect 436112 3482 436140 57258
rect 437492 3482 437520 75210
rect 438860 68400 438912 68406
rect 438860 68342 438912 68348
rect 438872 3482 438900 68342
rect 440240 64252 440292 64258
rect 440240 64194 440292 64200
rect 440252 3482 440280 64194
rect 441632 3482 441660 76502
rect 443000 71120 443052 71126
rect 443000 71062 443052 71068
rect 434732 3454 435864 3482
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 435836 480 435864 3454
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 71062
rect 443092 20052 443144 20058
rect 443092 19994 443144 20000
rect 443104 3482 443132 19994
rect 444392 3482 444420 95950
rect 446416 20058 446444 100098
rect 493324 100020 493376 100026
rect 493324 99962 493376 99968
rect 462320 98728 462372 98734
rect 462320 98670 462372 98676
rect 455420 97368 455472 97374
rect 455420 97310 455472 97316
rect 448520 78056 448572 78062
rect 448520 77998 448572 78004
rect 447140 62892 447192 62898
rect 447140 62834 447192 62840
rect 446404 20052 446456 20058
rect 446404 19994 446456 20000
rect 446588 4140 446640 4146
rect 446588 4082 446640 4088
rect 443104 3454 444236 3482
rect 444392 3454 445432 3482
rect 444208 480 444236 3454
rect 445404 480 445432 3454
rect 446600 480 446628 4082
rect 447152 3482 447180 62834
rect 448532 3482 448560 77998
rect 451280 61464 451332 61470
rect 451280 61406 451332 61412
rect 450176 4072 450228 4078
rect 450176 4014 450228 4020
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 4014
rect 451292 480 451320 61406
rect 454040 21480 454092 21486
rect 454040 21422 454092 21428
rect 451372 16040 451424 16046
rect 451372 15982 451424 15988
rect 451384 3482 451412 15982
rect 453672 4004 453724 4010
rect 453672 3946 453724 3952
rect 451384 3454 452516 3482
rect 452488 480 452516 3454
rect 453684 480 453712 3946
rect 454052 3482 454080 21422
rect 455432 3482 455460 97310
rect 459652 82204 459704 82210
rect 459652 82146 459704 82152
rect 458180 36644 458232 36650
rect 458180 36586 458232 36592
rect 457260 3868 457312 3874
rect 457260 3810 457312 3816
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3810
rect 458192 3482 458220 36586
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 82146
rect 460940 60036 460992 60042
rect 460940 59978 460992 59984
rect 460848 3936 460900 3942
rect 460848 3878 460900 3884
rect 460860 480 460888 3878
rect 460952 3482 460980 59978
rect 462332 3482 462360 98670
rect 485780 98660 485832 98666
rect 485780 98602 485832 98608
rect 482284 83564 482336 83570
rect 482284 83506 482336 83512
rect 480260 79416 480312 79422
rect 480260 79358 480312 79364
rect 469220 61396 469272 61402
rect 469220 61338 469272 61344
rect 465080 58744 465132 58750
rect 465080 58686 465132 58692
rect 464436 3800 464488 3806
rect 464436 3742 464488 3748
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3742
rect 465092 3482 465120 58686
rect 467932 22840 467984 22846
rect 467932 22782 467984 22788
rect 466460 19984 466512 19990
rect 466460 19926 466512 19932
rect 466472 3482 466500 19926
rect 467840 3732 467892 3738
rect 467840 3674 467892 3680
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 3210 467880 3674
rect 467944 3398 467972 22782
rect 469232 3482 469260 61338
rect 476120 39432 476172 39438
rect 476120 39374 476172 39380
rect 471980 24200 472032 24206
rect 471980 24142 472032 24148
rect 471520 3664 471572 3670
rect 471520 3606 471572 3612
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 3182 467972 3210
rect 467944 480 467972 3182
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3606
rect 471992 3482 472020 24142
rect 473360 21412 473412 21418
rect 473360 21354 473412 21360
rect 473372 3482 473400 21354
rect 475108 3596 475160 3602
rect 475108 3538 475160 3544
rect 471992 3454 472756 3482
rect 473372 3454 473952 3482
rect 472728 480 472756 3454
rect 473924 480 473952 3454
rect 475120 480 475148 3538
rect 476132 3482 476160 39374
rect 478880 38004 478932 38010
rect 478880 37946 478932 37952
rect 477592 36576 477644 36582
rect 477592 36518 477644 36524
rect 477604 3482 477632 36518
rect 476132 3454 476344 3482
rect 476316 480 476344 3454
rect 477512 3454 477632 3482
rect 478696 3528 478748 3534
rect 478696 3470 478748 3476
rect 478892 3482 478920 37946
rect 480272 3482 480300 79358
rect 482296 9194 482324 83506
rect 484400 25628 484452 25634
rect 484400 25570 484452 25576
rect 482204 9166 482324 9194
rect 482204 7342 482232 9166
rect 482192 7336 482244 7342
rect 482192 7278 482244 7284
rect 483480 4888 483532 4894
rect 483480 4830 483532 4836
rect 477512 480 477540 3454
rect 478708 480 478736 3470
rect 478892 3454 479932 3482
rect 480272 3454 481128 3482
rect 479904 480 479932 3454
rect 481100 480 481128 3454
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 482296 480 482324 3402
rect 483492 480 483520 4830
rect 484412 3482 484440 25570
rect 485792 7546 485820 98602
rect 488540 60104 488592 60110
rect 488540 60046 488592 60052
rect 487160 26988 487212 26994
rect 487160 26930 487212 26936
rect 485872 14544 485924 14550
rect 485872 14486 485924 14492
rect 485780 7540 485832 7546
rect 485780 7482 485832 7488
rect 485884 7426 485912 14486
rect 487172 12442 487200 26930
rect 488552 12442 488580 60046
rect 491300 28348 491352 28354
rect 491300 28290 491352 28296
rect 491312 19310 491340 28290
rect 492680 22772 492732 22778
rect 492680 22714 492732 22720
rect 492692 19310 492720 22714
rect 491300 19304 491352 19310
rect 491300 19246 491352 19252
rect 492680 19304 492732 19310
rect 492680 19246 492732 19252
rect 487160 12436 487212 12442
rect 487160 12378 487212 12384
rect 488172 12436 488224 12442
rect 488172 12378 488224 12384
rect 488540 12436 488592 12442
rect 488540 12378 488592 12384
rect 489368 12436 489420 12442
rect 489368 12378 489420 12384
rect 486976 7540 487028 7546
rect 486976 7482 487028 7488
rect 485792 7398 485912 7426
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 480 485820 7398
rect 486988 480 487016 7482
rect 488184 480 488212 12378
rect 489380 480 489408 12378
rect 491760 9716 491812 9722
rect 491760 9658 491812 9664
rect 492956 9716 493008 9722
rect 492956 9658 493008 9664
rect 490564 6248 490616 6254
rect 490564 6190 490616 6196
rect 490576 480 490604 6190
rect 491772 480 491800 9658
rect 492968 480 492996 9658
rect 493336 4826 493364 99962
rect 496820 97300 496872 97306
rect 496820 97242 496872 97248
rect 495440 58676 495492 58682
rect 495440 58618 495492 58624
rect 494060 42152 494112 42158
rect 494060 42094 494112 42100
rect 494072 7682 494100 42094
rect 494152 7744 494204 7750
rect 494152 7686 494204 7692
rect 494060 7676 494112 7682
rect 494060 7618 494112 7624
rect 493324 4820 493376 4826
rect 493324 4762 493376 4768
rect 494164 480 494192 7686
rect 495348 7676 495400 7682
rect 495348 7618 495400 7624
rect 495360 480 495388 7618
rect 495452 3482 495480 58618
rect 496832 3482 496860 97242
rect 500960 95940 501012 95946
rect 500960 95882 501012 95888
rect 498200 43512 498252 43518
rect 498200 43454 498252 43460
rect 498212 3482 498240 43454
rect 499580 24132 499632 24138
rect 499580 24074 499632 24080
rect 499592 3482 499620 24074
rect 500972 3482 501000 95882
rect 503720 94580 503772 94586
rect 503720 94522 503772 94528
rect 502340 44940 502392 44946
rect 502340 44882 502392 44888
rect 502352 3482 502380 44882
rect 502432 39364 502484 39370
rect 502432 39306 502484 39312
rect 502444 3602 502472 39306
rect 502432 3596 502484 3602
rect 502432 3538 502484 3544
rect 503628 3596 503680 3602
rect 503628 3538 503680 3544
rect 495452 3454 496584 3482
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 499592 3454 500172 3482
rect 500972 3454 501276 3482
rect 502352 3454 502472 3482
rect 496556 480 496584 3454
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 500144 480 500172 3454
rect 501248 480 501276 3454
rect 502444 480 502472 3454
rect 503640 480 503668 3538
rect 503732 3482 503760 94522
rect 514760 93152 514812 93158
rect 514760 93094 514812 93100
rect 512000 49088 512052 49094
rect 512000 49030 512052 49036
rect 509240 47660 509292 47666
rect 509240 47602 509292 47608
rect 509252 46918 509280 47602
rect 509240 46912 509292 46918
rect 509240 46854 509292 46860
rect 505100 46300 505152 46306
rect 505100 46242 505152 46248
rect 505112 12442 505140 46242
rect 506480 37936 506532 37942
rect 506480 37878 506532 37884
rect 506492 12442 506520 37878
rect 509240 37324 509292 37330
rect 509240 37266 509292 37272
rect 509252 27606 509280 37266
rect 509240 27600 509292 27606
rect 509240 27542 509292 27548
rect 510712 25560 510764 25566
rect 510712 25502 510764 25508
rect 510724 19394 510752 25502
rect 510632 19366 510752 19394
rect 510632 19310 510660 19366
rect 510620 19304 510672 19310
rect 510620 19246 510672 19252
rect 505100 12436 505152 12442
rect 505100 12378 505152 12384
rect 506020 12436 506072 12442
rect 506020 12378 506072 12384
rect 506480 12436 506532 12442
rect 506480 12378 506532 12384
rect 507216 12436 507268 12442
rect 507216 12378 507268 12384
rect 503732 3454 504864 3482
rect 504836 480 504864 3454
rect 506032 480 506060 12378
rect 507228 480 507256 12378
rect 509608 9716 509660 9722
rect 509608 9658 509660 9664
rect 510804 9716 510856 9722
rect 510804 9658 510856 9664
rect 508412 9036 508464 9042
rect 508412 8978 508464 8984
rect 508424 480 508452 8978
rect 509620 480 509648 9658
rect 510816 480 510844 9658
rect 512012 7682 512040 49030
rect 513380 26920 513432 26926
rect 513380 26862 513432 26868
rect 513392 12442 513420 26862
rect 514772 12442 514800 93094
rect 518900 91792 518952 91798
rect 518900 91734 518952 91740
rect 518912 85542 518940 91734
rect 521660 90364 521712 90370
rect 521660 90306 521712 90312
rect 518900 85536 518952 85542
rect 518900 85478 518952 85484
rect 518900 75948 518952 75954
rect 518900 75890 518952 75896
rect 518912 66230 518940 75890
rect 518900 66224 518952 66230
rect 518900 66166 518952 66172
rect 518900 56636 518952 56642
rect 518900 56578 518952 56584
rect 518912 46918 518940 56578
rect 518900 46912 518952 46918
rect 518900 46854 518952 46860
rect 517520 42084 517572 42090
rect 517520 42026 517572 42032
rect 516140 31136 516192 31142
rect 516140 31078 516192 31084
rect 516152 19310 516180 31078
rect 516140 19304 516192 19310
rect 516140 19246 516192 19252
rect 517532 12510 517560 42026
rect 518900 37324 518952 37330
rect 518900 37266 518952 37272
rect 518912 27606 518940 37266
rect 520280 32496 520332 32502
rect 520280 32438 520332 32444
rect 518900 27600 518952 27606
rect 518900 27542 518952 27548
rect 518900 18012 518952 18018
rect 518900 17954 518952 17960
rect 518912 12510 518940 17954
rect 517520 12504 517572 12510
rect 517520 12446 517572 12452
rect 518900 12504 518952 12510
rect 518900 12446 518952 12452
rect 513380 12436 513432 12442
rect 513380 12378 513432 12384
rect 514392 12436 514444 12442
rect 514392 12378 514444 12384
rect 514760 12436 514812 12442
rect 514760 12378 514812 12384
rect 515588 12436 515640 12442
rect 515588 12378 515640 12384
rect 512092 10396 512144 10402
rect 512092 10338 512144 10344
rect 512000 7676 512052 7682
rect 512000 7618 512052 7624
rect 512104 1442 512132 10338
rect 513196 7676 513248 7682
rect 513196 7618 513248 7624
rect 512012 1414 512132 1442
rect 512012 480 512040 1414
rect 513208 480 513236 7618
rect 514404 480 514432 12378
rect 515600 480 515628 12378
rect 517888 12368 517940 12374
rect 517888 12310 517940 12316
rect 519084 12368 519136 12374
rect 519084 12310 519136 12316
rect 516784 9716 516836 9722
rect 516784 9658 516836 9664
rect 516796 480 516824 9658
rect 517900 9654 517928 12310
rect 519096 9654 519124 12310
rect 517888 9648 517940 9654
rect 517888 9590 517940 9596
rect 519084 9648 519136 9654
rect 519084 9590 519136 9596
rect 517888 604 517940 610
rect 517888 546 517940 552
rect 519084 604 519136 610
rect 519084 546 519136 552
rect 517900 480 517928 546
rect 519096 480 519124 546
rect 520292 480 520320 32438
rect 521672 12442 521700 90306
rect 528560 89004 528612 89010
rect 528560 88946 528612 88952
rect 527180 50448 527232 50454
rect 527180 50390 527232 50396
rect 527192 46918 527220 50390
rect 527180 46912 527232 46918
rect 527180 46854 527232 46860
rect 527180 37324 527232 37330
rect 527180 37266 527232 37272
rect 523040 33856 523092 33862
rect 523040 33798 523092 33804
rect 523052 12442 523080 33798
rect 524512 28280 524564 28286
rect 524512 28222 524564 28228
rect 524524 19394 524552 28222
rect 527192 27606 527220 37266
rect 527180 27600 527232 27606
rect 527180 27542 527232 27548
rect 524432 19366 524552 19394
rect 524432 12510 524460 19366
rect 527180 18012 527232 18018
rect 527180 17954 527232 17960
rect 527192 14890 527220 17954
rect 527180 14884 527232 14890
rect 527180 14826 527232 14832
rect 527364 14884 527416 14890
rect 527364 14826 527416 14832
rect 524420 12504 524472 12510
rect 524420 12446 524472 12452
rect 521660 12436 521712 12442
rect 521660 12378 521712 12384
rect 522672 12436 522724 12442
rect 522672 12378 522724 12384
rect 523040 12436 523092 12442
rect 523040 12378 523092 12384
rect 523868 12436 523920 12442
rect 523868 12378 523920 12384
rect 521476 6180 521528 6186
rect 521476 6122 521528 6128
rect 521488 480 521516 6122
rect 522684 480 522712 12378
rect 523880 480 523908 12378
rect 525064 12368 525116 12374
rect 525064 12310 525116 12316
rect 527376 12322 527404 14826
rect 525076 9654 525104 12310
rect 527376 12294 527496 12322
rect 526260 11824 526312 11830
rect 526260 11766 526312 11772
rect 525064 9648 525116 9654
rect 525064 9590 525116 9596
rect 525064 9512 525116 9518
rect 525064 9454 525116 9460
rect 525076 480 525104 9454
rect 526272 480 526300 11766
rect 527468 9654 527496 12294
rect 527456 9648 527508 9654
rect 527456 9590 527508 9596
rect 527456 9512 527508 9518
rect 527456 9454 527508 9460
rect 527468 480 527496 9454
rect 528572 7614 528600 88946
rect 532700 86284 532752 86290
rect 532700 86226 532752 86232
rect 532712 85542 532740 86226
rect 532700 85536 532752 85542
rect 532700 85478 532752 85484
rect 536840 84856 536892 84862
rect 536840 84798 536892 84804
rect 532700 75948 532752 75954
rect 532700 75890 532752 75896
rect 532712 66230 532740 75890
rect 532700 66224 532752 66230
rect 532700 66166 532752 66172
rect 532700 56636 532752 56642
rect 532700 56578 532752 56584
rect 529940 51740 529992 51746
rect 529940 51682 529992 51688
rect 529952 12442 529980 51682
rect 532712 46918 532740 56578
rect 534080 53100 534132 53106
rect 534080 53042 534132 53048
rect 532700 46912 532752 46918
rect 532700 46854 532752 46860
rect 531320 43444 531372 43450
rect 531320 43386 531372 43392
rect 531332 12442 531360 43386
rect 532700 37324 532752 37330
rect 532700 37266 532752 37272
rect 532712 27606 532740 37266
rect 532700 27600 532752 27606
rect 532700 27542 532752 27548
rect 529940 12436 529992 12442
rect 529940 12378 529992 12384
rect 531044 12436 531096 12442
rect 531044 12378 531096 12384
rect 531320 12436 531372 12442
rect 531320 12378 531372 12384
rect 532240 12436 532292 12442
rect 532240 12378 532292 12384
rect 528560 7608 528612 7614
rect 528560 7550 528612 7556
rect 529848 7608 529900 7614
rect 529848 7550 529900 7556
rect 528652 7540 528704 7546
rect 528652 7482 528704 7488
rect 528664 480 528692 7482
rect 529860 480 529888 7550
rect 531056 480 531084 12378
rect 532252 480 532280 12378
rect 533436 9716 533488 9722
rect 533436 9658 533488 9664
rect 533448 480 533476 9658
rect 534092 3482 534120 53042
rect 535460 44872 535512 44878
rect 535460 44814 535512 44820
rect 535472 3482 535500 44814
rect 536852 3482 536880 84798
rect 539600 83496 539652 83502
rect 539600 83438 539652 83444
rect 536932 54528 536984 54534
rect 536932 54470 536984 54476
rect 536944 3602 536972 54470
rect 538220 46232 538272 46238
rect 538220 46174 538272 46180
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 538128 3596 538180 3602
rect 538128 3538 538180 3544
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 3538
rect 538232 3346 538260 46174
rect 539612 3346 539640 83438
rect 550640 82136 550692 82142
rect 550640 82078 550692 82084
rect 550652 77217 550680 82078
rect 550638 77208 550694 77217
rect 550638 77143 550694 77152
rect 550914 77208 550970 77217
rect 550914 77143 550970 77152
rect 545120 72480 545172 72486
rect 545120 72422 545172 72428
rect 542360 47592 542412 47598
rect 542360 47534 542412 47540
rect 540980 35216 541032 35222
rect 540980 35158 541032 35164
rect 540992 3346 541020 35158
rect 542372 3346 542400 47534
rect 544108 13116 544160 13122
rect 544108 13058 544160 13064
rect 538232 3318 539364 3346
rect 539612 3318 540560 3346
rect 540992 3318 541756 3346
rect 542372 3318 542952 3346
rect 539336 480 539364 3318
rect 540532 480 540560 3318
rect 541728 480 541756 3318
rect 542924 480 542952 3318
rect 544120 480 544148 13058
rect 545132 12510 545160 72422
rect 547880 71052 547932 71058
rect 547880 70994 547932 71000
rect 547892 19310 547920 70994
rect 550928 67658 550956 77143
rect 554780 69692 554832 69698
rect 554780 69634 554832 69640
rect 550640 67652 550692 67658
rect 550640 67594 550692 67600
rect 550916 67652 550968 67658
rect 550916 67594 550968 67600
rect 550652 58177 550680 67594
rect 550638 58168 550694 58177
rect 550638 58103 550694 58112
rect 550638 58032 550694 58041
rect 550638 57967 550694 57976
rect 549260 49020 549312 49026
rect 549260 48962 549312 48968
rect 547880 19304 547932 19310
rect 547880 19246 547932 19252
rect 548892 19304 548944 19310
rect 548892 19246 548944 19252
rect 546500 17264 546552 17270
rect 546500 17206 546552 17212
rect 545120 12504 545172 12510
rect 545120 12446 545172 12452
rect 545304 12368 545356 12374
rect 545304 12310 545356 12316
rect 545316 9654 545344 12310
rect 545304 9648 545356 9654
rect 545304 9590 545356 9596
rect 546512 7614 546540 17206
rect 548904 9654 548932 19246
rect 549272 12442 549300 48962
rect 550652 19310 550680 57967
rect 552020 55888 552072 55894
rect 552020 55830 552072 55836
rect 550640 19304 550692 19310
rect 550640 19246 550692 19252
rect 552032 14498 552060 55830
rect 553400 31068 553452 31074
rect 553400 31010 553452 31016
rect 553412 19310 553440 31010
rect 553400 19304 553452 19310
rect 553400 19246 553452 19252
rect 552032 14470 552152 14498
rect 549260 12436 549312 12442
rect 549260 12378 549312 12384
rect 550088 12436 550140 12442
rect 550088 12378 550140 12384
rect 550100 9654 550128 12378
rect 552124 12374 552152 14470
rect 551192 12368 551244 12374
rect 551192 12310 551244 12316
rect 552112 12368 552164 12374
rect 552112 12310 552164 12316
rect 552388 12368 552440 12374
rect 552388 12310 552440 12316
rect 548892 9648 548944 9654
rect 548892 9590 548944 9596
rect 550088 9648 550140 9654
rect 550088 9590 550140 9596
rect 546592 8968 546644 8974
rect 546592 8910 546644 8916
rect 546500 7608 546552 7614
rect 546500 7550 546552 7556
rect 546604 7426 546632 8910
rect 547696 7608 547748 7614
rect 547696 7550 547748 7556
rect 546512 7398 546632 7426
rect 545304 604 545356 610
rect 545304 546 545356 552
rect 545316 480 545344 546
rect 546512 480 546540 7398
rect 547708 480 547736 7550
rect 548892 604 548944 610
rect 548892 546 548944 552
rect 550088 604 550140 610
rect 550088 546 550140 552
rect 548904 480 548932 546
rect 550100 480 550128 546
rect 551204 480 551232 12310
rect 552400 480 552428 12310
rect 553584 9716 553636 9722
rect 553584 9658 553636 9664
rect 553596 480 553624 9658
rect 554792 7614 554820 69634
rect 554872 18624 554924 18630
rect 554872 18566 554924 18572
rect 554780 7608 554832 7614
rect 554780 7550 554832 7556
rect 554884 7426 554912 18566
rect 555436 17950 555464 104858
rect 574100 94512 574152 94518
rect 574100 94454 574152 94460
rect 557540 80708 557592 80714
rect 557540 80650 557592 80656
rect 555424 17944 555476 17950
rect 555424 17886 555476 17892
rect 557552 12442 557580 80650
rect 564440 79348 564492 79354
rect 564440 79290 564492 79296
rect 563060 68332 563112 68338
rect 563060 68274 563112 68280
rect 560300 32428 560352 32434
rect 560300 32370 560352 32376
rect 560312 19310 560340 32370
rect 560300 19304 560352 19310
rect 560300 19246 560352 19252
rect 560760 19304 560812 19310
rect 560760 19246 560812 19252
rect 557540 12436 557592 12442
rect 557540 12378 557592 12384
rect 558368 12436 558420 12442
rect 558368 12378 558420 12384
rect 557172 10328 557224 10334
rect 557172 10270 557224 10276
rect 555976 7608 556028 7614
rect 555976 7550 556028 7556
rect 554792 7398 554912 7426
rect 554792 480 554820 7398
rect 555988 480 556016 7550
rect 557184 480 557212 10270
rect 558380 480 558408 12378
rect 559564 4820 559616 4826
rect 559564 4762 559616 4768
rect 559576 480 559604 4762
rect 560772 480 560800 19246
rect 561956 14476 562008 14482
rect 561956 14418 562008 14424
rect 561968 480 561996 14418
rect 563072 7426 563100 68274
rect 563152 33788 563204 33794
rect 563152 33730 563204 33736
rect 563164 7614 563192 33730
rect 564452 12442 564480 79290
rect 568580 77988 568632 77994
rect 568580 77930 568632 77936
rect 565820 66904 565872 66910
rect 565820 66846 565872 66852
rect 565832 12442 565860 66846
rect 567936 50380 567988 50386
rect 567936 50322 567988 50328
rect 567948 48278 567976 50322
rect 568592 48521 568620 77930
rect 571340 75200 571392 75206
rect 571340 75142 571392 75148
rect 569960 56636 570012 56642
rect 569960 56578 570012 56584
rect 568578 48512 568634 48521
rect 568578 48447 568634 48456
rect 568578 48376 568634 48385
rect 568578 48311 568634 48320
rect 567936 48272 567988 48278
rect 567936 48214 567988 48220
rect 567844 38684 567896 38690
rect 567844 38626 567896 38632
rect 567856 31754 567884 38626
rect 567844 31748 567896 31754
rect 567844 31690 567896 31696
rect 568028 31748 568080 31754
rect 568028 31690 568080 31696
rect 568040 27606 568068 31690
rect 568028 27600 568080 27606
rect 568028 27542 568080 27548
rect 568028 18012 568080 18018
rect 568028 17954 568080 17960
rect 564440 12436 564492 12442
rect 564440 12378 564492 12384
rect 565544 12436 565596 12442
rect 565544 12378 565596 12384
rect 565820 12436 565872 12442
rect 565820 12378 565872 12384
rect 566740 12436 566792 12442
rect 566740 12378 566792 12384
rect 563152 7608 563204 7614
rect 563152 7550 563204 7556
rect 564348 7608 564400 7614
rect 564348 7550 564400 7556
rect 563072 7398 563192 7426
rect 563164 480 563192 7398
rect 564360 480 564388 7550
rect 565556 480 565584 12378
rect 566752 480 566780 12378
rect 567844 11756 567896 11762
rect 567844 11698 567896 11704
rect 567856 480 567884 11698
rect 568040 8265 568068 17954
rect 568592 12510 568620 48311
rect 569972 46918 570000 56578
rect 569960 46912 570012 46918
rect 569960 46854 570012 46860
rect 569960 37324 570012 37330
rect 569960 37266 570012 37272
rect 569972 27606 570000 37266
rect 569960 27600 570012 27606
rect 569960 27542 570012 27548
rect 568580 12504 568632 12510
rect 568580 12446 568632 12452
rect 569040 12436 569092 12442
rect 569040 12378 569092 12384
rect 568026 8256 568082 8265
rect 568026 8191 568082 8200
rect 568210 8120 568266 8129
rect 568210 8055 568266 8064
rect 568224 3602 568252 8055
rect 568212 3596 568264 3602
rect 568212 3538 568264 3544
rect 569052 480 569080 12378
rect 570236 9716 570288 9722
rect 570236 9658 570288 9664
rect 570248 480 570276 9658
rect 571352 7614 571380 75142
rect 572720 57248 572772 57254
rect 572720 57190 572772 57196
rect 571432 20052 571484 20058
rect 571432 19994 571484 20000
rect 571340 7608 571392 7614
rect 571340 7550 571392 7556
rect 571444 480 571472 19994
rect 572628 7608 572680 7614
rect 572628 7550 572680 7556
rect 572640 480 572668 7550
rect 572732 3618 572760 57190
rect 574112 3618 574140 94454
rect 575480 73840 575532 73846
rect 575480 73782 575532 73788
rect 575492 3618 575520 73782
rect 578896 64569 578924 125598
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 578882 64560 578938 64569
rect 578882 64495 578938 64504
rect 576860 64184 576912 64190
rect 576860 64126 576912 64132
rect 572732 3590 573864 3618
rect 574112 3590 575060 3618
rect 575492 3590 576256 3618
rect 573836 480 573864 3590
rect 575032 480 575060 3590
rect 576228 480 576256 3590
rect 576872 610 576900 64126
rect 578884 62824 578936 62830
rect 578884 62766 578936 62772
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 576860 604 576912 610
rect 576860 546 576912 552
rect 577412 604 577464 610
rect 577412 546 577464 552
rect 577424 480 577452 546
rect 578620 480 578648 3470
rect 578896 3194 578924 62766
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 578976 15904 579028 15910
rect 578976 15846 579028 15852
rect 578988 3534 579016 15846
rect 578976 3528 579028 3534
rect 578976 3470 579028 3476
rect 579804 3528 579856 3534
rect 579804 3470 579856 3476
rect 578884 3188 578936 3194
rect 578884 3130 578936 3136
rect 579816 480 579844 3470
rect 582196 3324 582248 3330
rect 582196 3266 582248 3272
rect 581000 3188 581052 3194
rect 581000 3130 581052 3136
rect 581012 480 581040 3130
rect 582208 480 582236 3266
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667936 3478 667992
rect 3054 653520 3110 653576
rect 3238 624824 3294 624880
rect 3330 595992 3386 596048
rect 3146 481072 3202 481128
rect 3054 452376 3110 452432
rect 3330 423700 3386 423736
rect 3330 423680 3332 423700
rect 3332 423680 3384 423700
rect 3384 423680 3386 423700
rect 3514 610408 3570 610464
rect 3146 394984 3202 395040
rect 4066 567296 4122 567352
rect 3606 553016 3662 553072
rect 3422 380568 3478 380624
rect 3054 337456 3110 337512
rect 3514 366152 3570 366208
rect 3422 294344 3478 294400
rect 4066 538600 4122 538656
rect 8114 531256 8170 531312
rect 8390 531256 8446 531312
rect 8114 511944 8170 512000
rect 8390 511944 8446 512000
rect 3882 509904 3938 509960
rect 3698 495488 3754 495544
rect 7930 482976 7986 483032
rect 8206 482976 8262 483032
rect 3790 437960 3846 438016
rect 3606 323040 3662 323096
rect 3514 280064 3570 280120
rect 3422 251232 3478 251288
rect 3698 308760 3754 308816
rect 72974 608504 73030 608560
rect 73158 608504 73214 608560
rect 72698 531256 72754 531312
rect 72882 531256 72938 531312
rect 72606 511944 72662 512000
rect 72790 511944 72846 512000
rect 137834 531256 137890 531312
rect 138110 531256 138166 531312
rect 137834 511944 137890 512000
rect 138110 511944 138166 512000
rect 137650 482976 137706 483032
rect 137926 482976 137982 483032
rect 154210 482976 154266 483032
rect 154486 482976 154542 483032
rect 137466 463664 137522 463720
rect 137650 463664 137706 463720
rect 218150 560224 218206 560280
rect 218334 560224 218390 560280
rect 234710 560224 234766 560280
rect 234894 560224 234950 560280
rect 218150 540912 218206 540968
rect 218334 540912 218390 540968
rect 234710 540912 234766 540968
rect 234894 540912 234950 540968
rect 218150 521600 218206 521656
rect 218334 521600 218390 521656
rect 234710 521600 234766 521656
rect 234894 521600 234950 521656
rect 217966 502288 218022 502344
rect 218242 502324 218244 502344
rect 218244 502324 218296 502344
rect 218296 502324 218298 502344
rect 218242 502288 218298 502324
rect 234526 502288 234582 502344
rect 234802 502324 234804 502344
rect 234804 502324 234856 502344
rect 234856 502324 234858 502344
rect 234802 502288 234858 502324
rect 217966 492632 218022 492688
rect 218150 492632 218206 492688
rect 234526 492632 234582 492688
rect 234710 492632 234766 492688
rect 282918 683168 282974 683224
rect 283286 683168 283342 683224
rect 299662 569880 299718 569936
rect 299570 560360 299626 560416
rect 299570 560224 299626 560280
rect 299754 560224 299810 560280
rect 283102 521600 283158 521656
rect 283286 521600 283342 521656
rect 299662 521600 299718 521656
rect 299846 521600 299902 521656
rect 282918 502288 282974 502344
rect 283194 502324 283196 502344
rect 283196 502324 283248 502344
rect 283248 502324 283250 502344
rect 283194 502288 283250 502324
rect 299478 502288 299534 502344
rect 299754 502324 299756 502344
rect 299756 502324 299808 502344
rect 299808 502324 299810 502344
rect 299754 502288 299810 502324
rect 282918 492632 282974 492688
rect 283102 492652 283158 492688
rect 283102 492632 283104 492652
rect 283104 492632 283156 492652
rect 283156 492632 283158 492652
rect 299478 492632 299534 492688
rect 299662 492652 299718 492688
rect 299662 492632 299664 492652
rect 299664 492632 299716 492652
rect 299716 492632 299718 492652
rect 282918 454008 282974 454064
rect 283194 454008 283250 454064
rect 347870 560224 347926 560280
rect 348054 560224 348110 560280
rect 364430 560224 364486 560280
rect 364614 560224 364670 560280
rect 347870 540912 347926 540968
rect 348054 540912 348110 540968
rect 364430 540912 364486 540968
rect 364614 540912 364670 540968
rect 347870 521600 347926 521656
rect 348054 521600 348110 521656
rect 364430 521600 364486 521656
rect 364614 521600 364670 521656
rect 347962 502324 347964 502344
rect 347964 502324 348016 502344
rect 348016 502324 348018 502344
rect 347962 502288 348018 502324
rect 364246 502288 364302 502344
rect 364522 502324 364524 502344
rect 364524 502324 364576 502344
rect 364576 502324 364578 502344
rect 364522 502288 364578 502324
rect 347870 492632 347926 492688
rect 364246 492632 364302 492688
rect 364430 492632 364486 492688
rect 412822 521600 412878 521656
rect 413006 521600 413062 521656
rect 429382 521600 429438 521656
rect 429566 521600 429622 521656
rect 412638 502288 412694 502344
rect 412914 502324 412916 502344
rect 412916 502324 412968 502344
rect 412968 502324 412970 502344
rect 412914 502288 412970 502324
rect 429198 502288 429254 502344
rect 429474 502324 429476 502344
rect 429476 502324 429528 502344
rect 429528 502324 429530 502344
rect 429474 502288 429530 502324
rect 412638 492632 412694 492688
rect 412822 492652 412878 492688
rect 412822 492632 412824 492652
rect 412824 492632 412876 492652
rect 412876 492632 412878 492652
rect 429198 492632 429254 492688
rect 429382 492652 429438 492688
rect 429382 492632 429384 492652
rect 429384 492632 429436 492652
rect 429436 492632 429438 492652
rect 412638 454008 412694 454064
rect 412914 454008 412970 454064
rect 429198 454008 429254 454064
rect 429474 454008 429530 454064
rect 477590 560224 477646 560280
rect 477774 560224 477830 560280
rect 494150 560224 494206 560280
rect 494334 560224 494390 560280
rect 477590 540912 477646 540968
rect 477774 540912 477830 540968
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 477590 521600 477646 521656
rect 477774 521600 477830 521656
rect 494150 521600 494206 521656
rect 494334 521600 494390 521656
rect 477406 502288 477462 502344
rect 477682 502324 477684 502344
rect 477684 502324 477736 502344
rect 477736 502324 477738 502344
rect 477682 502288 477738 502324
rect 493966 502288 494022 502344
rect 494242 502324 494244 502344
rect 494244 502324 494296 502344
rect 494296 502324 494298 502344
rect 494242 502288 494298 502324
rect 477406 492632 477462 492688
rect 477590 492632 477646 492688
rect 493966 492632 494022 492688
rect 494150 492632 494206 492688
rect 580170 697992 580226 698048
rect 542358 683168 542414 683224
rect 542726 683168 542782 683224
rect 542542 521600 542598 521656
rect 542726 521600 542782 521656
rect 542358 502288 542414 502344
rect 542634 502324 542636 502344
rect 542636 502324 542688 502344
rect 542688 502324 542690 502344
rect 542634 502288 542690 502324
rect 542358 492632 542414 492688
rect 542542 492652 542598 492688
rect 542542 492632 542544 492652
rect 542544 492632 542596 492652
rect 542596 492632 542598 492652
rect 542358 454008 542414 454064
rect 542634 454008 542690 454064
rect 401598 418784 401654 418840
rect 78678 418512 78734 418568
rect 401598 411712 401654 411768
rect 78678 410896 78734 410952
rect 401598 404504 401654 404560
rect 78678 403280 78734 403336
rect 401598 397432 401654 397488
rect 78678 395664 78734 395720
rect 401598 390360 401654 390416
rect 78678 388048 78734 388104
rect 401598 383152 401654 383208
rect 78678 380432 78734 380488
rect 401598 376080 401654 376136
rect 78678 372816 78734 372872
rect 401598 369008 401654 369064
rect 78678 365200 78734 365256
rect 401598 361800 401654 361856
rect 78678 357584 78734 357640
rect 401598 354728 401654 354784
rect 78678 349968 78734 350024
rect 401598 347692 401600 347712
rect 401600 347692 401652 347712
rect 401652 347692 401654 347712
rect 401598 347656 401654 347692
rect 78678 342216 78734 342272
rect 401598 340448 401654 340504
rect 78678 334600 78734 334656
rect 401598 333376 401654 333432
rect 78678 327020 78680 327040
rect 78680 327020 78732 327040
rect 78732 327020 78734 327040
rect 78678 326984 78734 327020
rect 401598 326304 401654 326360
rect 78678 319368 78734 319424
rect 401598 319096 401654 319152
rect 401598 312024 401654 312080
rect 78678 311788 78680 311808
rect 78680 311788 78732 311808
rect 78732 311788 78734 311808
rect 78678 311752 78734 311788
rect 401598 304816 401654 304872
rect 78678 304136 78734 304192
rect 401598 297744 401654 297800
rect 78678 296520 78734 296576
rect 401598 290672 401654 290728
rect 78678 288904 78734 288960
rect 401598 283464 401654 283520
rect 78678 281288 78734 281344
rect 401598 276392 401654 276448
rect 78678 273672 78734 273728
rect 401598 269320 401654 269376
rect 78678 266056 78734 266112
rect 3606 265648 3662 265704
rect 401598 262148 401600 262168
rect 401600 262148 401652 262168
rect 401652 262148 401654 262168
rect 401598 262112 401654 262148
rect 78678 258304 78734 258360
rect 401598 255076 401600 255096
rect 401600 255076 401652 255096
rect 401652 255076 401654 255096
rect 401598 255040 401654 255076
rect 78678 250688 78734 250744
rect 402242 247968 402298 248024
rect 78678 243072 78734 243128
rect 401598 240760 401654 240816
rect 3514 236952 3570 237008
rect 78678 235456 78734 235512
rect 401598 233688 401654 233744
rect 78678 227840 78734 227896
rect 401598 226616 401654 226672
rect 2962 222536 3018 222592
rect 78678 220224 78734 220280
rect 401598 219408 401654 219464
rect 79322 212608 79378 212664
rect 401598 212372 401600 212392
rect 401600 212372 401652 212392
rect 401652 212372 401654 212392
rect 401598 212336 401654 212372
rect 3422 208120 3478 208176
rect 559102 521600 559158 521656
rect 559286 521600 559342 521656
rect 558918 502288 558974 502344
rect 559194 502324 559196 502344
rect 559196 502324 559248 502344
rect 559248 502324 559250 502344
rect 559194 502288 559250 502324
rect 558918 492632 558974 492688
rect 559102 492652 559158 492688
rect 559102 492632 559104 492652
rect 559104 492632 559156 492652
rect 559156 492632 559158 492652
rect 558918 454008 558974 454064
rect 559194 454008 559250 454064
rect 580262 686296 580318 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 580170 545536 580226 545592
rect 578882 533840 578938 533896
rect 580170 510312 580226 510368
rect 580170 498616 580226 498672
rect 579894 486784 579950 486840
rect 580170 463392 580226 463448
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 580354 451696 580410 451752
rect 580262 404776 580318 404832
rect 580170 392944 580226 393000
rect 580170 369552 580226 369608
rect 579894 357856 579950 357912
rect 580170 346024 580226 346080
rect 578882 322632 578938 322688
rect 579618 310800 579674 310856
rect 578882 299104 578938 299160
rect 580170 275712 580226 275768
rect 579802 263880 579858 263936
rect 580170 252184 580226 252240
rect 580170 228792 580226 228848
rect 580262 216960 580318 217016
rect 401598 205128 401654 205184
rect 79322 204992 79378 205048
rect 580354 205264 580410 205320
rect 401598 198056 401654 198112
rect 79414 197376 79470 197432
rect 3146 193840 3202 193896
rect 79322 189760 79378 189816
rect 3238 179424 3294 179480
rect 78678 166776 78734 166832
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 401598 190984 401654 191040
rect 401598 183776 401654 183832
rect 79506 182008 79562 182064
rect 79414 174392 79470 174448
rect 79322 159160 79378 159216
rect 78678 143928 78734 143984
rect 78678 121080 78734 121136
rect 3514 78920 3570 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 580170 181872 580226 181928
rect 402242 176704 402298 176760
rect 580170 170040 580226 170096
rect 402242 169632 402298 169688
rect 402334 162424 402390 162480
rect 402242 155352 402298 155408
rect 79690 151544 79746 151600
rect 79598 136312 79654 136368
rect 79506 128696 79562 128752
rect 79414 113464 79470 113520
rect 79322 105848 79378 105904
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 401598 126928 401654 126984
rect 579802 158344 579858 158400
rect 402610 148280 402666 148336
rect 402518 141072 402574 141128
rect 402426 134000 402482 134056
rect 402334 119720 402390 119776
rect 402242 112648 402298 112704
rect 401598 105576 401654 105632
rect 3422 7112 3478 7168
rect 91926 85448 91982 85504
rect 92202 85448 92258 85504
rect 96250 96600 96306 96656
rect 96434 96600 96490 96656
rect 96342 80688 96398 80744
rect 96342 67632 96398 67688
rect 104530 96600 104586 96656
rect 104714 96600 104770 96656
rect 151450 96600 151506 96656
rect 151634 96600 151690 96656
rect 151634 80144 151690 80200
rect 151542 77288 151598 77344
rect 197726 67496 197782 67552
rect 198002 67496 198058 67552
rect 198554 29008 198610 29064
rect 198738 29008 198794 29064
rect 215022 64912 215078 64968
rect 215206 64912 215262 64968
rect 215022 60696 215078 60752
rect 215022 48320 215078 48376
rect 227074 77288 227130 77344
rect 227258 77288 227314 77344
rect 227258 67768 227314 67824
rect 227258 67632 227314 67688
rect 227442 61376 227498 61432
rect 227350 48320 227406 48376
rect 239770 96600 239826 96656
rect 239954 96600 240010 96656
rect 274362 96600 274418 96656
rect 274546 96600 274602 96656
rect 341706 77288 341762 77344
rect 341890 77288 341946 77344
rect 341890 67768 341946 67824
rect 341890 67632 341946 67688
rect 370686 86944 370742 87000
rect 370870 86944 370926 87000
rect 580170 134816 580226 134872
rect 550638 77152 550694 77208
rect 550914 77152 550970 77208
rect 550638 58112 550694 58168
rect 550638 57976 550694 58032
rect 568578 48456 568634 48512
rect 568578 48320 568634 48376
rect 568026 8200 568082 8256
rect 568210 8064 568266 8120
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 578882 64504 578938 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 282913 683226 282979 683229
rect 283281 683226 283347 683229
rect 282913 683224 283347 683226
rect 282913 683168 282918 683224
rect 282974 683168 283286 683224
rect 283342 683168 283347 683224
rect 282913 683166 283347 683168
rect 282913 683163 282979 683166
rect 283281 683163 283347 683166
rect 542353 683226 542419 683229
rect 542721 683226 542787 683229
rect 542353 683224 542787 683226
rect 542353 683168 542358 683224
rect 542414 683168 542726 683224
rect 542782 683168 542787 683224
rect 542353 683166 542787 683168
rect 542353 683163 542419 683166
rect 542721 683163 542787 683166
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3233 624882 3299 624885
rect -960 624880 3299 624882
rect -960 624824 3238 624880
rect 3294 624824 3299 624880
rect -960 624822 3299 624824
rect -960 624732 480 624822
rect 3233 624819 3299 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3509 610466 3575 610469
rect -960 610464 3575 610466
rect -960 610408 3514 610464
rect 3570 610408 3575 610464
rect -960 610406 3575 610408
rect -960 610316 480 610406
rect 3509 610403 3575 610406
rect 72969 608562 73035 608565
rect 73153 608562 73219 608565
rect 72969 608560 73219 608562
rect 72969 608504 72974 608560
rect 73030 608504 73158 608560
rect 73214 608504 73219 608560
rect 72969 608502 73219 608504
rect 72969 608499 73035 608502
rect 73153 608499 73219 608502
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 299657 569940 299723 569941
rect 299606 569938 299612 569940
rect 299566 569878 299612 569938
rect 299676 569936 299723 569940
rect 299718 569880 299723 569936
rect 299606 569876 299612 569878
rect 299676 569876 299723 569880
rect 299657 569875 299723 569876
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 299565 560420 299631 560421
rect 299565 560418 299612 560420
rect 299520 560416 299612 560418
rect 299520 560360 299570 560416
rect 299520 560358 299612 560360
rect 299565 560356 299612 560358
rect 299676 560356 299682 560420
rect 299565 560355 299631 560356
rect 218145 560282 218211 560285
rect 218329 560282 218395 560285
rect 218145 560280 218395 560282
rect 218145 560224 218150 560280
rect 218206 560224 218334 560280
rect 218390 560224 218395 560280
rect 218145 560222 218395 560224
rect 218145 560219 218211 560222
rect 218329 560219 218395 560222
rect 234705 560282 234771 560285
rect 234889 560282 234955 560285
rect 234705 560280 234955 560282
rect 234705 560224 234710 560280
rect 234766 560224 234894 560280
rect 234950 560224 234955 560280
rect 234705 560222 234955 560224
rect 234705 560219 234771 560222
rect 234889 560219 234955 560222
rect 299565 560282 299631 560285
rect 299749 560282 299815 560285
rect 299565 560280 299815 560282
rect 299565 560224 299570 560280
rect 299626 560224 299754 560280
rect 299810 560224 299815 560280
rect 299565 560222 299815 560224
rect 299565 560219 299631 560222
rect 299749 560219 299815 560222
rect 347865 560282 347931 560285
rect 348049 560282 348115 560285
rect 347865 560280 348115 560282
rect 347865 560224 347870 560280
rect 347926 560224 348054 560280
rect 348110 560224 348115 560280
rect 347865 560222 348115 560224
rect 347865 560219 347931 560222
rect 348049 560219 348115 560222
rect 364425 560282 364491 560285
rect 364609 560282 364675 560285
rect 364425 560280 364675 560282
rect 364425 560224 364430 560280
rect 364486 560224 364614 560280
rect 364670 560224 364675 560280
rect 364425 560222 364675 560224
rect 364425 560219 364491 560222
rect 364609 560219 364675 560222
rect 477585 560282 477651 560285
rect 477769 560282 477835 560285
rect 477585 560280 477835 560282
rect 477585 560224 477590 560280
rect 477646 560224 477774 560280
rect 477830 560224 477835 560280
rect 477585 560222 477835 560224
rect 477585 560219 477651 560222
rect 477769 560219 477835 560222
rect 494145 560282 494211 560285
rect 494329 560282 494395 560285
rect 494145 560280 494395 560282
rect 494145 560224 494150 560280
rect 494206 560224 494334 560280
rect 494390 560224 494395 560280
rect 494145 560222 494395 560224
rect 494145 560219 494211 560222
rect 494329 560219 494395 560222
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3601 553074 3667 553077
rect -960 553072 3667 553074
rect -960 553016 3606 553072
rect 3662 553016 3667 553072
rect -960 553014 3667 553016
rect -960 552924 480 553014
rect 3601 553011 3667 553014
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218145 540970 218211 540973
rect 218329 540970 218395 540973
rect 218145 540968 218395 540970
rect 218145 540912 218150 540968
rect 218206 540912 218334 540968
rect 218390 540912 218395 540968
rect 218145 540910 218395 540912
rect 218145 540907 218211 540910
rect 218329 540907 218395 540910
rect 234705 540970 234771 540973
rect 234889 540970 234955 540973
rect 234705 540968 234955 540970
rect 234705 540912 234710 540968
rect 234766 540912 234894 540968
rect 234950 540912 234955 540968
rect 234705 540910 234955 540912
rect 234705 540907 234771 540910
rect 234889 540907 234955 540910
rect 347865 540970 347931 540973
rect 348049 540970 348115 540973
rect 347865 540968 348115 540970
rect 347865 540912 347870 540968
rect 347926 540912 348054 540968
rect 348110 540912 348115 540968
rect 347865 540910 348115 540912
rect 347865 540907 347931 540910
rect 348049 540907 348115 540910
rect 364425 540970 364491 540973
rect 364609 540970 364675 540973
rect 364425 540968 364675 540970
rect 364425 540912 364430 540968
rect 364486 540912 364614 540968
rect 364670 540912 364675 540968
rect 364425 540910 364675 540912
rect 364425 540907 364491 540910
rect 364609 540907 364675 540910
rect 477585 540970 477651 540973
rect 477769 540970 477835 540973
rect 477585 540968 477835 540970
rect 477585 540912 477590 540968
rect 477646 540912 477774 540968
rect 477830 540912 477835 540968
rect 477585 540910 477835 540912
rect 477585 540907 477651 540910
rect 477769 540907 477835 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -960 538658 480 538748
rect 4061 538658 4127 538661
rect -960 538656 4127 538658
rect -960 538600 4066 538656
rect 4122 538600 4127 538656
rect -960 538598 4127 538600
rect -960 538508 480 538598
rect 4061 538595 4127 538598
rect 578877 533898 578943 533901
rect 583520 533898 584960 533988
rect 578877 533896 584960 533898
rect 578877 533840 578882 533896
rect 578938 533840 584960 533896
rect 578877 533838 584960 533840
rect 578877 533835 578943 533838
rect 583520 533748 584960 533838
rect 8109 531314 8175 531317
rect 8385 531314 8451 531317
rect 8109 531312 8451 531314
rect 8109 531256 8114 531312
rect 8170 531256 8390 531312
rect 8446 531256 8451 531312
rect 8109 531254 8451 531256
rect 8109 531251 8175 531254
rect 8385 531251 8451 531254
rect 72693 531314 72759 531317
rect 72877 531314 72943 531317
rect 72693 531312 72943 531314
rect 72693 531256 72698 531312
rect 72754 531256 72882 531312
rect 72938 531256 72943 531312
rect 72693 531254 72943 531256
rect 72693 531251 72759 531254
rect 72877 531251 72943 531254
rect 137829 531314 137895 531317
rect 138105 531314 138171 531317
rect 137829 531312 138171 531314
rect 137829 531256 137834 531312
rect 137890 531256 138110 531312
rect 138166 531256 138171 531312
rect 137829 531254 138171 531256
rect 137829 531251 137895 531254
rect 138105 531251 138171 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 218145 521658 218211 521661
rect 218329 521658 218395 521661
rect 218145 521656 218395 521658
rect 218145 521600 218150 521656
rect 218206 521600 218334 521656
rect 218390 521600 218395 521656
rect 218145 521598 218395 521600
rect 218145 521595 218211 521598
rect 218329 521595 218395 521598
rect 234705 521658 234771 521661
rect 234889 521658 234955 521661
rect 234705 521656 234955 521658
rect 234705 521600 234710 521656
rect 234766 521600 234894 521656
rect 234950 521600 234955 521656
rect 234705 521598 234955 521600
rect 234705 521595 234771 521598
rect 234889 521595 234955 521598
rect 283097 521658 283163 521661
rect 283281 521658 283347 521661
rect 283097 521656 283347 521658
rect 283097 521600 283102 521656
rect 283158 521600 283286 521656
rect 283342 521600 283347 521656
rect 283097 521598 283347 521600
rect 283097 521595 283163 521598
rect 283281 521595 283347 521598
rect 299657 521658 299723 521661
rect 299841 521658 299907 521661
rect 299657 521656 299907 521658
rect 299657 521600 299662 521656
rect 299718 521600 299846 521656
rect 299902 521600 299907 521656
rect 299657 521598 299907 521600
rect 299657 521595 299723 521598
rect 299841 521595 299907 521598
rect 347865 521658 347931 521661
rect 348049 521658 348115 521661
rect 347865 521656 348115 521658
rect 347865 521600 347870 521656
rect 347926 521600 348054 521656
rect 348110 521600 348115 521656
rect 347865 521598 348115 521600
rect 347865 521595 347931 521598
rect 348049 521595 348115 521598
rect 364425 521658 364491 521661
rect 364609 521658 364675 521661
rect 364425 521656 364675 521658
rect 364425 521600 364430 521656
rect 364486 521600 364614 521656
rect 364670 521600 364675 521656
rect 364425 521598 364675 521600
rect 364425 521595 364491 521598
rect 364609 521595 364675 521598
rect 412817 521658 412883 521661
rect 413001 521658 413067 521661
rect 412817 521656 413067 521658
rect 412817 521600 412822 521656
rect 412878 521600 413006 521656
rect 413062 521600 413067 521656
rect 412817 521598 413067 521600
rect 412817 521595 412883 521598
rect 413001 521595 413067 521598
rect 429377 521658 429443 521661
rect 429561 521658 429627 521661
rect 429377 521656 429627 521658
rect 429377 521600 429382 521656
rect 429438 521600 429566 521656
rect 429622 521600 429627 521656
rect 429377 521598 429627 521600
rect 429377 521595 429443 521598
rect 429561 521595 429627 521598
rect 477585 521658 477651 521661
rect 477769 521658 477835 521661
rect 477585 521656 477835 521658
rect 477585 521600 477590 521656
rect 477646 521600 477774 521656
rect 477830 521600 477835 521656
rect 477585 521598 477835 521600
rect 477585 521595 477651 521598
rect 477769 521595 477835 521598
rect 494145 521658 494211 521661
rect 494329 521658 494395 521661
rect 494145 521656 494395 521658
rect 494145 521600 494150 521656
rect 494206 521600 494334 521656
rect 494390 521600 494395 521656
rect 494145 521598 494395 521600
rect 494145 521595 494211 521598
rect 494329 521595 494395 521598
rect 542537 521658 542603 521661
rect 542721 521658 542787 521661
rect 542537 521656 542787 521658
rect 542537 521600 542542 521656
rect 542598 521600 542726 521656
rect 542782 521600 542787 521656
rect 542537 521598 542787 521600
rect 542537 521595 542603 521598
rect 542721 521595 542787 521598
rect 559097 521658 559163 521661
rect 559281 521658 559347 521661
rect 559097 521656 559347 521658
rect 559097 521600 559102 521656
rect 559158 521600 559286 521656
rect 559342 521600 559347 521656
rect 559097 521598 559347 521600
rect 559097 521595 559163 521598
rect 559281 521595 559347 521598
rect 8109 512002 8175 512005
rect 8385 512002 8451 512005
rect 8109 512000 8451 512002
rect 8109 511944 8114 512000
rect 8170 511944 8390 512000
rect 8446 511944 8451 512000
rect 8109 511942 8451 511944
rect 8109 511939 8175 511942
rect 8385 511939 8451 511942
rect 72601 512002 72667 512005
rect 72785 512002 72851 512005
rect 72601 512000 72851 512002
rect 72601 511944 72606 512000
rect 72662 511944 72790 512000
rect 72846 511944 72851 512000
rect 72601 511942 72851 511944
rect 72601 511939 72667 511942
rect 72785 511939 72851 511942
rect 137829 512002 137895 512005
rect 138105 512002 138171 512005
rect 137829 512000 138171 512002
rect 137829 511944 137834 512000
rect 137890 511944 138110 512000
rect 138166 511944 138171 512000
rect 137829 511942 138171 511944
rect 137829 511939 137895 511942
rect 138105 511939 138171 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3877 509962 3943 509965
rect -960 509960 3943 509962
rect -960 509904 3882 509960
rect 3938 509904 3943 509960
rect -960 509902 3943 509904
rect -960 509812 480 509902
rect 3877 509899 3943 509902
rect 217961 502346 218027 502349
rect 218237 502346 218303 502349
rect 217961 502344 218303 502346
rect 217961 502288 217966 502344
rect 218022 502288 218242 502344
rect 218298 502288 218303 502344
rect 217961 502286 218303 502288
rect 217961 502283 218027 502286
rect 218237 502283 218303 502286
rect 234521 502346 234587 502349
rect 234797 502346 234863 502349
rect 234521 502344 234863 502346
rect 234521 502288 234526 502344
rect 234582 502288 234802 502344
rect 234858 502288 234863 502344
rect 234521 502286 234863 502288
rect 234521 502283 234587 502286
rect 234797 502283 234863 502286
rect 282913 502346 282979 502349
rect 283189 502346 283255 502349
rect 282913 502344 283255 502346
rect 282913 502288 282918 502344
rect 282974 502288 283194 502344
rect 283250 502288 283255 502344
rect 282913 502286 283255 502288
rect 282913 502283 282979 502286
rect 283189 502283 283255 502286
rect 299473 502346 299539 502349
rect 299749 502346 299815 502349
rect 299473 502344 299815 502346
rect 299473 502288 299478 502344
rect 299534 502288 299754 502344
rect 299810 502288 299815 502344
rect 299473 502286 299815 502288
rect 299473 502283 299539 502286
rect 299749 502283 299815 502286
rect 347814 502284 347820 502348
rect 347884 502346 347890 502348
rect 347957 502346 348023 502349
rect 347884 502344 348023 502346
rect 347884 502288 347962 502344
rect 348018 502288 348023 502344
rect 347884 502286 348023 502288
rect 347884 502284 347890 502286
rect 347957 502283 348023 502286
rect 364241 502346 364307 502349
rect 364517 502346 364583 502349
rect 364241 502344 364583 502346
rect 364241 502288 364246 502344
rect 364302 502288 364522 502344
rect 364578 502288 364583 502344
rect 364241 502286 364583 502288
rect 364241 502283 364307 502286
rect 364517 502283 364583 502286
rect 412633 502346 412699 502349
rect 412909 502346 412975 502349
rect 412633 502344 412975 502346
rect 412633 502288 412638 502344
rect 412694 502288 412914 502344
rect 412970 502288 412975 502344
rect 412633 502286 412975 502288
rect 412633 502283 412699 502286
rect 412909 502283 412975 502286
rect 429193 502346 429259 502349
rect 429469 502346 429535 502349
rect 429193 502344 429535 502346
rect 429193 502288 429198 502344
rect 429254 502288 429474 502344
rect 429530 502288 429535 502344
rect 429193 502286 429535 502288
rect 429193 502283 429259 502286
rect 429469 502283 429535 502286
rect 477401 502346 477467 502349
rect 477677 502346 477743 502349
rect 477401 502344 477743 502346
rect 477401 502288 477406 502344
rect 477462 502288 477682 502344
rect 477738 502288 477743 502344
rect 477401 502286 477743 502288
rect 477401 502283 477467 502286
rect 477677 502283 477743 502286
rect 493961 502346 494027 502349
rect 494237 502346 494303 502349
rect 493961 502344 494303 502346
rect 493961 502288 493966 502344
rect 494022 502288 494242 502344
rect 494298 502288 494303 502344
rect 493961 502286 494303 502288
rect 493961 502283 494027 502286
rect 494237 502283 494303 502286
rect 542353 502346 542419 502349
rect 542629 502346 542695 502349
rect 542353 502344 542695 502346
rect 542353 502288 542358 502344
rect 542414 502288 542634 502344
rect 542690 502288 542695 502344
rect 542353 502286 542695 502288
rect 542353 502283 542419 502286
rect 542629 502283 542695 502286
rect 558913 502346 558979 502349
rect 559189 502346 559255 502349
rect 558913 502344 559255 502346
rect 558913 502288 558918 502344
rect 558974 502288 559194 502344
rect 559250 502288 559255 502344
rect 558913 502286 559255 502288
rect 558913 502283 558979 502286
rect 559189 502283 559255 502286
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3693 495546 3759 495549
rect -960 495544 3759 495546
rect -960 495488 3698 495544
rect 3754 495488 3759 495544
rect -960 495486 3759 495488
rect -960 495396 480 495486
rect 3693 495483 3759 495486
rect 217961 492690 218027 492693
rect 218145 492690 218211 492693
rect 217961 492688 218211 492690
rect 217961 492632 217966 492688
rect 218022 492632 218150 492688
rect 218206 492632 218211 492688
rect 217961 492630 218211 492632
rect 217961 492627 218027 492630
rect 218145 492627 218211 492630
rect 234521 492690 234587 492693
rect 234705 492690 234771 492693
rect 234521 492688 234771 492690
rect 234521 492632 234526 492688
rect 234582 492632 234710 492688
rect 234766 492632 234771 492688
rect 234521 492630 234771 492632
rect 234521 492627 234587 492630
rect 234705 492627 234771 492630
rect 282913 492690 282979 492693
rect 283097 492690 283163 492693
rect 282913 492688 283163 492690
rect 282913 492632 282918 492688
rect 282974 492632 283102 492688
rect 283158 492632 283163 492688
rect 282913 492630 283163 492632
rect 282913 492627 282979 492630
rect 283097 492627 283163 492630
rect 299473 492690 299539 492693
rect 299657 492690 299723 492693
rect 347865 492692 347931 492693
rect 299473 492688 299723 492690
rect 299473 492632 299478 492688
rect 299534 492632 299662 492688
rect 299718 492632 299723 492688
rect 299473 492630 299723 492632
rect 299473 492627 299539 492630
rect 299657 492627 299723 492630
rect 347814 492628 347820 492692
rect 347884 492690 347931 492692
rect 364241 492690 364307 492693
rect 364425 492690 364491 492693
rect 347884 492688 347976 492690
rect 347926 492632 347976 492688
rect 347884 492630 347976 492632
rect 364241 492688 364491 492690
rect 364241 492632 364246 492688
rect 364302 492632 364430 492688
rect 364486 492632 364491 492688
rect 364241 492630 364491 492632
rect 347884 492628 347931 492630
rect 347865 492627 347931 492628
rect 364241 492627 364307 492630
rect 364425 492627 364491 492630
rect 412633 492690 412699 492693
rect 412817 492690 412883 492693
rect 412633 492688 412883 492690
rect 412633 492632 412638 492688
rect 412694 492632 412822 492688
rect 412878 492632 412883 492688
rect 412633 492630 412883 492632
rect 412633 492627 412699 492630
rect 412817 492627 412883 492630
rect 429193 492690 429259 492693
rect 429377 492690 429443 492693
rect 429193 492688 429443 492690
rect 429193 492632 429198 492688
rect 429254 492632 429382 492688
rect 429438 492632 429443 492688
rect 429193 492630 429443 492632
rect 429193 492627 429259 492630
rect 429377 492627 429443 492630
rect 477401 492690 477467 492693
rect 477585 492690 477651 492693
rect 477401 492688 477651 492690
rect 477401 492632 477406 492688
rect 477462 492632 477590 492688
rect 477646 492632 477651 492688
rect 477401 492630 477651 492632
rect 477401 492627 477467 492630
rect 477585 492627 477651 492630
rect 493961 492690 494027 492693
rect 494145 492690 494211 492693
rect 493961 492688 494211 492690
rect 493961 492632 493966 492688
rect 494022 492632 494150 492688
rect 494206 492632 494211 492688
rect 493961 492630 494211 492632
rect 493961 492627 494027 492630
rect 494145 492627 494211 492630
rect 542353 492690 542419 492693
rect 542537 492690 542603 492693
rect 542353 492688 542603 492690
rect 542353 492632 542358 492688
rect 542414 492632 542542 492688
rect 542598 492632 542603 492688
rect 542353 492630 542603 492632
rect 542353 492627 542419 492630
rect 542537 492627 542603 492630
rect 558913 492690 558979 492693
rect 559097 492690 559163 492693
rect 558913 492688 559163 492690
rect 558913 492632 558918 492688
rect 558974 492632 559102 492688
rect 559158 492632 559163 492688
rect 558913 492630 559163 492632
rect 558913 492627 558979 492630
rect 559097 492627 559163 492630
rect 579889 486842 579955 486845
rect 583520 486842 584960 486932
rect 579889 486840 584960 486842
rect 579889 486784 579894 486840
rect 579950 486784 584960 486840
rect 579889 486782 584960 486784
rect 579889 486779 579955 486782
rect 583520 486692 584960 486782
rect 7925 483034 7991 483037
rect 8201 483034 8267 483037
rect 7925 483032 8267 483034
rect 7925 482976 7930 483032
rect 7986 482976 8206 483032
rect 8262 482976 8267 483032
rect 7925 482974 8267 482976
rect 7925 482971 7991 482974
rect 8201 482971 8267 482974
rect 137645 483034 137711 483037
rect 137921 483034 137987 483037
rect 137645 483032 137987 483034
rect 137645 482976 137650 483032
rect 137706 482976 137926 483032
rect 137982 482976 137987 483032
rect 137645 482974 137987 482976
rect 137645 482971 137711 482974
rect 137921 482971 137987 482974
rect 154205 483034 154271 483037
rect 154481 483034 154547 483037
rect 154205 483032 154547 483034
rect 154205 482976 154210 483032
rect 154266 482976 154486 483032
rect 154542 482976 154547 483032
rect 154205 482974 154547 482976
rect 154205 482971 154271 482974
rect 154481 482971 154547 482974
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 137461 463722 137527 463725
rect 137645 463722 137711 463725
rect 137461 463720 137711 463722
rect 137461 463664 137466 463720
rect 137522 463664 137650 463720
rect 137706 463664 137711 463720
rect 137461 463662 137711 463664
rect 137461 463659 137527 463662
rect 137645 463659 137711 463662
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 282913 454066 282979 454069
rect 283189 454066 283255 454069
rect 282913 454064 283255 454066
rect 282913 454008 282918 454064
rect 282974 454008 283194 454064
rect 283250 454008 283255 454064
rect 282913 454006 283255 454008
rect 282913 454003 282979 454006
rect 283189 454003 283255 454006
rect 412633 454066 412699 454069
rect 412909 454066 412975 454069
rect 412633 454064 412975 454066
rect 412633 454008 412638 454064
rect 412694 454008 412914 454064
rect 412970 454008 412975 454064
rect 412633 454006 412975 454008
rect 412633 454003 412699 454006
rect 412909 454003 412975 454006
rect 429193 454066 429259 454069
rect 429469 454066 429535 454069
rect 429193 454064 429535 454066
rect 429193 454008 429198 454064
rect 429254 454008 429474 454064
rect 429530 454008 429535 454064
rect 429193 454006 429535 454008
rect 429193 454003 429259 454006
rect 429469 454003 429535 454006
rect 542353 454066 542419 454069
rect 542629 454066 542695 454069
rect 542353 454064 542695 454066
rect 542353 454008 542358 454064
rect 542414 454008 542634 454064
rect 542690 454008 542695 454064
rect 542353 454006 542695 454008
rect 542353 454003 542419 454006
rect 542629 454003 542695 454006
rect 558913 454066 558979 454069
rect 559189 454066 559255 454069
rect 558913 454064 559255 454066
rect 558913 454008 558918 454064
rect 558974 454008 559194 454064
rect 559250 454008 559255 454064
rect 558913 454006 559255 454008
rect 558913 454003 558979 454006
rect 559189 454003 559255 454006
rect -960 452434 480 452524
rect 3049 452434 3115 452437
rect -960 452432 3115 452434
rect -960 452376 3054 452432
rect 3110 452376 3115 452432
rect -960 452374 3115 452376
rect -960 452284 480 452374
rect 3049 452371 3115 452374
rect 580349 451754 580415 451757
rect 583520 451754 584960 451844
rect 580349 451752 584960 451754
rect 580349 451696 580354 451752
rect 580410 451696 584960 451752
rect 580349 451694 584960 451696
rect 580349 451691 580415 451694
rect 583520 451604 584960 451694
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3785 438018 3851 438021
rect -960 438016 3851 438018
rect -960 437960 3790 438016
rect 3846 437960 3851 438016
rect -960 437958 3851 437960
rect -960 437868 480 437958
rect 3785 437955 3851 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 401593 418842 401659 418845
rect 400292 418840 401659 418842
rect 400292 418784 401598 418840
rect 401654 418784 401659 418840
rect 400292 418782 401659 418784
rect 401593 418779 401659 418782
rect 78673 418570 78739 418573
rect 78673 418568 82156 418570
rect 78673 418512 78678 418568
rect 78734 418512 82156 418568
rect 78673 418510 82156 418512
rect 78673 418507 78739 418510
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 401593 411770 401659 411773
rect 400292 411768 401659 411770
rect 400292 411712 401598 411768
rect 401654 411712 401659 411768
rect 400292 411710 401659 411712
rect 401593 411707 401659 411710
rect 78673 410954 78739 410957
rect 78673 410952 82156 410954
rect 78673 410896 78678 410952
rect 78734 410896 82156 410952
rect 78673 410894 82156 410896
rect 78673 410891 78739 410894
rect -960 409172 480 409412
rect 580257 404834 580323 404837
rect 583520 404834 584960 404924
rect 580257 404832 584960 404834
rect 580257 404776 580262 404832
rect 580318 404776 584960 404832
rect 580257 404774 584960 404776
rect 580257 404771 580323 404774
rect 583520 404684 584960 404774
rect 401593 404562 401659 404565
rect 400292 404560 401659 404562
rect 400292 404504 401598 404560
rect 401654 404504 401659 404560
rect 400292 404502 401659 404504
rect 401593 404499 401659 404502
rect 78673 403338 78739 403341
rect 78673 403336 82156 403338
rect 78673 403280 78678 403336
rect 78734 403280 82156 403336
rect 78673 403278 82156 403280
rect 78673 403275 78739 403278
rect 401593 397490 401659 397493
rect 400292 397488 401659 397490
rect 400292 397432 401598 397488
rect 401654 397432 401659 397488
rect 400292 397430 401659 397432
rect 401593 397427 401659 397430
rect 78673 395722 78739 395725
rect 78673 395720 82156 395722
rect 78673 395664 78678 395720
rect 78734 395664 82156 395720
rect 78673 395662 82156 395664
rect 78673 395659 78739 395662
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 401593 390418 401659 390421
rect 400292 390416 401659 390418
rect 400292 390360 401598 390416
rect 401654 390360 401659 390416
rect 400292 390358 401659 390360
rect 401593 390355 401659 390358
rect 78673 388106 78739 388109
rect 78673 388104 82156 388106
rect 78673 388048 78678 388104
rect 78734 388048 82156 388104
rect 78673 388046 82156 388048
rect 78673 388043 78739 388046
rect 401593 383210 401659 383213
rect 400292 383208 401659 383210
rect 400292 383152 401598 383208
rect 401654 383152 401659 383208
rect 400292 383150 401659 383152
rect 401593 383147 401659 383150
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 78673 380490 78739 380493
rect 78673 380488 82156 380490
rect 78673 380432 78678 380488
rect 78734 380432 82156 380488
rect 78673 380430 82156 380432
rect 78673 380427 78739 380430
rect 401593 376138 401659 376141
rect 400292 376136 401659 376138
rect 400292 376080 401598 376136
rect 401654 376080 401659 376136
rect 400292 376078 401659 376080
rect 401593 376075 401659 376078
rect 78673 372874 78739 372877
rect 78673 372872 82156 372874
rect 78673 372816 78678 372872
rect 78734 372816 82156 372872
rect 78673 372814 82156 372816
rect 78673 372811 78739 372814
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect 401593 369066 401659 369069
rect 400292 369064 401659 369066
rect 400292 369008 401598 369064
rect 401654 369008 401659 369064
rect 400292 369006 401659 369008
rect 401593 369003 401659 369006
rect -960 366210 480 366300
rect 3509 366210 3575 366213
rect -960 366208 3575 366210
rect -960 366152 3514 366208
rect 3570 366152 3575 366208
rect -960 366150 3575 366152
rect -960 366060 480 366150
rect 3509 366147 3575 366150
rect 78673 365258 78739 365261
rect 78673 365256 82156 365258
rect 78673 365200 78678 365256
rect 78734 365200 82156 365256
rect 78673 365198 82156 365200
rect 78673 365195 78739 365198
rect 401593 361858 401659 361861
rect 400292 361856 401659 361858
rect 400292 361800 401598 361856
rect 401654 361800 401659 361856
rect 400292 361798 401659 361800
rect 401593 361795 401659 361798
rect 579889 357914 579955 357917
rect 583520 357914 584960 358004
rect 579889 357912 584960 357914
rect 579889 357856 579894 357912
rect 579950 357856 584960 357912
rect 579889 357854 584960 357856
rect 579889 357851 579955 357854
rect 583520 357764 584960 357854
rect 78673 357642 78739 357645
rect 78673 357640 82156 357642
rect 78673 357584 78678 357640
rect 78734 357584 82156 357640
rect 78673 357582 82156 357584
rect 78673 357579 78739 357582
rect 401593 354786 401659 354789
rect 400292 354784 401659 354786
rect 400292 354728 401598 354784
rect 401654 354728 401659 354784
rect 400292 354726 401659 354728
rect 401593 354723 401659 354726
rect -960 351780 480 352020
rect 78673 350026 78739 350029
rect 78673 350024 82156 350026
rect 78673 349968 78678 350024
rect 78734 349968 82156 350024
rect 78673 349966 82156 349968
rect 78673 349963 78739 349966
rect 401593 347714 401659 347717
rect 400292 347712 401659 347714
rect 400292 347656 401598 347712
rect 401654 347656 401659 347712
rect 400292 347654 401659 347656
rect 401593 347651 401659 347654
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 78673 342274 78739 342277
rect 78673 342272 82156 342274
rect 78673 342216 78678 342272
rect 78734 342216 82156 342272
rect 78673 342214 82156 342216
rect 78673 342211 78739 342214
rect 401593 340506 401659 340509
rect 400292 340504 401659 340506
rect 400292 340448 401598 340504
rect 401654 340448 401659 340504
rect 400292 340446 401659 340448
rect 401593 340443 401659 340446
rect -960 337514 480 337604
rect 3049 337514 3115 337517
rect -960 337512 3115 337514
rect -960 337456 3054 337512
rect 3110 337456 3115 337512
rect -960 337454 3115 337456
rect -960 337364 480 337454
rect 3049 337451 3115 337454
rect 78673 334658 78739 334661
rect 78673 334656 82156 334658
rect 78673 334600 78678 334656
rect 78734 334600 82156 334656
rect 78673 334598 82156 334600
rect 78673 334595 78739 334598
rect 583520 334236 584960 334476
rect 401593 333434 401659 333437
rect 400292 333432 401659 333434
rect 400292 333376 401598 333432
rect 401654 333376 401659 333432
rect 400292 333374 401659 333376
rect 401593 333371 401659 333374
rect 78673 327042 78739 327045
rect 78673 327040 82156 327042
rect 78673 326984 78678 327040
rect 78734 326984 82156 327040
rect 78673 326982 82156 326984
rect 78673 326979 78739 326982
rect 401593 326362 401659 326365
rect 400292 326360 401659 326362
rect 400292 326304 401598 326360
rect 401654 326304 401659 326360
rect 400292 326302 401659 326304
rect 401593 326299 401659 326302
rect -960 323098 480 323188
rect 3601 323098 3667 323101
rect -960 323096 3667 323098
rect -960 323040 3606 323096
rect 3662 323040 3667 323096
rect -960 323038 3667 323040
rect -960 322948 480 323038
rect 3601 323035 3667 323038
rect 578877 322690 578943 322693
rect 583520 322690 584960 322780
rect 578877 322688 584960 322690
rect 578877 322632 578882 322688
rect 578938 322632 584960 322688
rect 578877 322630 584960 322632
rect 578877 322627 578943 322630
rect 583520 322540 584960 322630
rect 78673 319426 78739 319429
rect 78673 319424 82156 319426
rect 78673 319368 78678 319424
rect 78734 319368 82156 319424
rect 78673 319366 82156 319368
rect 78673 319363 78739 319366
rect 401593 319154 401659 319157
rect 400292 319152 401659 319154
rect 400292 319096 401598 319152
rect 401654 319096 401659 319152
rect 400292 319094 401659 319096
rect 401593 319091 401659 319094
rect 401593 312082 401659 312085
rect 400292 312080 401659 312082
rect 400292 312024 401598 312080
rect 401654 312024 401659 312080
rect 400292 312022 401659 312024
rect 401593 312019 401659 312022
rect 78673 311810 78739 311813
rect 78673 311808 82156 311810
rect 78673 311752 78678 311808
rect 78734 311752 82156 311808
rect 78673 311750 82156 311752
rect 78673 311747 78739 311750
rect 579613 310858 579679 310861
rect 583520 310858 584960 310948
rect 579613 310856 584960 310858
rect 579613 310800 579618 310856
rect 579674 310800 584960 310856
rect 579613 310798 584960 310800
rect 579613 310795 579679 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3693 308818 3759 308821
rect -960 308816 3759 308818
rect -960 308760 3698 308816
rect 3754 308760 3759 308816
rect -960 308758 3759 308760
rect -960 308668 480 308758
rect 3693 308755 3759 308758
rect 401593 304874 401659 304877
rect 400292 304872 401659 304874
rect 400292 304816 401598 304872
rect 401654 304816 401659 304872
rect 400292 304814 401659 304816
rect 401593 304811 401659 304814
rect 78673 304194 78739 304197
rect 78673 304192 82156 304194
rect 78673 304136 78678 304192
rect 78734 304136 82156 304192
rect 78673 304134 82156 304136
rect 78673 304131 78739 304134
rect 578877 299162 578943 299165
rect 583520 299162 584960 299252
rect 578877 299160 584960 299162
rect 578877 299104 578882 299160
rect 578938 299104 584960 299160
rect 578877 299102 584960 299104
rect 578877 299099 578943 299102
rect 583520 299012 584960 299102
rect 401593 297802 401659 297805
rect 400292 297800 401659 297802
rect 400292 297744 401598 297800
rect 401654 297744 401659 297800
rect 400292 297742 401659 297744
rect 401593 297739 401659 297742
rect 78673 296578 78739 296581
rect 78673 296576 82156 296578
rect 78673 296520 78678 296576
rect 78734 296520 82156 296576
rect 78673 296518 82156 296520
rect 78673 296515 78739 296518
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 401593 290730 401659 290733
rect 400292 290728 401659 290730
rect 400292 290672 401598 290728
rect 401654 290672 401659 290728
rect 400292 290670 401659 290672
rect 401593 290667 401659 290670
rect 78673 288962 78739 288965
rect 78673 288960 82156 288962
rect 78673 288904 78678 288960
rect 78734 288904 82156 288960
rect 78673 288902 82156 288904
rect 78673 288899 78739 288902
rect 583520 287316 584960 287556
rect 401593 283522 401659 283525
rect 400292 283520 401659 283522
rect 400292 283464 401598 283520
rect 401654 283464 401659 283520
rect 400292 283462 401659 283464
rect 401593 283459 401659 283462
rect 78673 281346 78739 281349
rect 78673 281344 82156 281346
rect 78673 281288 78678 281344
rect 78734 281288 82156 281344
rect 78673 281286 82156 281288
rect 78673 281283 78739 281286
rect -960 280122 480 280212
rect 3509 280122 3575 280125
rect -960 280120 3575 280122
rect -960 280064 3514 280120
rect 3570 280064 3575 280120
rect -960 280062 3575 280064
rect -960 279972 480 280062
rect 3509 280059 3575 280062
rect 401593 276450 401659 276453
rect 400292 276448 401659 276450
rect 400292 276392 401598 276448
rect 401654 276392 401659 276448
rect 400292 276390 401659 276392
rect 401593 276387 401659 276390
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 78673 273730 78739 273733
rect 78673 273728 82156 273730
rect 78673 273672 78678 273728
rect 78734 273672 82156 273728
rect 78673 273670 82156 273672
rect 78673 273667 78739 273670
rect 401593 269378 401659 269381
rect 400292 269376 401659 269378
rect 400292 269320 401598 269376
rect 401654 269320 401659 269376
rect 400292 269318 401659 269320
rect 401593 269315 401659 269318
rect 78673 266114 78739 266117
rect 78673 266112 82156 266114
rect 78673 266056 78678 266112
rect 78734 266056 82156 266112
rect 78673 266054 82156 266056
rect 78673 266051 78739 266054
rect -960 265706 480 265796
rect 3601 265706 3667 265709
rect -960 265704 3667 265706
rect -960 265648 3606 265704
rect 3662 265648 3667 265704
rect -960 265646 3667 265648
rect -960 265556 480 265646
rect 3601 265643 3667 265646
rect 579797 263938 579863 263941
rect 583520 263938 584960 264028
rect 579797 263936 584960 263938
rect 579797 263880 579802 263936
rect 579858 263880 584960 263936
rect 579797 263878 584960 263880
rect 579797 263875 579863 263878
rect 583520 263788 584960 263878
rect 401593 262170 401659 262173
rect 400292 262168 401659 262170
rect 400292 262112 401598 262168
rect 401654 262112 401659 262168
rect 400292 262110 401659 262112
rect 401593 262107 401659 262110
rect 78673 258362 78739 258365
rect 78673 258360 82156 258362
rect 78673 258304 78678 258360
rect 78734 258304 82156 258360
rect 78673 258302 82156 258304
rect 78673 258299 78739 258302
rect 401593 255098 401659 255101
rect 400292 255096 401659 255098
rect 400292 255040 401598 255096
rect 401654 255040 401659 255096
rect 400292 255038 401659 255040
rect 401593 255035 401659 255038
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 78673 250746 78739 250749
rect 78673 250744 82156 250746
rect 78673 250688 78678 250744
rect 78734 250688 82156 250744
rect 78673 250686 82156 250688
rect 78673 250683 78739 250686
rect 402237 248026 402303 248029
rect 400292 248024 402303 248026
rect 400292 247968 402242 248024
rect 402298 247968 402303 248024
rect 400292 247966 402303 247968
rect 402237 247963 402303 247966
rect 78673 243130 78739 243133
rect 78673 243128 82156 243130
rect 78673 243072 78678 243128
rect 78734 243072 82156 243128
rect 78673 243070 82156 243072
rect 78673 243067 78739 243070
rect 401593 240818 401659 240821
rect 400292 240816 401659 240818
rect 400292 240760 401598 240816
rect 401654 240760 401659 240816
rect 400292 240758 401659 240760
rect 401593 240755 401659 240758
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 78673 235514 78739 235517
rect 78673 235512 82156 235514
rect 78673 235456 78678 235512
rect 78734 235456 82156 235512
rect 78673 235454 82156 235456
rect 78673 235451 78739 235454
rect 401593 233746 401659 233749
rect 400292 233744 401659 233746
rect 400292 233688 401598 233744
rect 401654 233688 401659 233744
rect 400292 233686 401659 233688
rect 401593 233683 401659 233686
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 78673 227898 78739 227901
rect 78673 227896 82156 227898
rect 78673 227840 78678 227896
rect 78734 227840 82156 227896
rect 78673 227838 82156 227840
rect 78673 227835 78739 227838
rect 401593 226674 401659 226677
rect 400292 226672 401659 226674
rect 400292 226616 401598 226672
rect 401654 226616 401659 226672
rect 400292 226614 401659 226616
rect 401593 226611 401659 226614
rect -960 222594 480 222684
rect 2957 222594 3023 222597
rect -960 222592 3023 222594
rect -960 222536 2962 222592
rect 3018 222536 3023 222592
rect -960 222534 3023 222536
rect -960 222444 480 222534
rect 2957 222531 3023 222534
rect 78673 220282 78739 220285
rect 78673 220280 82156 220282
rect 78673 220224 78678 220280
rect 78734 220224 82156 220280
rect 78673 220222 82156 220224
rect 78673 220219 78739 220222
rect 401593 219466 401659 219469
rect 400292 219464 401659 219466
rect 400292 219408 401598 219464
rect 401654 219408 401659 219464
rect 400292 219406 401659 219408
rect 401593 219403 401659 219406
rect 580257 217018 580323 217021
rect 583520 217018 584960 217108
rect 580257 217016 584960 217018
rect 580257 216960 580262 217016
rect 580318 216960 584960 217016
rect 580257 216958 584960 216960
rect 580257 216955 580323 216958
rect 583520 216868 584960 216958
rect 79317 212666 79383 212669
rect 79317 212664 82156 212666
rect 79317 212608 79322 212664
rect 79378 212608 82156 212664
rect 79317 212606 82156 212608
rect 79317 212603 79383 212606
rect 401593 212394 401659 212397
rect 400292 212392 401659 212394
rect 400292 212336 401598 212392
rect 401654 212336 401659 212392
rect 400292 212334 401659 212336
rect 401593 212331 401659 212334
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 580349 205322 580415 205325
rect 583520 205322 584960 205412
rect 580349 205320 584960 205322
rect 580349 205264 580354 205320
rect 580410 205264 584960 205320
rect 580349 205262 584960 205264
rect 580349 205259 580415 205262
rect 401593 205186 401659 205189
rect 400292 205184 401659 205186
rect 400292 205128 401598 205184
rect 401654 205128 401659 205184
rect 583520 205172 584960 205262
rect 400292 205126 401659 205128
rect 401593 205123 401659 205126
rect 79317 205050 79383 205053
rect 79317 205048 82156 205050
rect 79317 204992 79322 205048
rect 79378 204992 82156 205048
rect 79317 204990 82156 204992
rect 79317 204987 79383 204990
rect 401593 198114 401659 198117
rect 400292 198112 401659 198114
rect 400292 198056 401598 198112
rect 401654 198056 401659 198112
rect 400292 198054 401659 198056
rect 401593 198051 401659 198054
rect 79409 197434 79475 197437
rect 79409 197432 82156 197434
rect 79409 197376 79414 197432
rect 79470 197376 82156 197432
rect 79409 197374 82156 197376
rect 79409 197371 79475 197374
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 401593 191042 401659 191045
rect 400292 191040 401659 191042
rect 400292 190984 401598 191040
rect 401654 190984 401659 191040
rect 400292 190982 401659 190984
rect 401593 190979 401659 190982
rect 79317 189818 79383 189821
rect 79317 189816 82156 189818
rect 79317 189760 79322 189816
rect 79378 189760 82156 189816
rect 79317 189758 82156 189760
rect 79317 189755 79383 189758
rect 401593 183834 401659 183837
rect 400292 183832 401659 183834
rect 400292 183776 401598 183832
rect 401654 183776 401659 183832
rect 400292 183774 401659 183776
rect 401593 183771 401659 183774
rect 79501 182066 79567 182069
rect 79501 182064 82156 182066
rect 79501 182008 79506 182064
rect 79562 182008 82156 182064
rect 79501 182006 82156 182008
rect 79501 182003 79567 182006
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 402237 176762 402303 176765
rect 400292 176760 402303 176762
rect 400292 176704 402242 176760
rect 402298 176704 402303 176760
rect 400292 176702 402303 176704
rect 402237 176699 402303 176702
rect 79409 174450 79475 174453
rect 79409 174448 82156 174450
rect 79409 174392 79414 174448
rect 79470 174392 82156 174448
rect 79409 174390 82156 174392
rect 79409 174387 79475 174390
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 402237 169690 402303 169693
rect 400292 169688 402303 169690
rect 400292 169632 402242 169688
rect 402298 169632 402303 169688
rect 400292 169630 402303 169632
rect 402237 169627 402303 169630
rect 78673 166834 78739 166837
rect 78673 166832 82156 166834
rect 78673 166776 78678 166832
rect 78734 166776 82156 166832
rect 78673 166774 82156 166776
rect 78673 166771 78739 166774
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 402329 162482 402395 162485
rect 400292 162480 402395 162482
rect 400292 162424 402334 162480
rect 402390 162424 402395 162480
rect 400292 162422 402395 162424
rect 402329 162419 402395 162422
rect 79317 159218 79383 159221
rect 79317 159216 82156 159218
rect 79317 159160 79322 159216
rect 79378 159160 82156 159216
rect 79317 159158 82156 159160
rect 79317 159155 79383 159158
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 402237 155410 402303 155413
rect 400292 155408 402303 155410
rect 400292 155352 402242 155408
rect 402298 155352 402303 155408
rect 400292 155350 402303 155352
rect 402237 155347 402303 155350
rect 79685 151602 79751 151605
rect 79685 151600 82156 151602
rect 79685 151544 79690 151600
rect 79746 151544 82156 151600
rect 79685 151542 82156 151544
rect 79685 151539 79751 151542
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 402605 148338 402671 148341
rect 400292 148336 402671 148338
rect 400292 148280 402610 148336
rect 402666 148280 402671 148336
rect 400292 148278 402671 148280
rect 402605 148275 402671 148278
rect 583520 146556 584960 146796
rect 78673 143986 78739 143989
rect 78673 143984 82156 143986
rect 78673 143928 78678 143984
rect 78734 143928 82156 143984
rect 78673 143926 82156 143928
rect 78673 143923 78739 143926
rect 402513 141130 402579 141133
rect 400292 141128 402579 141130
rect 400292 141072 402518 141128
rect 402574 141072 402579 141128
rect 400292 141070 402579 141072
rect 402513 141067 402579 141070
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 79593 136370 79659 136373
rect 79593 136368 82156 136370
rect 79593 136312 79598 136368
rect 79654 136312 82156 136368
rect 79593 136310 82156 136312
rect 79593 136307 79659 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 402421 134058 402487 134061
rect 400292 134056 402487 134058
rect 400292 134000 402426 134056
rect 402482 134000 402487 134056
rect 400292 133998 402487 134000
rect 402421 133995 402487 133998
rect 79501 128754 79567 128757
rect 79501 128752 82156 128754
rect 79501 128696 79506 128752
rect 79562 128696 82156 128752
rect 79501 128694 82156 128696
rect 79501 128691 79567 128694
rect 401593 126986 401659 126989
rect 400292 126984 401659 126986
rect 400292 126928 401598 126984
rect 401654 126928 401659 126984
rect 400292 126926 401659 126928
rect 401593 126923 401659 126926
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 78673 121138 78739 121141
rect 78673 121136 82156 121138
rect 78673 121080 78678 121136
rect 78734 121080 82156 121136
rect 78673 121078 82156 121080
rect 78673 121075 78739 121078
rect 402329 119778 402395 119781
rect 400292 119776 402395 119778
rect 400292 119720 402334 119776
rect 402390 119720 402395 119776
rect 400292 119718 402395 119720
rect 402329 119715 402395 119718
rect 79409 113522 79475 113525
rect 79409 113520 82156 113522
rect 79409 113464 79414 113520
rect 79470 113464 82156 113520
rect 79409 113462 82156 113464
rect 79409 113459 79475 113462
rect 402237 112706 402303 112709
rect 400292 112704 402303 112706
rect 400292 112648 402242 112704
rect 402298 112648 402303 112704
rect 400292 112646 402303 112648
rect 402237 112643 402303 112646
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 79317 105906 79383 105909
rect 79317 105904 82156 105906
rect 79317 105848 79322 105904
rect 79378 105848 82156 105904
rect 79317 105846 82156 105848
rect 79317 105843 79383 105846
rect 401593 105634 401659 105637
rect 400292 105632 401659 105634
rect 400292 105576 401598 105632
rect 401654 105576 401659 105632
rect 400292 105574 401659 105576
rect 401593 105571 401659 105574
rect 583520 99636 584960 99876
rect 96245 96658 96311 96661
rect 96429 96658 96495 96661
rect 96245 96656 96495 96658
rect 96245 96600 96250 96656
rect 96306 96600 96434 96656
rect 96490 96600 96495 96656
rect 96245 96598 96495 96600
rect 96245 96595 96311 96598
rect 96429 96595 96495 96598
rect 104525 96658 104591 96661
rect 104709 96658 104775 96661
rect 104525 96656 104775 96658
rect 104525 96600 104530 96656
rect 104586 96600 104714 96656
rect 104770 96600 104775 96656
rect 104525 96598 104775 96600
rect 104525 96595 104591 96598
rect 104709 96595 104775 96598
rect 151445 96658 151511 96661
rect 151629 96658 151695 96661
rect 151445 96656 151695 96658
rect 151445 96600 151450 96656
rect 151506 96600 151634 96656
rect 151690 96600 151695 96656
rect 151445 96598 151695 96600
rect 151445 96595 151511 96598
rect 151629 96595 151695 96598
rect 239765 96658 239831 96661
rect 239949 96658 240015 96661
rect 239765 96656 240015 96658
rect 239765 96600 239770 96656
rect 239826 96600 239954 96656
rect 240010 96600 240015 96656
rect 239765 96598 240015 96600
rect 239765 96595 239831 96598
rect 239949 96595 240015 96598
rect 274357 96658 274423 96661
rect 274541 96658 274607 96661
rect 274357 96656 274607 96658
rect 274357 96600 274362 96656
rect 274418 96600 274546 96656
rect 274602 96600 274607 96656
rect 274357 96598 274607 96600
rect 274357 96595 274423 96598
rect 274541 96595 274607 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 370681 87002 370747 87005
rect 370865 87002 370931 87005
rect 370681 87000 370931 87002
rect 370681 86944 370686 87000
rect 370742 86944 370870 87000
rect 370926 86944 370931 87000
rect 370681 86942 370931 86944
rect 370681 86939 370747 86942
rect 370865 86939 370931 86942
rect 91921 85506 91987 85509
rect 92197 85506 92263 85509
rect 91921 85504 92263 85506
rect 91921 85448 91926 85504
rect 91982 85448 92202 85504
rect 92258 85448 92263 85504
rect 91921 85446 92263 85448
rect 91921 85443 91987 85446
rect 92197 85443 92263 85446
rect 96337 80748 96403 80749
rect 96286 80746 96292 80748
rect 96246 80686 96292 80746
rect 96356 80744 96403 80748
rect 96398 80688 96403 80744
rect 96286 80684 96292 80686
rect 96356 80684 96403 80688
rect 96337 80683 96403 80684
rect 151486 80140 151492 80204
rect 151556 80202 151562 80204
rect 151629 80202 151695 80205
rect 151556 80200 151695 80202
rect 151556 80144 151634 80200
rect 151690 80144 151695 80200
rect 151556 80142 151695 80144
rect 151556 80140 151562 80142
rect 151629 80139 151695 80142
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 151537 77348 151603 77349
rect 151486 77284 151492 77348
rect 151556 77346 151603 77348
rect 227069 77346 227135 77349
rect 227253 77346 227319 77349
rect 151556 77344 151648 77346
rect 151598 77288 151648 77344
rect 151556 77286 151648 77288
rect 227069 77344 227319 77346
rect 227069 77288 227074 77344
rect 227130 77288 227258 77344
rect 227314 77288 227319 77344
rect 227069 77286 227319 77288
rect 151556 77284 151603 77286
rect 151537 77283 151603 77284
rect 227069 77283 227135 77286
rect 227253 77283 227319 77286
rect 341701 77346 341767 77349
rect 341885 77346 341951 77349
rect 341701 77344 341951 77346
rect 341701 77288 341706 77344
rect 341762 77288 341890 77344
rect 341946 77288 341951 77344
rect 341701 77286 341951 77288
rect 341701 77283 341767 77286
rect 341885 77283 341951 77286
rect 550633 77210 550699 77213
rect 550909 77210 550975 77213
rect 550633 77208 550975 77210
rect 550633 77152 550638 77208
rect 550694 77152 550914 77208
rect 550970 77152 550975 77208
rect 550633 77150 550975 77152
rect 550633 77147 550699 77150
rect 550909 77147 550975 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 96286 67764 96292 67828
rect 96356 67826 96362 67828
rect 96356 67766 96538 67826
rect 96356 67764 96362 67766
rect 96337 67690 96403 67693
rect 96478 67690 96538 67766
rect 227253 67824 227319 67829
rect 227253 67768 227258 67824
rect 227314 67768 227319 67824
rect 227253 67763 227319 67768
rect 341885 67824 341951 67829
rect 341885 67768 341890 67824
rect 341946 67768 341951 67824
rect 341885 67763 341951 67768
rect 227256 67693 227316 67763
rect 341888 67693 341948 67763
rect 96337 67688 96538 67690
rect 96337 67632 96342 67688
rect 96398 67632 96538 67688
rect 96337 67630 96538 67632
rect 227253 67688 227319 67693
rect 227253 67632 227258 67688
rect 227314 67632 227319 67688
rect 96337 67627 96403 67630
rect 227253 67627 227319 67632
rect 341885 67688 341951 67693
rect 341885 67632 341890 67688
rect 341946 67632 341951 67688
rect 341885 67627 341951 67632
rect 197721 67554 197787 67557
rect 197997 67554 198063 67557
rect 197721 67552 198063 67554
rect 197721 67496 197726 67552
rect 197782 67496 198002 67552
rect 198058 67496 198063 67552
rect 197721 67494 198063 67496
rect 197721 67491 197787 67494
rect 197997 67491 198063 67494
rect 215017 64970 215083 64973
rect 215201 64970 215267 64973
rect 215017 64968 215267 64970
rect 215017 64912 215022 64968
rect 215078 64912 215206 64968
rect 215262 64912 215267 64968
rect 215017 64910 215267 64912
rect 215017 64907 215083 64910
rect 215201 64907 215267 64910
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 578877 64562 578943 64565
rect 583520 64562 584960 64652
rect 578877 64560 584960 64562
rect 578877 64504 578882 64560
rect 578938 64504 584960 64560
rect 578877 64502 584960 64504
rect 578877 64499 578943 64502
rect 583520 64412 584960 64502
rect 227437 61436 227503 61437
rect 227437 61434 227484 61436
rect 227392 61432 227484 61434
rect 227392 61376 227442 61432
rect 227392 61374 227484 61376
rect 227437 61372 227484 61374
rect 227548 61372 227554 61436
rect 227437 61371 227503 61372
rect 215017 60754 215083 60757
rect 215150 60754 215156 60756
rect 215017 60752 215156 60754
rect 215017 60696 215022 60752
rect 215078 60696 215156 60752
rect 215017 60694 215156 60696
rect 215017 60691 215083 60694
rect 215150 60692 215156 60694
rect 215220 60692 215226 60756
rect 550633 58170 550699 58173
rect 550590 58168 550699 58170
rect 550590 58112 550638 58168
rect 550694 58112 550699 58168
rect 550590 58107 550699 58112
rect 550590 58037 550650 58107
rect 550590 58032 550699 58037
rect 550590 57976 550638 58032
rect 550694 57976 550699 58032
rect 550590 57974 550699 57976
rect 550633 57971 550699 57974
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 568573 48514 568639 48517
rect 568438 48512 568639 48514
rect 568438 48456 568578 48512
rect 568634 48456 568639 48512
rect 568438 48454 568639 48456
rect 215017 48378 215083 48381
rect 215150 48378 215156 48380
rect 215017 48376 215156 48378
rect 215017 48320 215022 48376
rect 215078 48320 215156 48376
rect 215017 48318 215156 48320
rect 215017 48315 215083 48318
rect 215150 48316 215156 48318
rect 215220 48316 215226 48380
rect 227345 48378 227411 48381
rect 227478 48378 227484 48380
rect 227345 48376 227484 48378
rect 227345 48320 227350 48376
rect 227406 48320 227484 48376
rect 227345 48318 227484 48320
rect 227345 48315 227411 48318
rect 227478 48316 227484 48318
rect 227548 48316 227554 48380
rect 568438 48378 568498 48454
rect 568573 48451 568639 48454
rect 568573 48378 568639 48381
rect 568438 48376 568639 48378
rect 568438 48320 568578 48376
rect 568634 48320 568639 48376
rect 568438 48318 568639 48320
rect 568573 48315 568639 48318
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 198549 29066 198615 29069
rect 198733 29066 198799 29069
rect 198549 29064 198799 29066
rect 198549 29008 198554 29064
rect 198610 29008 198738 29064
rect 198794 29008 198799 29064
rect 198549 29006 198799 29008
rect 198549 29003 198615 29006
rect 198733 29003 198799 29006
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 568021 8258 568087 8261
rect 567886 8256 568087 8258
rect 567886 8200 568026 8256
rect 568082 8200 568087 8256
rect 567886 8198 568087 8200
rect 567886 8122 567946 8198
rect 568021 8195 568087 8198
rect 568205 8122 568271 8125
rect 567886 8120 568271 8122
rect 567886 8064 568210 8120
rect 568266 8064 568271 8120
rect 567886 8062 568271 8064
rect 568205 8059 568271 8062
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< via3 >>
rect 299612 569936 299676 569940
rect 299612 569880 299662 569936
rect 299662 569880 299676 569936
rect 299612 569876 299676 569880
rect 299612 560416 299676 560420
rect 299612 560360 299626 560416
rect 299626 560360 299676 560416
rect 299612 560356 299676 560360
rect 347820 502284 347884 502348
rect 347820 492688 347884 492692
rect 347820 492632 347870 492688
rect 347870 492632 347884 492688
rect 347820 492628 347884 492632
rect 96292 80744 96356 80748
rect 96292 80688 96342 80744
rect 96342 80688 96356 80744
rect 96292 80684 96356 80688
rect 151492 80140 151556 80204
rect 151492 77344 151556 77348
rect 151492 77288 151542 77344
rect 151542 77288 151556 77344
rect 151492 77284 151556 77288
rect 96292 67764 96356 67828
rect 227484 61432 227548 61436
rect 227484 61376 227498 61432
rect 227498 61376 227548 61432
rect 227484 61372 227548 61376
rect 215156 60692 215220 60756
rect 215156 48316 215220 48380
rect 227484 48316 227548 48380
<< metal4 >>
rect -4876 707718 -4276 707740
rect -4876 707482 -4694 707718
rect -4458 707482 -4276 707718
rect -4876 707398 -4276 707482
rect -4876 707162 -4694 707398
rect -4458 707162 -4276 707398
rect -4876 672054 -4276 707162
rect -4876 671818 -4694 672054
rect -4458 671818 -4276 672054
rect -4876 671734 -4276 671818
rect -4876 671498 -4694 671734
rect -4458 671498 -4276 671734
rect -4876 636054 -4276 671498
rect -4876 635818 -4694 636054
rect -4458 635818 -4276 636054
rect -4876 635734 -4276 635818
rect -4876 635498 -4694 635734
rect -4458 635498 -4276 635734
rect -4876 600054 -4276 635498
rect -4876 599818 -4694 600054
rect -4458 599818 -4276 600054
rect -4876 599734 -4276 599818
rect -4876 599498 -4694 599734
rect -4458 599498 -4276 599734
rect -4876 564054 -4276 599498
rect -4876 563818 -4694 564054
rect -4458 563818 -4276 564054
rect -4876 563734 -4276 563818
rect -4876 563498 -4694 563734
rect -4458 563498 -4276 563734
rect -4876 528054 -4276 563498
rect -4876 527818 -4694 528054
rect -4458 527818 -4276 528054
rect -4876 527734 -4276 527818
rect -4876 527498 -4694 527734
rect -4458 527498 -4276 527734
rect -4876 492054 -4276 527498
rect -4876 491818 -4694 492054
rect -4458 491818 -4276 492054
rect -4876 491734 -4276 491818
rect -4876 491498 -4694 491734
rect -4458 491498 -4276 491734
rect -4876 456054 -4276 491498
rect -4876 455818 -4694 456054
rect -4458 455818 -4276 456054
rect -4876 455734 -4276 455818
rect -4876 455498 -4694 455734
rect -4458 455498 -4276 455734
rect -4876 420054 -4276 455498
rect -4876 419818 -4694 420054
rect -4458 419818 -4276 420054
rect -4876 419734 -4276 419818
rect -4876 419498 -4694 419734
rect -4458 419498 -4276 419734
rect -4876 384054 -4276 419498
rect -4876 383818 -4694 384054
rect -4458 383818 -4276 384054
rect -4876 383734 -4276 383818
rect -4876 383498 -4694 383734
rect -4458 383498 -4276 383734
rect -4876 348054 -4276 383498
rect -4876 347818 -4694 348054
rect -4458 347818 -4276 348054
rect -4876 347734 -4276 347818
rect -4876 347498 -4694 347734
rect -4458 347498 -4276 347734
rect -4876 312054 -4276 347498
rect -4876 311818 -4694 312054
rect -4458 311818 -4276 312054
rect -4876 311734 -4276 311818
rect -4876 311498 -4694 311734
rect -4458 311498 -4276 311734
rect -4876 276054 -4276 311498
rect -4876 275818 -4694 276054
rect -4458 275818 -4276 276054
rect -4876 275734 -4276 275818
rect -4876 275498 -4694 275734
rect -4458 275498 -4276 275734
rect -4876 240054 -4276 275498
rect -4876 239818 -4694 240054
rect -4458 239818 -4276 240054
rect -4876 239734 -4276 239818
rect -4876 239498 -4694 239734
rect -4458 239498 -4276 239734
rect -4876 204054 -4276 239498
rect -4876 203818 -4694 204054
rect -4458 203818 -4276 204054
rect -4876 203734 -4276 203818
rect -4876 203498 -4694 203734
rect -4458 203498 -4276 203734
rect -4876 168054 -4276 203498
rect -4876 167818 -4694 168054
rect -4458 167818 -4276 168054
rect -4876 167734 -4276 167818
rect -4876 167498 -4694 167734
rect -4458 167498 -4276 167734
rect -4876 132054 -4276 167498
rect -4876 131818 -4694 132054
rect -4458 131818 -4276 132054
rect -4876 131734 -4276 131818
rect -4876 131498 -4694 131734
rect -4458 131498 -4276 131734
rect -4876 96054 -4276 131498
rect -4876 95818 -4694 96054
rect -4458 95818 -4276 96054
rect -4876 95734 -4276 95818
rect -4876 95498 -4694 95734
rect -4458 95498 -4276 95734
rect -4876 60054 -4276 95498
rect -4876 59818 -4694 60054
rect -4458 59818 -4276 60054
rect -4876 59734 -4276 59818
rect -4876 59498 -4694 59734
rect -4458 59498 -4276 59734
rect -4876 24054 -4276 59498
rect -4876 23818 -4694 24054
rect -4458 23818 -4276 24054
rect -4876 23734 -4276 23818
rect -4876 23498 -4694 23734
rect -4458 23498 -4276 23734
rect -4876 -3226 -4276 23498
rect -3916 706758 -3316 706780
rect -3916 706522 -3734 706758
rect -3498 706522 -3316 706758
rect -3916 706438 -3316 706522
rect -3916 706202 -3734 706438
rect -3498 706202 -3316 706438
rect -3916 690054 -3316 706202
rect 4404 706758 5004 707740
rect 4404 706522 4586 706758
rect 4822 706522 5004 706758
rect 4404 706438 5004 706522
rect 4404 706202 4586 706438
rect 4822 706202 5004 706438
rect -3916 689818 -3734 690054
rect -3498 689818 -3316 690054
rect -3916 689734 -3316 689818
rect -3916 689498 -3734 689734
rect -3498 689498 -3316 689734
rect -3916 654054 -3316 689498
rect -3916 653818 -3734 654054
rect -3498 653818 -3316 654054
rect -3916 653734 -3316 653818
rect -3916 653498 -3734 653734
rect -3498 653498 -3316 653734
rect -3916 618054 -3316 653498
rect -3916 617818 -3734 618054
rect -3498 617818 -3316 618054
rect -3916 617734 -3316 617818
rect -3916 617498 -3734 617734
rect -3498 617498 -3316 617734
rect -3916 582054 -3316 617498
rect -3916 581818 -3734 582054
rect -3498 581818 -3316 582054
rect -3916 581734 -3316 581818
rect -3916 581498 -3734 581734
rect -3498 581498 -3316 581734
rect -3916 546054 -3316 581498
rect -3916 545818 -3734 546054
rect -3498 545818 -3316 546054
rect -3916 545734 -3316 545818
rect -3916 545498 -3734 545734
rect -3498 545498 -3316 545734
rect -3916 510054 -3316 545498
rect -3916 509818 -3734 510054
rect -3498 509818 -3316 510054
rect -3916 509734 -3316 509818
rect -3916 509498 -3734 509734
rect -3498 509498 -3316 509734
rect -3916 474054 -3316 509498
rect -3916 473818 -3734 474054
rect -3498 473818 -3316 474054
rect -3916 473734 -3316 473818
rect -3916 473498 -3734 473734
rect -3498 473498 -3316 473734
rect -3916 438054 -3316 473498
rect -3916 437818 -3734 438054
rect -3498 437818 -3316 438054
rect -3916 437734 -3316 437818
rect -3916 437498 -3734 437734
rect -3498 437498 -3316 437734
rect -3916 402054 -3316 437498
rect -3916 401818 -3734 402054
rect -3498 401818 -3316 402054
rect -3916 401734 -3316 401818
rect -3916 401498 -3734 401734
rect -3498 401498 -3316 401734
rect -3916 366054 -3316 401498
rect -3916 365818 -3734 366054
rect -3498 365818 -3316 366054
rect -3916 365734 -3316 365818
rect -3916 365498 -3734 365734
rect -3498 365498 -3316 365734
rect -3916 330054 -3316 365498
rect -3916 329818 -3734 330054
rect -3498 329818 -3316 330054
rect -3916 329734 -3316 329818
rect -3916 329498 -3734 329734
rect -3498 329498 -3316 329734
rect -3916 294054 -3316 329498
rect -3916 293818 -3734 294054
rect -3498 293818 -3316 294054
rect -3916 293734 -3316 293818
rect -3916 293498 -3734 293734
rect -3498 293498 -3316 293734
rect -3916 258054 -3316 293498
rect -3916 257818 -3734 258054
rect -3498 257818 -3316 258054
rect -3916 257734 -3316 257818
rect -3916 257498 -3734 257734
rect -3498 257498 -3316 257734
rect -3916 222054 -3316 257498
rect -3916 221818 -3734 222054
rect -3498 221818 -3316 222054
rect -3916 221734 -3316 221818
rect -3916 221498 -3734 221734
rect -3498 221498 -3316 221734
rect -3916 186054 -3316 221498
rect -3916 185818 -3734 186054
rect -3498 185818 -3316 186054
rect -3916 185734 -3316 185818
rect -3916 185498 -3734 185734
rect -3498 185498 -3316 185734
rect -3916 150054 -3316 185498
rect -3916 149818 -3734 150054
rect -3498 149818 -3316 150054
rect -3916 149734 -3316 149818
rect -3916 149498 -3734 149734
rect -3498 149498 -3316 149734
rect -3916 114054 -3316 149498
rect -3916 113818 -3734 114054
rect -3498 113818 -3316 114054
rect -3916 113734 -3316 113818
rect -3916 113498 -3734 113734
rect -3498 113498 -3316 113734
rect -3916 78054 -3316 113498
rect -3916 77818 -3734 78054
rect -3498 77818 -3316 78054
rect -3916 77734 -3316 77818
rect -3916 77498 -3734 77734
rect -3498 77498 -3316 77734
rect -3916 42054 -3316 77498
rect -3916 41818 -3734 42054
rect -3498 41818 -3316 42054
rect -3916 41734 -3316 41818
rect -3916 41498 -3734 41734
rect -3498 41498 -3316 41734
rect -3916 6054 -3316 41498
rect -3916 5818 -3734 6054
rect -3498 5818 -3316 6054
rect -3916 5734 -3316 5818
rect -3916 5498 -3734 5734
rect -3498 5498 -3316 5734
rect -3916 -2266 -3316 5498
rect -2956 705798 -2356 705820
rect -2956 705562 -2774 705798
rect -2538 705562 -2356 705798
rect -2956 705478 -2356 705562
rect -2956 705242 -2774 705478
rect -2538 705242 -2356 705478
rect -2956 668454 -2356 705242
rect -2956 668218 -2774 668454
rect -2538 668218 -2356 668454
rect -2956 668134 -2356 668218
rect -2956 667898 -2774 668134
rect -2538 667898 -2356 668134
rect -2956 632454 -2356 667898
rect -2956 632218 -2774 632454
rect -2538 632218 -2356 632454
rect -2956 632134 -2356 632218
rect -2956 631898 -2774 632134
rect -2538 631898 -2356 632134
rect -2956 596454 -2356 631898
rect -2956 596218 -2774 596454
rect -2538 596218 -2356 596454
rect -2956 596134 -2356 596218
rect -2956 595898 -2774 596134
rect -2538 595898 -2356 596134
rect -2956 560454 -2356 595898
rect -2956 560218 -2774 560454
rect -2538 560218 -2356 560454
rect -2956 560134 -2356 560218
rect -2956 559898 -2774 560134
rect -2538 559898 -2356 560134
rect -2956 524454 -2356 559898
rect -2956 524218 -2774 524454
rect -2538 524218 -2356 524454
rect -2956 524134 -2356 524218
rect -2956 523898 -2774 524134
rect -2538 523898 -2356 524134
rect -2956 488454 -2356 523898
rect -2956 488218 -2774 488454
rect -2538 488218 -2356 488454
rect -2956 488134 -2356 488218
rect -2956 487898 -2774 488134
rect -2538 487898 -2356 488134
rect -2956 452454 -2356 487898
rect -2956 452218 -2774 452454
rect -2538 452218 -2356 452454
rect -2956 452134 -2356 452218
rect -2956 451898 -2774 452134
rect -2538 451898 -2356 452134
rect -2956 416454 -2356 451898
rect -2956 416218 -2774 416454
rect -2538 416218 -2356 416454
rect -2956 416134 -2356 416218
rect -2956 415898 -2774 416134
rect -2538 415898 -2356 416134
rect -2956 380454 -2356 415898
rect -2956 380218 -2774 380454
rect -2538 380218 -2356 380454
rect -2956 380134 -2356 380218
rect -2956 379898 -2774 380134
rect -2538 379898 -2356 380134
rect -2956 344454 -2356 379898
rect -2956 344218 -2774 344454
rect -2538 344218 -2356 344454
rect -2956 344134 -2356 344218
rect -2956 343898 -2774 344134
rect -2538 343898 -2356 344134
rect -2956 308454 -2356 343898
rect -2956 308218 -2774 308454
rect -2538 308218 -2356 308454
rect -2956 308134 -2356 308218
rect -2956 307898 -2774 308134
rect -2538 307898 -2356 308134
rect -2956 272454 -2356 307898
rect -2956 272218 -2774 272454
rect -2538 272218 -2356 272454
rect -2956 272134 -2356 272218
rect -2956 271898 -2774 272134
rect -2538 271898 -2356 272134
rect -2956 236454 -2356 271898
rect -2956 236218 -2774 236454
rect -2538 236218 -2356 236454
rect -2956 236134 -2356 236218
rect -2956 235898 -2774 236134
rect -2538 235898 -2356 236134
rect -2956 200454 -2356 235898
rect -2956 200218 -2774 200454
rect -2538 200218 -2356 200454
rect -2956 200134 -2356 200218
rect -2956 199898 -2774 200134
rect -2538 199898 -2356 200134
rect -2956 164454 -2356 199898
rect -2956 164218 -2774 164454
rect -2538 164218 -2356 164454
rect -2956 164134 -2356 164218
rect -2956 163898 -2774 164134
rect -2538 163898 -2356 164134
rect -2956 128454 -2356 163898
rect -2956 128218 -2774 128454
rect -2538 128218 -2356 128454
rect -2956 128134 -2356 128218
rect -2956 127898 -2774 128134
rect -2538 127898 -2356 128134
rect -2956 92454 -2356 127898
rect -2956 92218 -2774 92454
rect -2538 92218 -2356 92454
rect -2956 92134 -2356 92218
rect -2956 91898 -2774 92134
rect -2538 91898 -2356 92134
rect -2956 56454 -2356 91898
rect -2956 56218 -2774 56454
rect -2538 56218 -2356 56454
rect -2956 56134 -2356 56218
rect -2956 55898 -2774 56134
rect -2538 55898 -2356 56134
rect -2956 20454 -2356 55898
rect -2956 20218 -2774 20454
rect -2538 20218 -2356 20454
rect -2956 20134 -2356 20218
rect -2956 19898 -2774 20134
rect -2538 19898 -2356 20134
rect -2956 -1306 -2356 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705820
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2956 -1542 -2774 -1306
rect -2538 -1542 -2356 -1306
rect -2956 -1626 -2356 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 -2356 -1626
rect -2956 -1884 -2356 -1862
rect 804 -1884 1404 -902
rect 4404 690054 5004 706202
rect 22404 707718 23004 707740
rect 22404 707482 22586 707718
rect 22822 707482 23004 707718
rect 22404 707398 23004 707482
rect 22404 707162 22586 707398
rect 22822 707162 23004 707398
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3916 -2502 -3734 -2266
rect -3498 -2502 -3316 -2266
rect -3916 -2586 -3316 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 -3316 -2586
rect -3916 -2844 -3316 -2822
rect 4404 -2266 5004 5498
rect 18804 705798 19404 705820
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668454 19404 705242
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1306 19404 19898
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1884 19404 -1862
rect 22404 672054 23004 707162
rect 40404 706758 41004 707740
rect 40404 706522 40586 706758
rect 40822 706522 41004 706758
rect 40404 706438 41004 706522
rect 40404 706202 40586 706438
rect 40822 706202 41004 706438
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 4404 -2502 4586 -2266
rect 4822 -2502 5004 -2266
rect 4404 -2586 5004 -2502
rect 4404 -2822 4586 -2586
rect 4822 -2822 5004 -2586
rect -4876 -3462 -4694 -3226
rect -4458 -3462 -4276 -3226
rect -4876 -3546 -4276 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 -4276 -3546
rect -4876 -3804 -4276 -3782
rect 4404 -3804 5004 -2822
rect 22404 -3226 23004 23498
rect 36804 704838 37404 705820
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1884 37404 -902
rect 40404 690054 41004 706202
rect 58404 707718 59004 707740
rect 58404 707482 58586 707718
rect 58822 707482 59004 707718
rect 58404 707398 59004 707482
rect 58404 707162 58586 707398
rect 58822 707162 59004 707398
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 22404 -3462 22586 -3226
rect 22822 -3462 23004 -3226
rect 22404 -3546 23004 -3462
rect 22404 -3782 22586 -3546
rect 22822 -3782 23004 -3546
rect 22404 -3804 23004 -3782
rect 40404 -2266 41004 5498
rect 54804 705798 55404 705820
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668454 55404 705242
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1306 55404 19898
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1884 55404 -1862
rect 58404 672054 59004 707162
rect 76404 706758 77004 707740
rect 76404 706522 76586 706758
rect 76822 706522 77004 706758
rect 76404 706438 77004 706522
rect 76404 706202 76586 706438
rect 76822 706202 77004 706438
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 40404 -2502 40586 -2266
rect 40822 -2502 41004 -2266
rect 40404 -2586 41004 -2502
rect 40404 -2822 40586 -2586
rect 40822 -2822 41004 -2586
rect 40404 -3804 41004 -2822
rect 58404 -3226 59004 23498
rect 72804 704838 73404 705820
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1884 73404 -902
rect 76404 690054 77004 706202
rect 94404 707718 95004 707740
rect 94404 707482 94586 707718
rect 94822 707482 95004 707718
rect 94404 707398 95004 707482
rect 94404 707162 94586 707398
rect 94822 707162 95004 707398
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 90804 705798 91404 705820
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668454 91404 705242
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 422437 91404 451898
rect 94404 672054 95004 707162
rect 112404 706758 113004 707740
rect 112404 706522 112586 706758
rect 112822 706522 113004 706758
rect 112404 706438 113004 706522
rect 112404 706202 112586 706438
rect 112822 706202 113004 706438
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 422437 95004 455498
rect 108804 704838 109404 705820
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 422437 109404 433898
rect 112404 690054 113004 706202
rect 130404 707718 131004 707740
rect 130404 707482 130586 707718
rect 130822 707482 131004 707718
rect 130404 707398 131004 707482
rect 130404 707162 130586 707398
rect 130822 707162 131004 707398
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 422437 113004 437498
rect 126804 705798 127404 705820
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668454 127404 705242
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 422437 127404 451898
rect 130404 672054 131004 707162
rect 148404 706758 149004 707740
rect 148404 706522 148586 706758
rect 148822 706522 149004 706758
rect 148404 706438 149004 706522
rect 148404 706202 148586 706438
rect 148822 706202 149004 706438
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 422437 131004 455498
rect 144804 704838 145404 705820
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 422437 145404 433898
rect 148404 690054 149004 706202
rect 166404 707718 167004 707740
rect 166404 707482 166586 707718
rect 166822 707482 167004 707718
rect 166404 707398 167004 707482
rect 166404 707162 166586 707398
rect 166822 707162 167004 707398
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 422437 149004 437498
rect 162804 705798 163404 705820
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668454 163404 705242
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 422437 163404 451898
rect 166404 672054 167004 707162
rect 184404 706758 185004 707740
rect 184404 706522 184586 706758
rect 184822 706522 185004 706758
rect 184404 706438 185004 706522
rect 184404 706202 184586 706438
rect 184822 706202 185004 706438
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 422437 167004 455498
rect 180804 704838 181404 705820
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 422437 181404 433898
rect 184404 690054 185004 706202
rect 202404 707718 203004 707740
rect 202404 707482 202586 707718
rect 202822 707482 203004 707718
rect 202404 707398 203004 707482
rect 202404 707162 202586 707398
rect 202822 707162 203004 707398
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 422437 185004 437498
rect 198804 705798 199404 705820
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668454 199404 705242
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 422437 199404 451898
rect 202404 672054 203004 707162
rect 220404 706758 221004 707740
rect 220404 706522 220586 706758
rect 220822 706522 221004 706758
rect 220404 706438 221004 706522
rect 220404 706202 220586 706438
rect 220822 706202 221004 706438
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 422437 203004 455498
rect 216804 704838 217404 705820
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 422437 217404 433898
rect 220404 690054 221004 706202
rect 238404 707718 239004 707740
rect 238404 707482 238586 707718
rect 238822 707482 239004 707718
rect 238404 707398 239004 707482
rect 238404 707162 238586 707398
rect 238822 707162 239004 707398
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 422437 221004 437498
rect 234804 705798 235404 705820
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668454 235404 705242
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 422437 235404 451898
rect 238404 672054 239004 707162
rect 256404 706758 257004 707740
rect 256404 706522 256586 706758
rect 256822 706522 257004 706758
rect 256404 706438 257004 706522
rect 256404 706202 256586 706438
rect 256822 706202 257004 706438
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 422437 239004 455498
rect 252804 704838 253404 705820
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 422437 253404 433898
rect 256404 690054 257004 706202
rect 274404 707718 275004 707740
rect 274404 707482 274586 707718
rect 274822 707482 275004 707718
rect 274404 707398 275004 707482
rect 274404 707162 274586 707398
rect 274822 707162 275004 707398
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 422437 257004 437498
rect 270804 705798 271404 705820
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668454 271404 705242
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 422437 271404 451898
rect 274404 672054 275004 707162
rect 292404 706758 293004 707740
rect 292404 706522 292586 706758
rect 292822 706522 293004 706758
rect 292404 706438 293004 706522
rect 292404 706202 292586 706438
rect 292822 706202 293004 706438
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 422437 275004 455498
rect 288804 704838 289404 705820
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 422437 289404 433898
rect 292404 690054 293004 706202
rect 310404 707718 311004 707740
rect 310404 707482 310586 707718
rect 310822 707482 311004 707718
rect 310404 707398 311004 707482
rect 310404 707162 310586 707398
rect 310822 707162 311004 707398
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 306804 705798 307404 705820
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668454 307404 705242
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 299611 569940 299677 569941
rect 299611 569876 299612 569940
rect 299676 569876 299677 569940
rect 299611 569875 299677 569876
rect 299614 560421 299674 569875
rect 306804 560454 307404 595898
rect 299611 560420 299677 560421
rect 299611 560356 299612 560420
rect 299676 560356 299677 560420
rect 299611 560355 299677 560356
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 422437 293004 437498
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 422437 307404 451898
rect 310404 672054 311004 707162
rect 328404 706758 329004 707740
rect 328404 706522 328586 706758
rect 328822 706522 329004 706758
rect 328404 706438 329004 706522
rect 328404 706202 328586 706438
rect 328822 706202 329004 706438
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 422437 311004 455498
rect 324804 704838 325404 705820
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 422437 325404 433898
rect 328404 690054 329004 706202
rect 346404 707718 347004 707740
rect 346404 707482 346586 707718
rect 346822 707482 347004 707718
rect 346404 707398 347004 707482
rect 346404 707162 346586 707398
rect 346822 707162 347004 707398
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 422437 329004 437498
rect 342804 705798 343404 705820
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668454 343404 705242
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 422437 343404 451898
rect 346404 672054 347004 707162
rect 364404 706758 365004 707740
rect 364404 706522 364586 706758
rect 364822 706522 365004 706758
rect 364404 706438 365004 706522
rect 364404 706202 364586 706438
rect 364822 706202 365004 706438
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 360804 704838 361404 705820
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 347819 502348 347885 502349
rect 347819 502284 347820 502348
rect 347884 502284 347885 502348
rect 347819 502283 347885 502284
rect 347822 492693 347882 502283
rect 347819 492692 347885 492693
rect 347819 492628 347820 492692
rect 347884 492628 347885 492692
rect 347819 492627 347885 492628
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 422437 347004 455498
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 422437 361404 433898
rect 364404 690054 365004 706202
rect 382404 707718 383004 707740
rect 382404 707482 382586 707718
rect 382822 707482 383004 707718
rect 382404 707398 383004 707482
rect 382404 707162 382586 707398
rect 382822 707162 383004 707398
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 422437 365004 437498
rect 378804 705798 379404 705820
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668454 379404 705242
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 422437 379404 451898
rect 382404 672054 383004 707162
rect 400404 706758 401004 707740
rect 400404 706522 400586 706758
rect 400822 706522 401004 706758
rect 400404 706438 401004 706522
rect 400404 706202 400586 706438
rect 400822 706202 401004 706438
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 422437 383004 455498
rect 396804 704838 397404 705820
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 422437 397404 433898
rect 400404 690054 401004 706202
rect 418404 707718 419004 707740
rect 418404 707482 418586 707718
rect 418822 707482 419004 707718
rect 418404 707398 419004 707482
rect 418404 707162 418586 707398
rect 418822 707162 419004 707398
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 101568 420054 101888 420076
rect 101568 419818 101610 420054
rect 101846 419818 101888 420054
rect 101568 419734 101888 419818
rect 101568 419498 101610 419734
rect 101846 419498 101888 419734
rect 101568 419476 101888 419498
rect 101568 416454 101888 416476
rect 101568 416218 101610 416454
rect 101846 416218 101888 416454
rect 101568 416134 101888 416218
rect 101568 415898 101610 416134
rect 101846 415898 101888 416134
rect 101568 415876 101888 415898
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 86208 402054 86528 402076
rect 86208 401818 86250 402054
rect 86486 401818 86528 402054
rect 86208 401734 86528 401818
rect 86208 401498 86250 401734
rect 86486 401498 86528 401734
rect 86208 401476 86528 401498
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 86208 398454 86528 398476
rect 86208 398218 86250 398454
rect 86486 398218 86528 398454
rect 86208 398134 86528 398218
rect 86208 397898 86250 398134
rect 86486 397898 86528 398134
rect 86208 397876 86528 397898
rect 101568 384054 101888 384076
rect 101568 383818 101610 384054
rect 101846 383818 101888 384054
rect 101568 383734 101888 383818
rect 101568 383498 101610 383734
rect 101846 383498 101888 383734
rect 101568 383476 101888 383498
rect 101568 380454 101888 380476
rect 101568 380218 101610 380454
rect 101846 380218 101888 380454
rect 101568 380134 101888 380218
rect 101568 379898 101610 380134
rect 101846 379898 101888 380134
rect 101568 379876 101888 379898
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 86208 366054 86528 366076
rect 86208 365818 86250 366054
rect 86486 365818 86528 366054
rect 86208 365734 86528 365818
rect 86208 365498 86250 365734
rect 86486 365498 86528 365734
rect 86208 365476 86528 365498
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 86208 362454 86528 362476
rect 86208 362218 86250 362454
rect 86486 362218 86528 362454
rect 86208 362134 86528 362218
rect 86208 361898 86250 362134
rect 86486 361898 86528 362134
rect 86208 361876 86528 361898
rect 101568 348054 101888 348076
rect 101568 347818 101610 348054
rect 101846 347818 101888 348054
rect 101568 347734 101888 347818
rect 101568 347498 101610 347734
rect 101846 347498 101888 347734
rect 101568 347476 101888 347498
rect 101568 344454 101888 344476
rect 101568 344218 101610 344454
rect 101846 344218 101888 344454
rect 101568 344134 101888 344218
rect 101568 343898 101610 344134
rect 101846 343898 101888 344134
rect 101568 343876 101888 343898
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 86208 330054 86528 330076
rect 86208 329818 86250 330054
rect 86486 329818 86528 330054
rect 86208 329734 86528 329818
rect 86208 329498 86250 329734
rect 86486 329498 86528 329734
rect 86208 329476 86528 329498
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 86208 326454 86528 326476
rect 86208 326218 86250 326454
rect 86486 326218 86528 326454
rect 86208 326134 86528 326218
rect 86208 325898 86250 326134
rect 86486 325898 86528 326134
rect 86208 325876 86528 325898
rect 101568 312054 101888 312076
rect 101568 311818 101610 312054
rect 101846 311818 101888 312054
rect 101568 311734 101888 311818
rect 101568 311498 101610 311734
rect 101846 311498 101888 311734
rect 101568 311476 101888 311498
rect 101568 308454 101888 308476
rect 101568 308218 101610 308454
rect 101846 308218 101888 308454
rect 101568 308134 101888 308218
rect 101568 307898 101610 308134
rect 101846 307898 101888 308134
rect 101568 307876 101888 307898
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 86208 294054 86528 294076
rect 86208 293818 86250 294054
rect 86486 293818 86528 294054
rect 86208 293734 86528 293818
rect 86208 293498 86250 293734
rect 86486 293498 86528 293734
rect 86208 293476 86528 293498
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 86208 290454 86528 290476
rect 86208 290218 86250 290454
rect 86486 290218 86528 290454
rect 86208 290134 86528 290218
rect 86208 289898 86250 290134
rect 86486 289898 86528 290134
rect 86208 289876 86528 289898
rect 101568 276054 101888 276076
rect 101568 275818 101610 276054
rect 101846 275818 101888 276054
rect 101568 275734 101888 275818
rect 101568 275498 101610 275734
rect 101846 275498 101888 275734
rect 101568 275476 101888 275498
rect 101568 272454 101888 272476
rect 101568 272218 101610 272454
rect 101846 272218 101888 272454
rect 101568 272134 101888 272218
rect 101568 271898 101610 272134
rect 101846 271898 101888 272134
rect 101568 271876 101888 271898
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 86208 258054 86528 258076
rect 86208 257818 86250 258054
rect 86486 257818 86528 258054
rect 86208 257734 86528 257818
rect 86208 257498 86250 257734
rect 86486 257498 86528 257734
rect 86208 257476 86528 257498
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 86208 254454 86528 254476
rect 86208 254218 86250 254454
rect 86486 254218 86528 254454
rect 86208 254134 86528 254218
rect 86208 253898 86250 254134
rect 86486 253898 86528 254134
rect 86208 253876 86528 253898
rect 101568 240054 101888 240076
rect 101568 239818 101610 240054
rect 101846 239818 101888 240054
rect 101568 239734 101888 239818
rect 101568 239498 101610 239734
rect 101846 239498 101888 239734
rect 101568 239476 101888 239498
rect 101568 236454 101888 236476
rect 101568 236218 101610 236454
rect 101846 236218 101888 236454
rect 101568 236134 101888 236218
rect 101568 235898 101610 236134
rect 101846 235898 101888 236134
rect 101568 235876 101888 235898
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 86208 222054 86528 222076
rect 86208 221818 86250 222054
rect 86486 221818 86528 222054
rect 86208 221734 86528 221818
rect 86208 221498 86250 221734
rect 86486 221498 86528 221734
rect 86208 221476 86528 221498
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 86208 218454 86528 218476
rect 86208 218218 86250 218454
rect 86486 218218 86528 218454
rect 86208 218134 86528 218218
rect 86208 217898 86250 218134
rect 86486 217898 86528 218134
rect 86208 217876 86528 217898
rect 101568 204054 101888 204076
rect 101568 203818 101610 204054
rect 101846 203818 101888 204054
rect 101568 203734 101888 203818
rect 101568 203498 101610 203734
rect 101846 203498 101888 203734
rect 101568 203476 101888 203498
rect 101568 200454 101888 200476
rect 101568 200218 101610 200454
rect 101846 200218 101888 200454
rect 101568 200134 101888 200218
rect 101568 199898 101610 200134
rect 101846 199898 101888 200134
rect 101568 199876 101888 199898
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 86208 186054 86528 186076
rect 86208 185818 86250 186054
rect 86486 185818 86528 186054
rect 86208 185734 86528 185818
rect 86208 185498 86250 185734
rect 86486 185498 86528 185734
rect 86208 185476 86528 185498
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 86208 182454 86528 182476
rect 86208 182218 86250 182454
rect 86486 182218 86528 182454
rect 86208 182134 86528 182218
rect 86208 181898 86250 182134
rect 86486 181898 86528 182134
rect 86208 181876 86528 181898
rect 101568 168054 101888 168076
rect 101568 167818 101610 168054
rect 101846 167818 101888 168054
rect 101568 167734 101888 167818
rect 101568 167498 101610 167734
rect 101846 167498 101888 167734
rect 101568 167476 101888 167498
rect 101568 164454 101888 164476
rect 101568 164218 101610 164454
rect 101846 164218 101888 164454
rect 101568 164134 101888 164218
rect 101568 163898 101610 164134
rect 101846 163898 101888 164134
rect 101568 163876 101888 163898
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 86208 150054 86528 150076
rect 86208 149818 86250 150054
rect 86486 149818 86528 150054
rect 86208 149734 86528 149818
rect 86208 149498 86250 149734
rect 86486 149498 86528 149734
rect 86208 149476 86528 149498
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 86208 146454 86528 146476
rect 86208 146218 86250 146454
rect 86486 146218 86528 146454
rect 86208 146134 86528 146218
rect 86208 145898 86250 146134
rect 86486 145898 86528 146134
rect 86208 145876 86528 145898
rect 101568 132054 101888 132076
rect 101568 131818 101610 132054
rect 101846 131818 101888 132054
rect 101568 131734 101888 131818
rect 101568 131498 101610 131734
rect 101846 131498 101888 131734
rect 101568 131476 101888 131498
rect 101568 128454 101888 128476
rect 101568 128218 101610 128454
rect 101846 128218 101888 128454
rect 101568 128134 101888 128218
rect 101568 127898 101610 128134
rect 101846 127898 101888 128134
rect 101568 127876 101888 127898
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 86208 114054 86528 114076
rect 86208 113818 86250 114054
rect 86486 113818 86528 114054
rect 86208 113734 86528 113818
rect 86208 113498 86250 113734
rect 86486 113498 86528 113734
rect 86208 113476 86528 113498
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 86208 110454 86528 110476
rect 86208 110218 86250 110454
rect 86486 110218 86528 110454
rect 86208 110134 86528 110218
rect 86208 109898 86250 110134
rect 86486 109898 86528 110134
rect 86208 109876 86528 109898
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 58404 -3462 58586 -3226
rect 58822 -3462 59004 -3226
rect 58404 -3546 59004 -3462
rect 58404 -3782 58586 -3546
rect 58822 -3782 59004 -3546
rect 58404 -3804 59004 -3782
rect 76404 -2266 77004 5498
rect 90804 92454 91404 102000
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1306 91404 19898
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1884 91404 -1862
rect 94404 96054 95004 102000
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 96291 80748 96357 80749
rect 96291 80684 96292 80748
rect 96356 80684 96357 80748
rect 96291 80683 96357 80684
rect 96294 67829 96354 80683
rect 108804 74454 109404 102000
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 96291 67828 96357 67829
rect 96291 67764 96292 67828
rect 96356 67764 96357 67828
rect 96291 67763 96357 67764
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 76404 -2502 76586 -2266
rect 76822 -2502 77004 -2266
rect 76404 -2586 77004 -2502
rect 76404 -2822 76586 -2586
rect 76822 -2822 77004 -2586
rect 76404 -3804 77004 -2822
rect 94404 -3226 95004 23498
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1884 109404 -902
rect 112404 78054 113004 102000
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 94404 -3462 94586 -3226
rect 94822 -3462 95004 -3226
rect 94404 -3546 95004 -3462
rect 94404 -3782 94586 -3546
rect 94822 -3782 95004 -3546
rect 94404 -3804 95004 -3782
rect 112404 -2266 113004 5498
rect 126804 92454 127404 102000
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1306 127404 19898
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1884 127404 -1862
rect 130404 96054 131004 102000
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 112404 -2502 112586 -2266
rect 112822 -2502 113004 -2266
rect 112404 -2586 113004 -2502
rect 112404 -2822 112586 -2586
rect 112822 -2822 113004 -2586
rect 112404 -3804 113004 -2822
rect 130404 -3226 131004 23498
rect 144804 74454 145404 102000
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1884 145404 -902
rect 148404 78054 149004 102000
rect 162804 92454 163404 102000
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 151491 80204 151557 80205
rect 151491 80140 151492 80204
rect 151556 80140 151557 80204
rect 151491 80139 151557 80140
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 151494 77349 151554 80139
rect 151491 77348 151557 77349
rect 151491 77284 151492 77348
rect 151556 77284 151557 77348
rect 151491 77283 151557 77284
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 130404 -3462 130586 -3226
rect 130822 -3462 131004 -3226
rect 130404 -3546 131004 -3462
rect 130404 -3782 130586 -3546
rect 130822 -3782 131004 -3546
rect 130404 -3804 131004 -3782
rect 148404 -2266 149004 5498
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1306 163404 19898
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1884 163404 -1862
rect 166404 96054 167004 102000
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 148404 -2502 148586 -2266
rect 148822 -2502 149004 -2266
rect 148404 -2586 149004 -2502
rect 148404 -2822 148586 -2586
rect 148822 -2822 149004 -2586
rect 148404 -3804 149004 -2822
rect 166404 -3226 167004 23498
rect 180804 74454 181404 102000
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1884 181404 -902
rect 184404 78054 185004 102000
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 166404 -3462 166586 -3226
rect 166822 -3462 167004 -3226
rect 166404 -3546 167004 -3462
rect 166404 -3782 166586 -3546
rect 166822 -3782 167004 -3546
rect 166404 -3804 167004 -3782
rect 184404 -2266 185004 5498
rect 198804 92454 199404 102000
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1306 199404 19898
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1884 199404 -1862
rect 202404 96054 203004 102000
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 216804 74454 217404 102000
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 215155 60756 215221 60757
rect 215155 60692 215156 60756
rect 215220 60692 215221 60756
rect 215155 60691 215221 60692
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 215158 48381 215218 60691
rect 215155 48380 215221 48381
rect 215155 48316 215156 48380
rect 215220 48316 215221 48380
rect 215155 48315 215221 48316
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 184404 -2502 184586 -2266
rect 184822 -2502 185004 -2266
rect 184404 -2586 185004 -2502
rect 184404 -2822 184586 -2586
rect 184822 -2822 185004 -2586
rect 184404 -3804 185004 -2822
rect 202404 -3226 203004 23498
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1884 217404 -902
rect 220404 78054 221004 102000
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 234804 92454 235404 102000
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 227483 61436 227549 61437
rect 227483 61372 227484 61436
rect 227548 61372 227549 61436
rect 227483 61371 227549 61372
rect 227486 48381 227546 61371
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 227483 48380 227549 48381
rect 227483 48316 227484 48380
rect 227548 48316 227549 48380
rect 227483 48315 227549 48316
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 202404 -3462 202586 -3226
rect 202822 -3462 203004 -3226
rect 202404 -3546 203004 -3462
rect 202404 -3782 202586 -3546
rect 202822 -3782 203004 -3546
rect 202404 -3804 203004 -3782
rect 220404 -2266 221004 5498
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1306 235404 19898
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1884 235404 -1862
rect 238404 96054 239004 102000
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 220404 -2502 220586 -2266
rect 220822 -2502 221004 -2266
rect 220404 -2586 221004 -2502
rect 220404 -2822 220586 -2586
rect 220822 -2822 221004 -2586
rect 220404 -3804 221004 -2822
rect 238404 -3226 239004 23498
rect 252804 74454 253404 102000
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1884 253404 -902
rect 256404 78054 257004 102000
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 238404 -3462 238586 -3226
rect 238822 -3462 239004 -3226
rect 238404 -3546 239004 -3462
rect 238404 -3782 238586 -3546
rect 238822 -3782 239004 -3546
rect 238404 -3804 239004 -3782
rect 256404 -2266 257004 5498
rect 270804 92454 271404 102000
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1306 271404 19898
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1884 271404 -1862
rect 274404 96054 275004 102000
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 256404 -2502 256586 -2266
rect 256822 -2502 257004 -2266
rect 256404 -2586 257004 -2502
rect 256404 -2822 256586 -2586
rect 256822 -2822 257004 -2586
rect 256404 -3804 257004 -2822
rect 274404 -3226 275004 23498
rect 288804 74454 289404 102000
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1884 289404 -902
rect 292404 78054 293004 102000
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 274404 -3462 274586 -3226
rect 274822 -3462 275004 -3226
rect 274404 -3546 275004 -3462
rect 274404 -3782 274586 -3546
rect 274822 -3782 275004 -3546
rect 274404 -3804 275004 -3782
rect 292404 -2266 293004 5498
rect 306804 92454 307404 102000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1306 307404 19898
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1884 307404 -1862
rect 310404 96054 311004 102000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 292404 -2502 292586 -2266
rect 292822 -2502 293004 -2266
rect 292404 -2586 293004 -2502
rect 292404 -2822 292586 -2586
rect 292822 -2822 293004 -2586
rect 292404 -3804 293004 -2822
rect 310404 -3226 311004 23498
rect 324804 74454 325404 102000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1884 325404 -902
rect 328404 78054 329004 102000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 310404 -3462 310586 -3226
rect 310822 -3462 311004 -3226
rect 310404 -3546 311004 -3462
rect 310404 -3782 310586 -3546
rect 310822 -3782 311004 -3546
rect 310404 -3804 311004 -3782
rect 328404 -2266 329004 5498
rect 342804 92454 343404 102000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1306 343404 19898
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1884 343404 -1862
rect 346404 96054 347004 102000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 328404 -2502 328586 -2266
rect 328822 -2502 329004 -2266
rect 328404 -2586 329004 -2502
rect 328404 -2822 328586 -2586
rect 328822 -2822 329004 -2586
rect 328404 -3804 329004 -2822
rect 346404 -3226 347004 23498
rect 360804 74454 361404 102000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1884 361404 -902
rect 364404 78054 365004 102000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 346404 -3462 346586 -3226
rect 346822 -3462 347004 -3226
rect 346404 -3546 347004 -3462
rect 346404 -3782 346586 -3546
rect 346822 -3782 347004 -3546
rect 346404 -3804 347004 -3782
rect 364404 -2266 365004 5498
rect 378804 92454 379404 102000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1306 379404 19898
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1884 379404 -1862
rect 382404 96054 383004 102000
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 364404 -2502 364586 -2266
rect 364822 -2502 365004 -2266
rect 364404 -2586 365004 -2502
rect 364404 -2822 364586 -2586
rect 364822 -2822 365004 -2586
rect 364404 -3804 365004 -2822
rect 382404 -3226 383004 23498
rect 396804 74454 397404 102000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1884 397404 -902
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 382404 -3462 382586 -3226
rect 382822 -3462 383004 -3226
rect 382404 -3546 383004 -3462
rect 382404 -3782 382586 -3546
rect 382822 -3782 383004 -3546
rect 382404 -3804 383004 -3782
rect 400404 -2266 401004 5498
rect 414804 705798 415404 705820
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668454 415404 705242
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1306 415404 19898
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1884 415404 -1862
rect 418404 672054 419004 707162
rect 436404 706758 437004 707740
rect 436404 706522 436586 706758
rect 436822 706522 437004 706758
rect 436404 706438 437004 706522
rect 436404 706202 436586 706438
rect 436822 706202 437004 706438
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 400404 -2502 400586 -2266
rect 400822 -2502 401004 -2266
rect 400404 -2586 401004 -2502
rect 400404 -2822 400586 -2586
rect 400822 -2822 401004 -2586
rect 400404 -3804 401004 -2822
rect 418404 -3226 419004 23498
rect 432804 704838 433404 705820
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1884 433404 -902
rect 436404 690054 437004 706202
rect 454404 707718 455004 707740
rect 454404 707482 454586 707718
rect 454822 707482 455004 707718
rect 454404 707398 455004 707482
rect 454404 707162 454586 707398
rect 454822 707162 455004 707398
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 418404 -3462 418586 -3226
rect 418822 -3462 419004 -3226
rect 418404 -3546 419004 -3462
rect 418404 -3782 418586 -3546
rect 418822 -3782 419004 -3546
rect 418404 -3804 419004 -3782
rect 436404 -2266 437004 5498
rect 450804 705798 451404 705820
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668454 451404 705242
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1306 451404 19898
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1884 451404 -1862
rect 454404 672054 455004 707162
rect 472404 706758 473004 707740
rect 472404 706522 472586 706758
rect 472822 706522 473004 706758
rect 472404 706438 473004 706522
rect 472404 706202 472586 706438
rect 472822 706202 473004 706438
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 436404 -2502 436586 -2266
rect 436822 -2502 437004 -2266
rect 436404 -2586 437004 -2502
rect 436404 -2822 436586 -2586
rect 436822 -2822 437004 -2586
rect 436404 -3804 437004 -2822
rect 454404 -3226 455004 23498
rect 468804 704838 469404 705820
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1884 469404 -902
rect 472404 690054 473004 706202
rect 490404 707718 491004 707740
rect 490404 707482 490586 707718
rect 490822 707482 491004 707718
rect 490404 707398 491004 707482
rect 490404 707162 490586 707398
rect 490822 707162 491004 707398
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 454404 -3462 454586 -3226
rect 454822 -3462 455004 -3226
rect 454404 -3546 455004 -3462
rect 454404 -3782 454586 -3546
rect 454822 -3782 455004 -3546
rect 454404 -3804 455004 -3782
rect 472404 -2266 473004 5498
rect 486804 705798 487404 705820
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668454 487404 705242
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1306 487404 19898
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1884 487404 -1862
rect 490404 672054 491004 707162
rect 508404 706758 509004 707740
rect 508404 706522 508586 706758
rect 508822 706522 509004 706758
rect 508404 706438 509004 706522
rect 508404 706202 508586 706438
rect 508822 706202 509004 706438
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 472404 -2502 472586 -2266
rect 472822 -2502 473004 -2266
rect 472404 -2586 473004 -2502
rect 472404 -2822 472586 -2586
rect 472822 -2822 473004 -2586
rect 472404 -3804 473004 -2822
rect 490404 -3226 491004 23498
rect 504804 704838 505404 705820
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1884 505404 -902
rect 508404 690054 509004 706202
rect 526404 707718 527004 707740
rect 526404 707482 526586 707718
rect 526822 707482 527004 707718
rect 526404 707398 527004 707482
rect 526404 707162 526586 707398
rect 526822 707162 527004 707398
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 490404 -3462 490586 -3226
rect 490822 -3462 491004 -3226
rect 490404 -3546 491004 -3462
rect 490404 -3782 490586 -3546
rect 490822 -3782 491004 -3546
rect 490404 -3804 491004 -3782
rect 508404 -2266 509004 5498
rect 522804 705798 523404 705820
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668454 523404 705242
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1306 523404 19898
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1884 523404 -1862
rect 526404 672054 527004 707162
rect 544404 706758 545004 707740
rect 544404 706522 544586 706758
rect 544822 706522 545004 706758
rect 544404 706438 545004 706522
rect 544404 706202 544586 706438
rect 544822 706202 545004 706438
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 508404 -2502 508586 -2266
rect 508822 -2502 509004 -2266
rect 508404 -2586 509004 -2502
rect 508404 -2822 508586 -2586
rect 508822 -2822 509004 -2586
rect 508404 -3804 509004 -2822
rect 526404 -3226 527004 23498
rect 540804 704838 541404 705820
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1884 541404 -902
rect 544404 690054 545004 706202
rect 562404 707718 563004 707740
rect 562404 707482 562586 707718
rect 562822 707482 563004 707718
rect 562404 707398 563004 707482
rect 562404 707162 562586 707398
rect 562822 707162 563004 707398
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 526404 -3462 526586 -3226
rect 526822 -3462 527004 -3226
rect 526404 -3546 527004 -3462
rect 526404 -3782 526586 -3546
rect 526822 -3782 527004 -3546
rect 526404 -3804 527004 -3782
rect 544404 -2266 545004 5498
rect 558804 705798 559404 705820
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668454 559404 705242
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1306 559404 19898
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1884 559404 -1862
rect 562404 672054 563004 707162
rect 580404 706758 581004 707740
rect 588200 707718 588800 707740
rect 588200 707482 588382 707718
rect 588618 707482 588800 707718
rect 588200 707398 588800 707482
rect 588200 707162 588382 707398
rect 588618 707162 588800 707398
rect 580404 706522 580586 706758
rect 580822 706522 581004 706758
rect 580404 706438 581004 706522
rect 580404 706202 580586 706438
rect 580822 706202 581004 706438
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 544404 -2502 544586 -2266
rect 544822 -2502 545004 -2266
rect 544404 -2586 545004 -2502
rect 544404 -2822 544586 -2586
rect 544822 -2822 545004 -2586
rect 544404 -3804 545004 -2822
rect 562404 -3226 563004 23498
rect 576804 704838 577404 705820
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1884 577404 -902
rect 580404 690054 581004 706202
rect 587240 706758 587840 706780
rect 587240 706522 587422 706758
rect 587658 706522 587840 706758
rect 587240 706438 587840 706522
rect 587240 706202 587422 706438
rect 587658 706202 587840 706438
rect 586280 705798 586880 705820
rect 586280 705562 586462 705798
rect 586698 705562 586880 705798
rect 586280 705478 586880 705562
rect 586280 705242 586462 705478
rect 586698 705242 586880 705478
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 562404 -3462 562586 -3226
rect 562822 -3462 563004 -3226
rect 562404 -3546 563004 -3462
rect 562404 -3782 562586 -3546
rect 562822 -3782 563004 -3546
rect 562404 -3804 563004 -3782
rect 580404 -2266 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586280 668454 586880 705242
rect 586280 668218 586462 668454
rect 586698 668218 586880 668454
rect 586280 668134 586880 668218
rect 586280 667898 586462 668134
rect 586698 667898 586880 668134
rect 586280 632454 586880 667898
rect 586280 632218 586462 632454
rect 586698 632218 586880 632454
rect 586280 632134 586880 632218
rect 586280 631898 586462 632134
rect 586698 631898 586880 632134
rect 586280 596454 586880 631898
rect 586280 596218 586462 596454
rect 586698 596218 586880 596454
rect 586280 596134 586880 596218
rect 586280 595898 586462 596134
rect 586698 595898 586880 596134
rect 586280 560454 586880 595898
rect 586280 560218 586462 560454
rect 586698 560218 586880 560454
rect 586280 560134 586880 560218
rect 586280 559898 586462 560134
rect 586698 559898 586880 560134
rect 586280 524454 586880 559898
rect 586280 524218 586462 524454
rect 586698 524218 586880 524454
rect 586280 524134 586880 524218
rect 586280 523898 586462 524134
rect 586698 523898 586880 524134
rect 586280 488454 586880 523898
rect 586280 488218 586462 488454
rect 586698 488218 586880 488454
rect 586280 488134 586880 488218
rect 586280 487898 586462 488134
rect 586698 487898 586880 488134
rect 586280 452454 586880 487898
rect 586280 452218 586462 452454
rect 586698 452218 586880 452454
rect 586280 452134 586880 452218
rect 586280 451898 586462 452134
rect 586698 451898 586880 452134
rect 586280 416454 586880 451898
rect 586280 416218 586462 416454
rect 586698 416218 586880 416454
rect 586280 416134 586880 416218
rect 586280 415898 586462 416134
rect 586698 415898 586880 416134
rect 586280 380454 586880 415898
rect 586280 380218 586462 380454
rect 586698 380218 586880 380454
rect 586280 380134 586880 380218
rect 586280 379898 586462 380134
rect 586698 379898 586880 380134
rect 586280 344454 586880 379898
rect 586280 344218 586462 344454
rect 586698 344218 586880 344454
rect 586280 344134 586880 344218
rect 586280 343898 586462 344134
rect 586698 343898 586880 344134
rect 586280 308454 586880 343898
rect 586280 308218 586462 308454
rect 586698 308218 586880 308454
rect 586280 308134 586880 308218
rect 586280 307898 586462 308134
rect 586698 307898 586880 308134
rect 586280 272454 586880 307898
rect 586280 272218 586462 272454
rect 586698 272218 586880 272454
rect 586280 272134 586880 272218
rect 586280 271898 586462 272134
rect 586698 271898 586880 272134
rect 586280 236454 586880 271898
rect 586280 236218 586462 236454
rect 586698 236218 586880 236454
rect 586280 236134 586880 236218
rect 586280 235898 586462 236134
rect 586698 235898 586880 236134
rect 586280 200454 586880 235898
rect 586280 200218 586462 200454
rect 586698 200218 586880 200454
rect 586280 200134 586880 200218
rect 586280 199898 586462 200134
rect 586698 199898 586880 200134
rect 586280 164454 586880 199898
rect 586280 164218 586462 164454
rect 586698 164218 586880 164454
rect 586280 164134 586880 164218
rect 586280 163898 586462 164134
rect 586698 163898 586880 164134
rect 586280 128454 586880 163898
rect 586280 128218 586462 128454
rect 586698 128218 586880 128454
rect 586280 128134 586880 128218
rect 586280 127898 586462 128134
rect 586698 127898 586880 128134
rect 586280 92454 586880 127898
rect 586280 92218 586462 92454
rect 586698 92218 586880 92454
rect 586280 92134 586880 92218
rect 586280 91898 586462 92134
rect 586698 91898 586880 92134
rect 586280 56454 586880 91898
rect 586280 56218 586462 56454
rect 586698 56218 586880 56454
rect 586280 56134 586880 56218
rect 586280 55898 586462 56134
rect 586698 55898 586880 56134
rect 586280 20454 586880 55898
rect 586280 20218 586462 20454
rect 586698 20218 586880 20454
rect 586280 20134 586880 20218
rect 586280 19898 586462 20134
rect 586698 19898 586880 20134
rect 586280 -1306 586880 19898
rect 586280 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect 586280 -1626 586880 -1542
rect 586280 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect 586280 -1884 586880 -1862
rect 587240 690054 587840 706202
rect 587240 689818 587422 690054
rect 587658 689818 587840 690054
rect 587240 689734 587840 689818
rect 587240 689498 587422 689734
rect 587658 689498 587840 689734
rect 587240 654054 587840 689498
rect 587240 653818 587422 654054
rect 587658 653818 587840 654054
rect 587240 653734 587840 653818
rect 587240 653498 587422 653734
rect 587658 653498 587840 653734
rect 587240 618054 587840 653498
rect 587240 617818 587422 618054
rect 587658 617818 587840 618054
rect 587240 617734 587840 617818
rect 587240 617498 587422 617734
rect 587658 617498 587840 617734
rect 587240 582054 587840 617498
rect 587240 581818 587422 582054
rect 587658 581818 587840 582054
rect 587240 581734 587840 581818
rect 587240 581498 587422 581734
rect 587658 581498 587840 581734
rect 587240 546054 587840 581498
rect 587240 545818 587422 546054
rect 587658 545818 587840 546054
rect 587240 545734 587840 545818
rect 587240 545498 587422 545734
rect 587658 545498 587840 545734
rect 587240 510054 587840 545498
rect 587240 509818 587422 510054
rect 587658 509818 587840 510054
rect 587240 509734 587840 509818
rect 587240 509498 587422 509734
rect 587658 509498 587840 509734
rect 587240 474054 587840 509498
rect 587240 473818 587422 474054
rect 587658 473818 587840 474054
rect 587240 473734 587840 473818
rect 587240 473498 587422 473734
rect 587658 473498 587840 473734
rect 587240 438054 587840 473498
rect 587240 437818 587422 438054
rect 587658 437818 587840 438054
rect 587240 437734 587840 437818
rect 587240 437498 587422 437734
rect 587658 437498 587840 437734
rect 587240 402054 587840 437498
rect 587240 401818 587422 402054
rect 587658 401818 587840 402054
rect 587240 401734 587840 401818
rect 587240 401498 587422 401734
rect 587658 401498 587840 401734
rect 587240 366054 587840 401498
rect 587240 365818 587422 366054
rect 587658 365818 587840 366054
rect 587240 365734 587840 365818
rect 587240 365498 587422 365734
rect 587658 365498 587840 365734
rect 587240 330054 587840 365498
rect 587240 329818 587422 330054
rect 587658 329818 587840 330054
rect 587240 329734 587840 329818
rect 587240 329498 587422 329734
rect 587658 329498 587840 329734
rect 587240 294054 587840 329498
rect 587240 293818 587422 294054
rect 587658 293818 587840 294054
rect 587240 293734 587840 293818
rect 587240 293498 587422 293734
rect 587658 293498 587840 293734
rect 587240 258054 587840 293498
rect 587240 257818 587422 258054
rect 587658 257818 587840 258054
rect 587240 257734 587840 257818
rect 587240 257498 587422 257734
rect 587658 257498 587840 257734
rect 587240 222054 587840 257498
rect 587240 221818 587422 222054
rect 587658 221818 587840 222054
rect 587240 221734 587840 221818
rect 587240 221498 587422 221734
rect 587658 221498 587840 221734
rect 587240 186054 587840 221498
rect 587240 185818 587422 186054
rect 587658 185818 587840 186054
rect 587240 185734 587840 185818
rect 587240 185498 587422 185734
rect 587658 185498 587840 185734
rect 587240 150054 587840 185498
rect 587240 149818 587422 150054
rect 587658 149818 587840 150054
rect 587240 149734 587840 149818
rect 587240 149498 587422 149734
rect 587658 149498 587840 149734
rect 587240 114054 587840 149498
rect 587240 113818 587422 114054
rect 587658 113818 587840 114054
rect 587240 113734 587840 113818
rect 587240 113498 587422 113734
rect 587658 113498 587840 113734
rect 587240 78054 587840 113498
rect 587240 77818 587422 78054
rect 587658 77818 587840 78054
rect 587240 77734 587840 77818
rect 587240 77498 587422 77734
rect 587658 77498 587840 77734
rect 587240 42054 587840 77498
rect 587240 41818 587422 42054
rect 587658 41818 587840 42054
rect 587240 41734 587840 41818
rect 587240 41498 587422 41734
rect 587658 41498 587840 41734
rect 587240 6054 587840 41498
rect 587240 5818 587422 6054
rect 587658 5818 587840 6054
rect 587240 5734 587840 5818
rect 587240 5498 587422 5734
rect 587658 5498 587840 5734
rect 580404 -2502 580586 -2266
rect 580822 -2502 581004 -2266
rect 580404 -2586 581004 -2502
rect 580404 -2822 580586 -2586
rect 580822 -2822 581004 -2586
rect 580404 -3804 581004 -2822
rect 587240 -2266 587840 5498
rect 587240 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect 587240 -2586 587840 -2502
rect 587240 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect 587240 -2844 587840 -2822
rect 588200 672054 588800 707162
rect 588200 671818 588382 672054
rect 588618 671818 588800 672054
rect 588200 671734 588800 671818
rect 588200 671498 588382 671734
rect 588618 671498 588800 671734
rect 588200 636054 588800 671498
rect 588200 635818 588382 636054
rect 588618 635818 588800 636054
rect 588200 635734 588800 635818
rect 588200 635498 588382 635734
rect 588618 635498 588800 635734
rect 588200 600054 588800 635498
rect 588200 599818 588382 600054
rect 588618 599818 588800 600054
rect 588200 599734 588800 599818
rect 588200 599498 588382 599734
rect 588618 599498 588800 599734
rect 588200 564054 588800 599498
rect 588200 563818 588382 564054
rect 588618 563818 588800 564054
rect 588200 563734 588800 563818
rect 588200 563498 588382 563734
rect 588618 563498 588800 563734
rect 588200 528054 588800 563498
rect 588200 527818 588382 528054
rect 588618 527818 588800 528054
rect 588200 527734 588800 527818
rect 588200 527498 588382 527734
rect 588618 527498 588800 527734
rect 588200 492054 588800 527498
rect 588200 491818 588382 492054
rect 588618 491818 588800 492054
rect 588200 491734 588800 491818
rect 588200 491498 588382 491734
rect 588618 491498 588800 491734
rect 588200 456054 588800 491498
rect 588200 455818 588382 456054
rect 588618 455818 588800 456054
rect 588200 455734 588800 455818
rect 588200 455498 588382 455734
rect 588618 455498 588800 455734
rect 588200 420054 588800 455498
rect 588200 419818 588382 420054
rect 588618 419818 588800 420054
rect 588200 419734 588800 419818
rect 588200 419498 588382 419734
rect 588618 419498 588800 419734
rect 588200 384054 588800 419498
rect 588200 383818 588382 384054
rect 588618 383818 588800 384054
rect 588200 383734 588800 383818
rect 588200 383498 588382 383734
rect 588618 383498 588800 383734
rect 588200 348054 588800 383498
rect 588200 347818 588382 348054
rect 588618 347818 588800 348054
rect 588200 347734 588800 347818
rect 588200 347498 588382 347734
rect 588618 347498 588800 347734
rect 588200 312054 588800 347498
rect 588200 311818 588382 312054
rect 588618 311818 588800 312054
rect 588200 311734 588800 311818
rect 588200 311498 588382 311734
rect 588618 311498 588800 311734
rect 588200 276054 588800 311498
rect 588200 275818 588382 276054
rect 588618 275818 588800 276054
rect 588200 275734 588800 275818
rect 588200 275498 588382 275734
rect 588618 275498 588800 275734
rect 588200 240054 588800 275498
rect 588200 239818 588382 240054
rect 588618 239818 588800 240054
rect 588200 239734 588800 239818
rect 588200 239498 588382 239734
rect 588618 239498 588800 239734
rect 588200 204054 588800 239498
rect 588200 203818 588382 204054
rect 588618 203818 588800 204054
rect 588200 203734 588800 203818
rect 588200 203498 588382 203734
rect 588618 203498 588800 203734
rect 588200 168054 588800 203498
rect 588200 167818 588382 168054
rect 588618 167818 588800 168054
rect 588200 167734 588800 167818
rect 588200 167498 588382 167734
rect 588618 167498 588800 167734
rect 588200 132054 588800 167498
rect 588200 131818 588382 132054
rect 588618 131818 588800 132054
rect 588200 131734 588800 131818
rect 588200 131498 588382 131734
rect 588618 131498 588800 131734
rect 588200 96054 588800 131498
rect 588200 95818 588382 96054
rect 588618 95818 588800 96054
rect 588200 95734 588800 95818
rect 588200 95498 588382 95734
rect 588618 95498 588800 95734
rect 588200 60054 588800 95498
rect 588200 59818 588382 60054
rect 588618 59818 588800 60054
rect 588200 59734 588800 59818
rect 588200 59498 588382 59734
rect 588618 59498 588800 59734
rect 588200 24054 588800 59498
rect 588200 23818 588382 24054
rect 588618 23818 588800 24054
rect 588200 23734 588800 23818
rect 588200 23498 588382 23734
rect 588618 23498 588800 23734
rect 588200 -3226 588800 23498
rect 588200 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect 588200 -3546 588800 -3462
rect 588200 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect 588200 -3804 588800 -3782
<< via4 >>
rect -4694 707482 -4458 707718
rect -4694 707162 -4458 707398
rect -4694 671818 -4458 672054
rect -4694 671498 -4458 671734
rect -4694 635818 -4458 636054
rect -4694 635498 -4458 635734
rect -4694 599818 -4458 600054
rect -4694 599498 -4458 599734
rect -4694 563818 -4458 564054
rect -4694 563498 -4458 563734
rect -4694 527818 -4458 528054
rect -4694 527498 -4458 527734
rect -4694 491818 -4458 492054
rect -4694 491498 -4458 491734
rect -4694 455818 -4458 456054
rect -4694 455498 -4458 455734
rect -4694 419818 -4458 420054
rect -4694 419498 -4458 419734
rect -4694 383818 -4458 384054
rect -4694 383498 -4458 383734
rect -4694 347818 -4458 348054
rect -4694 347498 -4458 347734
rect -4694 311818 -4458 312054
rect -4694 311498 -4458 311734
rect -4694 275818 -4458 276054
rect -4694 275498 -4458 275734
rect -4694 239818 -4458 240054
rect -4694 239498 -4458 239734
rect -4694 203818 -4458 204054
rect -4694 203498 -4458 203734
rect -4694 167818 -4458 168054
rect -4694 167498 -4458 167734
rect -4694 131818 -4458 132054
rect -4694 131498 -4458 131734
rect -4694 95818 -4458 96054
rect -4694 95498 -4458 95734
rect -4694 59818 -4458 60054
rect -4694 59498 -4458 59734
rect -4694 23818 -4458 24054
rect -4694 23498 -4458 23734
rect -3734 706522 -3498 706758
rect -3734 706202 -3498 706438
rect 4586 706522 4822 706758
rect 4586 706202 4822 706438
rect -3734 689818 -3498 690054
rect -3734 689498 -3498 689734
rect -3734 653818 -3498 654054
rect -3734 653498 -3498 653734
rect -3734 617818 -3498 618054
rect -3734 617498 -3498 617734
rect -3734 581818 -3498 582054
rect -3734 581498 -3498 581734
rect -3734 545818 -3498 546054
rect -3734 545498 -3498 545734
rect -3734 509818 -3498 510054
rect -3734 509498 -3498 509734
rect -3734 473818 -3498 474054
rect -3734 473498 -3498 473734
rect -3734 437818 -3498 438054
rect -3734 437498 -3498 437734
rect -3734 401818 -3498 402054
rect -3734 401498 -3498 401734
rect -3734 365818 -3498 366054
rect -3734 365498 -3498 365734
rect -3734 329818 -3498 330054
rect -3734 329498 -3498 329734
rect -3734 293818 -3498 294054
rect -3734 293498 -3498 293734
rect -3734 257818 -3498 258054
rect -3734 257498 -3498 257734
rect -3734 221818 -3498 222054
rect -3734 221498 -3498 221734
rect -3734 185818 -3498 186054
rect -3734 185498 -3498 185734
rect -3734 149818 -3498 150054
rect -3734 149498 -3498 149734
rect -3734 113818 -3498 114054
rect -3734 113498 -3498 113734
rect -3734 77818 -3498 78054
rect -3734 77498 -3498 77734
rect -3734 41818 -3498 42054
rect -3734 41498 -3498 41734
rect -3734 5818 -3498 6054
rect -3734 5498 -3498 5734
rect -2774 705562 -2538 705798
rect -2774 705242 -2538 705478
rect -2774 668218 -2538 668454
rect -2774 667898 -2538 668134
rect -2774 632218 -2538 632454
rect -2774 631898 -2538 632134
rect -2774 596218 -2538 596454
rect -2774 595898 -2538 596134
rect -2774 560218 -2538 560454
rect -2774 559898 -2538 560134
rect -2774 524218 -2538 524454
rect -2774 523898 -2538 524134
rect -2774 488218 -2538 488454
rect -2774 487898 -2538 488134
rect -2774 452218 -2538 452454
rect -2774 451898 -2538 452134
rect -2774 416218 -2538 416454
rect -2774 415898 -2538 416134
rect -2774 380218 -2538 380454
rect -2774 379898 -2538 380134
rect -2774 344218 -2538 344454
rect -2774 343898 -2538 344134
rect -2774 308218 -2538 308454
rect -2774 307898 -2538 308134
rect -2774 272218 -2538 272454
rect -2774 271898 -2538 272134
rect -2774 236218 -2538 236454
rect -2774 235898 -2538 236134
rect -2774 200218 -2538 200454
rect -2774 199898 -2538 200134
rect -2774 164218 -2538 164454
rect -2774 163898 -2538 164134
rect -2774 128218 -2538 128454
rect -2774 127898 -2538 128134
rect -2774 92218 -2538 92454
rect -2774 91898 -2538 92134
rect -2774 56218 -2538 56454
rect -2774 55898 -2538 56134
rect -2774 20218 -2538 20454
rect -2774 19898 -2538 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2774 -1542 -2538 -1306
rect -2774 -1862 -2538 -1626
rect 22586 707482 22822 707718
rect 22586 707162 22822 707398
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3734 -2502 -3498 -2266
rect -3734 -2822 -3498 -2586
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 40586 706522 40822 706758
rect 40586 706202 40822 706438
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 4586 -2502 4822 -2266
rect 4586 -2822 4822 -2586
rect -4694 -3462 -4458 -3226
rect -4694 -3782 -4458 -3546
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 58586 707482 58822 707718
rect 58586 707162 58822 707398
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 22586 -3462 22822 -3226
rect 22586 -3782 22822 -3546
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 76586 706522 76822 706758
rect 76586 706202 76822 706438
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 40586 -2502 40822 -2266
rect 40586 -2822 40822 -2586
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 94586 707482 94822 707718
rect 94586 707162 94822 707398
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 112586 706522 112822 706758
rect 112586 706202 112822 706438
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 130586 707482 130822 707718
rect 130586 707162 130822 707398
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 148586 706522 148822 706758
rect 148586 706202 148822 706438
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 166586 707482 166822 707718
rect 166586 707162 166822 707398
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 184586 706522 184822 706758
rect 184586 706202 184822 706438
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 202586 707482 202822 707718
rect 202586 707162 202822 707398
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 220586 706522 220822 706758
rect 220586 706202 220822 706438
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 238586 707482 238822 707718
rect 238586 707162 238822 707398
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 256586 706522 256822 706758
rect 256586 706202 256822 706438
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 274586 707482 274822 707718
rect 274586 707162 274822 707398
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 292586 706522 292822 706758
rect 292586 706202 292822 706438
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 310586 707482 310822 707718
rect 310586 707162 310822 707398
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 328586 706522 328822 706758
rect 328586 706202 328822 706438
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 346586 707482 346822 707718
rect 346586 707162 346822 707398
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 364586 706522 364822 706758
rect 364586 706202 364822 706438
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 382586 707482 382822 707718
rect 382586 707162 382822 707398
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 400586 706522 400822 706758
rect 400586 706202 400822 706438
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 418586 707482 418822 707718
rect 418586 707162 418822 707398
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 101610 419818 101846 420054
rect 101610 419498 101846 419734
rect 101610 416218 101846 416454
rect 101610 415898 101846 416134
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 86250 401818 86486 402054
rect 86250 401498 86486 401734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 86250 398218 86486 398454
rect 86250 397898 86486 398134
rect 101610 383818 101846 384054
rect 101610 383498 101846 383734
rect 101610 380218 101846 380454
rect 101610 379898 101846 380134
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 86250 365818 86486 366054
rect 86250 365498 86486 365734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 86250 362218 86486 362454
rect 86250 361898 86486 362134
rect 101610 347818 101846 348054
rect 101610 347498 101846 347734
rect 101610 344218 101846 344454
rect 101610 343898 101846 344134
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 86250 329818 86486 330054
rect 86250 329498 86486 329734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 86250 326218 86486 326454
rect 86250 325898 86486 326134
rect 101610 311818 101846 312054
rect 101610 311498 101846 311734
rect 101610 308218 101846 308454
rect 101610 307898 101846 308134
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 86250 293818 86486 294054
rect 86250 293498 86486 293734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 86250 290218 86486 290454
rect 86250 289898 86486 290134
rect 101610 275818 101846 276054
rect 101610 275498 101846 275734
rect 101610 272218 101846 272454
rect 101610 271898 101846 272134
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 86250 257818 86486 258054
rect 86250 257498 86486 257734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 86250 254218 86486 254454
rect 86250 253898 86486 254134
rect 101610 239818 101846 240054
rect 101610 239498 101846 239734
rect 101610 236218 101846 236454
rect 101610 235898 101846 236134
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 86250 221818 86486 222054
rect 86250 221498 86486 221734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 86250 218218 86486 218454
rect 86250 217898 86486 218134
rect 101610 203818 101846 204054
rect 101610 203498 101846 203734
rect 101610 200218 101846 200454
rect 101610 199898 101846 200134
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 86250 185818 86486 186054
rect 86250 185498 86486 185734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 86250 182218 86486 182454
rect 86250 181898 86486 182134
rect 101610 167818 101846 168054
rect 101610 167498 101846 167734
rect 101610 164218 101846 164454
rect 101610 163898 101846 164134
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 86250 149818 86486 150054
rect 86250 149498 86486 149734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 86250 146218 86486 146454
rect 86250 145898 86486 146134
rect 101610 131818 101846 132054
rect 101610 131498 101846 131734
rect 101610 128218 101846 128454
rect 101610 127898 101846 128134
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 86250 113818 86486 114054
rect 86250 113498 86486 113734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 86250 110218 86486 110454
rect 86250 109898 86486 110134
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 58586 -3462 58822 -3226
rect 58586 -3782 58822 -3546
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 76586 -2502 76822 -2266
rect 76586 -2822 76822 -2586
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 94586 -3462 94822 -3226
rect 94586 -3782 94822 -3546
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 112586 -2502 112822 -2266
rect 112586 -2822 112822 -2586
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 130586 -3462 130822 -3226
rect 130586 -3782 130822 -3546
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 148586 -2502 148822 -2266
rect 148586 -2822 148822 -2586
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 166586 -3462 166822 -3226
rect 166586 -3782 166822 -3546
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 184586 -2502 184822 -2266
rect 184586 -2822 184822 -2586
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 202586 -3462 202822 -3226
rect 202586 -3782 202822 -3546
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 220586 -2502 220822 -2266
rect 220586 -2822 220822 -2586
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 238586 -3462 238822 -3226
rect 238586 -3782 238822 -3546
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 256586 -2502 256822 -2266
rect 256586 -2822 256822 -2586
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 274586 -3462 274822 -3226
rect 274586 -3782 274822 -3546
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 292586 -2502 292822 -2266
rect 292586 -2822 292822 -2586
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 310586 -3462 310822 -3226
rect 310586 -3782 310822 -3546
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 328586 -2502 328822 -2266
rect 328586 -2822 328822 -2586
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 346586 -3462 346822 -3226
rect 346586 -3782 346822 -3546
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 364586 -2502 364822 -2266
rect 364586 -2822 364822 -2586
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 382586 -3462 382822 -3226
rect 382586 -3782 382822 -3546
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 436586 706522 436822 706758
rect 436586 706202 436822 706438
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 400586 -2502 400822 -2266
rect 400586 -2822 400822 -2586
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 454586 707482 454822 707718
rect 454586 707162 454822 707398
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 418586 -3462 418822 -3226
rect 418586 -3782 418822 -3546
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 472586 706522 472822 706758
rect 472586 706202 472822 706438
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 436586 -2502 436822 -2266
rect 436586 -2822 436822 -2586
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 490586 707482 490822 707718
rect 490586 707162 490822 707398
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 454586 -3462 454822 -3226
rect 454586 -3782 454822 -3546
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 508586 706522 508822 706758
rect 508586 706202 508822 706438
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 472586 -2502 472822 -2266
rect 472586 -2822 472822 -2586
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 526586 707482 526822 707718
rect 526586 707162 526822 707398
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 490586 -3462 490822 -3226
rect 490586 -3782 490822 -3546
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 544586 706522 544822 706758
rect 544586 706202 544822 706438
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 508586 -2502 508822 -2266
rect 508586 -2822 508822 -2586
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 562586 707482 562822 707718
rect 562586 707162 562822 707398
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 526586 -3462 526822 -3226
rect 526586 -3782 526822 -3546
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 588382 707482 588618 707718
rect 588382 707162 588618 707398
rect 580586 706522 580822 706758
rect 580586 706202 580822 706438
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 544586 -2502 544822 -2266
rect 544586 -2822 544822 -2586
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587422 706522 587658 706758
rect 587422 706202 587658 706438
rect 586462 705562 586698 705798
rect 586462 705242 586698 705478
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 562586 -3462 562822 -3226
rect 562586 -3782 562822 -3546
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586462 668218 586698 668454
rect 586462 667898 586698 668134
rect 586462 632218 586698 632454
rect 586462 631898 586698 632134
rect 586462 596218 586698 596454
rect 586462 595898 586698 596134
rect 586462 560218 586698 560454
rect 586462 559898 586698 560134
rect 586462 524218 586698 524454
rect 586462 523898 586698 524134
rect 586462 488218 586698 488454
rect 586462 487898 586698 488134
rect 586462 452218 586698 452454
rect 586462 451898 586698 452134
rect 586462 416218 586698 416454
rect 586462 415898 586698 416134
rect 586462 380218 586698 380454
rect 586462 379898 586698 380134
rect 586462 344218 586698 344454
rect 586462 343898 586698 344134
rect 586462 308218 586698 308454
rect 586462 307898 586698 308134
rect 586462 272218 586698 272454
rect 586462 271898 586698 272134
rect 586462 236218 586698 236454
rect 586462 235898 586698 236134
rect 586462 200218 586698 200454
rect 586462 199898 586698 200134
rect 586462 164218 586698 164454
rect 586462 163898 586698 164134
rect 586462 128218 586698 128454
rect 586462 127898 586698 128134
rect 586462 92218 586698 92454
rect 586462 91898 586698 92134
rect 586462 56218 586698 56454
rect 586462 55898 586698 56134
rect 586462 20218 586698 20454
rect 586462 19898 586698 20134
rect 586462 -1542 586698 -1306
rect 586462 -1862 586698 -1626
rect 587422 689818 587658 690054
rect 587422 689498 587658 689734
rect 587422 653818 587658 654054
rect 587422 653498 587658 653734
rect 587422 617818 587658 618054
rect 587422 617498 587658 617734
rect 587422 581818 587658 582054
rect 587422 581498 587658 581734
rect 587422 545818 587658 546054
rect 587422 545498 587658 545734
rect 587422 509818 587658 510054
rect 587422 509498 587658 509734
rect 587422 473818 587658 474054
rect 587422 473498 587658 473734
rect 587422 437818 587658 438054
rect 587422 437498 587658 437734
rect 587422 401818 587658 402054
rect 587422 401498 587658 401734
rect 587422 365818 587658 366054
rect 587422 365498 587658 365734
rect 587422 329818 587658 330054
rect 587422 329498 587658 329734
rect 587422 293818 587658 294054
rect 587422 293498 587658 293734
rect 587422 257818 587658 258054
rect 587422 257498 587658 257734
rect 587422 221818 587658 222054
rect 587422 221498 587658 221734
rect 587422 185818 587658 186054
rect 587422 185498 587658 185734
rect 587422 149818 587658 150054
rect 587422 149498 587658 149734
rect 587422 113818 587658 114054
rect 587422 113498 587658 113734
rect 587422 77818 587658 78054
rect 587422 77498 587658 77734
rect 587422 41818 587658 42054
rect 587422 41498 587658 41734
rect 587422 5818 587658 6054
rect 587422 5498 587658 5734
rect 580586 -2502 580822 -2266
rect 580586 -2822 580822 -2586
rect 587422 -2502 587658 -2266
rect 587422 -2822 587658 -2586
rect 588382 671818 588618 672054
rect 588382 671498 588618 671734
rect 588382 635818 588618 636054
rect 588382 635498 588618 635734
rect 588382 599818 588618 600054
rect 588382 599498 588618 599734
rect 588382 563818 588618 564054
rect 588382 563498 588618 563734
rect 588382 527818 588618 528054
rect 588382 527498 588618 527734
rect 588382 491818 588618 492054
rect 588382 491498 588618 491734
rect 588382 455818 588618 456054
rect 588382 455498 588618 455734
rect 588382 419818 588618 420054
rect 588382 419498 588618 419734
rect 588382 383818 588618 384054
rect 588382 383498 588618 383734
rect 588382 347818 588618 348054
rect 588382 347498 588618 347734
rect 588382 311818 588618 312054
rect 588382 311498 588618 311734
rect 588382 275818 588618 276054
rect 588382 275498 588618 275734
rect 588382 239818 588618 240054
rect 588382 239498 588618 239734
rect 588382 203818 588618 204054
rect 588382 203498 588618 203734
rect 588382 167818 588618 168054
rect 588382 167498 588618 167734
rect 588382 131818 588618 132054
rect 588382 131498 588618 131734
rect 588382 95818 588618 96054
rect 588382 95498 588618 95734
rect 588382 59818 588618 60054
rect 588382 59498 588618 59734
rect 588382 23818 588618 24054
rect 588382 23498 588618 23734
rect 588382 -3462 588618 -3226
rect 588382 -3782 588618 -3546
<< metal5 >>
rect -4876 707740 -4276 707742
rect 22404 707740 23004 707742
rect 58404 707740 59004 707742
rect 94404 707740 95004 707742
rect 130404 707740 131004 707742
rect 166404 707740 167004 707742
rect 202404 707740 203004 707742
rect 238404 707740 239004 707742
rect 274404 707740 275004 707742
rect 310404 707740 311004 707742
rect 346404 707740 347004 707742
rect 382404 707740 383004 707742
rect 418404 707740 419004 707742
rect 454404 707740 455004 707742
rect 490404 707740 491004 707742
rect 526404 707740 527004 707742
rect 562404 707740 563004 707742
rect 588200 707740 588800 707742
rect -4876 707718 588800 707740
rect -4876 707482 -4694 707718
rect -4458 707482 22586 707718
rect 22822 707482 58586 707718
rect 58822 707482 94586 707718
rect 94822 707482 130586 707718
rect 130822 707482 166586 707718
rect 166822 707482 202586 707718
rect 202822 707482 238586 707718
rect 238822 707482 274586 707718
rect 274822 707482 310586 707718
rect 310822 707482 346586 707718
rect 346822 707482 382586 707718
rect 382822 707482 418586 707718
rect 418822 707482 454586 707718
rect 454822 707482 490586 707718
rect 490822 707482 526586 707718
rect 526822 707482 562586 707718
rect 562822 707482 588382 707718
rect 588618 707482 588800 707718
rect -4876 707398 588800 707482
rect -4876 707162 -4694 707398
rect -4458 707162 22586 707398
rect 22822 707162 58586 707398
rect 58822 707162 94586 707398
rect 94822 707162 130586 707398
rect 130822 707162 166586 707398
rect 166822 707162 202586 707398
rect 202822 707162 238586 707398
rect 238822 707162 274586 707398
rect 274822 707162 310586 707398
rect 310822 707162 346586 707398
rect 346822 707162 382586 707398
rect 382822 707162 418586 707398
rect 418822 707162 454586 707398
rect 454822 707162 490586 707398
rect 490822 707162 526586 707398
rect 526822 707162 562586 707398
rect 562822 707162 588382 707398
rect 588618 707162 588800 707398
rect -4876 707140 588800 707162
rect -4876 707138 -4276 707140
rect 22404 707138 23004 707140
rect 58404 707138 59004 707140
rect 94404 707138 95004 707140
rect 130404 707138 131004 707140
rect 166404 707138 167004 707140
rect 202404 707138 203004 707140
rect 238404 707138 239004 707140
rect 274404 707138 275004 707140
rect 310404 707138 311004 707140
rect 346404 707138 347004 707140
rect 382404 707138 383004 707140
rect 418404 707138 419004 707140
rect 454404 707138 455004 707140
rect 490404 707138 491004 707140
rect 526404 707138 527004 707140
rect 562404 707138 563004 707140
rect 588200 707138 588800 707140
rect -3916 706780 -3316 706782
rect 4404 706780 5004 706782
rect 40404 706780 41004 706782
rect 76404 706780 77004 706782
rect 112404 706780 113004 706782
rect 148404 706780 149004 706782
rect 184404 706780 185004 706782
rect 220404 706780 221004 706782
rect 256404 706780 257004 706782
rect 292404 706780 293004 706782
rect 328404 706780 329004 706782
rect 364404 706780 365004 706782
rect 400404 706780 401004 706782
rect 436404 706780 437004 706782
rect 472404 706780 473004 706782
rect 508404 706780 509004 706782
rect 544404 706780 545004 706782
rect 580404 706780 581004 706782
rect 587240 706780 587840 706782
rect -3916 706758 587840 706780
rect -3916 706522 -3734 706758
rect -3498 706522 4586 706758
rect 4822 706522 40586 706758
rect 40822 706522 76586 706758
rect 76822 706522 112586 706758
rect 112822 706522 148586 706758
rect 148822 706522 184586 706758
rect 184822 706522 220586 706758
rect 220822 706522 256586 706758
rect 256822 706522 292586 706758
rect 292822 706522 328586 706758
rect 328822 706522 364586 706758
rect 364822 706522 400586 706758
rect 400822 706522 436586 706758
rect 436822 706522 472586 706758
rect 472822 706522 508586 706758
rect 508822 706522 544586 706758
rect 544822 706522 580586 706758
rect 580822 706522 587422 706758
rect 587658 706522 587840 706758
rect -3916 706438 587840 706522
rect -3916 706202 -3734 706438
rect -3498 706202 4586 706438
rect 4822 706202 40586 706438
rect 40822 706202 76586 706438
rect 76822 706202 112586 706438
rect 112822 706202 148586 706438
rect 148822 706202 184586 706438
rect 184822 706202 220586 706438
rect 220822 706202 256586 706438
rect 256822 706202 292586 706438
rect 292822 706202 328586 706438
rect 328822 706202 364586 706438
rect 364822 706202 400586 706438
rect 400822 706202 436586 706438
rect 436822 706202 472586 706438
rect 472822 706202 508586 706438
rect 508822 706202 544586 706438
rect 544822 706202 580586 706438
rect 580822 706202 587422 706438
rect 587658 706202 587840 706438
rect -3916 706180 587840 706202
rect -3916 706178 -3316 706180
rect 4404 706178 5004 706180
rect 40404 706178 41004 706180
rect 76404 706178 77004 706180
rect 112404 706178 113004 706180
rect 148404 706178 149004 706180
rect 184404 706178 185004 706180
rect 220404 706178 221004 706180
rect 256404 706178 257004 706180
rect 292404 706178 293004 706180
rect 328404 706178 329004 706180
rect 364404 706178 365004 706180
rect 400404 706178 401004 706180
rect 436404 706178 437004 706180
rect 472404 706178 473004 706180
rect 508404 706178 509004 706180
rect 544404 706178 545004 706180
rect 580404 706178 581004 706180
rect 587240 706178 587840 706180
rect -2956 705820 -2356 705822
rect 18804 705820 19404 705822
rect 54804 705820 55404 705822
rect 90804 705820 91404 705822
rect 126804 705820 127404 705822
rect 162804 705820 163404 705822
rect 198804 705820 199404 705822
rect 234804 705820 235404 705822
rect 270804 705820 271404 705822
rect 306804 705820 307404 705822
rect 342804 705820 343404 705822
rect 378804 705820 379404 705822
rect 414804 705820 415404 705822
rect 450804 705820 451404 705822
rect 486804 705820 487404 705822
rect 522804 705820 523404 705822
rect 558804 705820 559404 705822
rect 586280 705820 586880 705822
rect -2956 705798 586880 705820
rect -2956 705562 -2774 705798
rect -2538 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586462 705798
rect 586698 705562 586880 705798
rect -2956 705478 586880 705562
rect -2956 705242 -2774 705478
rect -2538 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586462 705478
rect 586698 705242 586880 705478
rect -2956 705220 586880 705242
rect -2956 705218 -2356 705220
rect 18804 705218 19404 705220
rect 54804 705218 55404 705220
rect 90804 705218 91404 705220
rect 126804 705218 127404 705220
rect 162804 705218 163404 705220
rect 198804 705218 199404 705220
rect 234804 705218 235404 705220
rect 270804 705218 271404 705220
rect 306804 705218 307404 705220
rect 342804 705218 343404 705220
rect 378804 705218 379404 705220
rect 414804 705218 415404 705220
rect 450804 705218 451404 705220
rect 486804 705218 487404 705220
rect 522804 705218 523404 705220
rect 558804 705218 559404 705220
rect 586280 705218 586880 705220
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -3916 690076 -3316 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587240 690076 587840 690078
rect -4876 690054 588800 690076
rect -4876 689818 -3734 690054
rect -3498 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587422 690054
rect 587658 689818 588800 690054
rect -4876 689734 588800 689818
rect -4876 689498 -3734 689734
rect -3498 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587422 689734
rect 587658 689498 588800 689734
rect -4876 689476 588800 689498
rect -3916 689474 -3316 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587240 689474 587840 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2956 686454 586880 686476
rect -2956 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586880 686454
rect -2956 686134 586880 686218
rect -2956 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586880 686134
rect -2956 685876 586880 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -4876 672076 -4276 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588200 672076 588800 672078
rect -4876 672054 588800 672076
rect -4876 671818 -4694 672054
rect -4458 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588382 672054
rect 588618 671818 588800 672054
rect -4876 671734 588800 671818
rect -4876 671498 -4694 671734
rect -4458 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588382 671734
rect 588618 671498 588800 671734
rect -4876 671476 588800 671498
rect -4876 671474 -4276 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588200 671474 588800 671476
rect -2956 668476 -2356 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586280 668476 586880 668478
rect -2956 668454 586880 668476
rect -2956 668218 -2774 668454
rect -2538 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586462 668454
rect 586698 668218 586880 668454
rect -2956 668134 586880 668218
rect -2956 667898 -2774 668134
rect -2538 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586462 668134
rect 586698 667898 586880 668134
rect -2956 667876 586880 667898
rect -2956 667874 -2356 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586280 667874 586880 667876
rect -3916 654076 -3316 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587240 654076 587840 654078
rect -4876 654054 588800 654076
rect -4876 653818 -3734 654054
rect -3498 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587422 654054
rect 587658 653818 588800 654054
rect -4876 653734 588800 653818
rect -4876 653498 -3734 653734
rect -3498 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587422 653734
rect 587658 653498 588800 653734
rect -4876 653476 588800 653498
rect -3916 653474 -3316 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587240 653474 587840 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2956 650454 586880 650476
rect -2956 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586880 650454
rect -2956 650134 586880 650218
rect -2956 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586880 650134
rect -2956 649876 586880 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -4876 636076 -4276 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588200 636076 588800 636078
rect -4876 636054 588800 636076
rect -4876 635818 -4694 636054
rect -4458 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588382 636054
rect 588618 635818 588800 636054
rect -4876 635734 588800 635818
rect -4876 635498 -4694 635734
rect -4458 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588382 635734
rect 588618 635498 588800 635734
rect -4876 635476 588800 635498
rect -4876 635474 -4276 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588200 635474 588800 635476
rect -2956 632476 -2356 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586280 632476 586880 632478
rect -2956 632454 586880 632476
rect -2956 632218 -2774 632454
rect -2538 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586462 632454
rect 586698 632218 586880 632454
rect -2956 632134 586880 632218
rect -2956 631898 -2774 632134
rect -2538 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586462 632134
rect 586698 631898 586880 632134
rect -2956 631876 586880 631898
rect -2956 631874 -2356 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586280 631874 586880 631876
rect -3916 618076 -3316 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587240 618076 587840 618078
rect -4876 618054 588800 618076
rect -4876 617818 -3734 618054
rect -3498 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587422 618054
rect 587658 617818 588800 618054
rect -4876 617734 588800 617818
rect -4876 617498 -3734 617734
rect -3498 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587422 617734
rect 587658 617498 588800 617734
rect -4876 617476 588800 617498
rect -3916 617474 -3316 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587240 617474 587840 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2956 614454 586880 614476
rect -2956 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586880 614454
rect -2956 614134 586880 614218
rect -2956 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586880 614134
rect -2956 613876 586880 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -4876 600076 -4276 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588200 600076 588800 600078
rect -4876 600054 588800 600076
rect -4876 599818 -4694 600054
rect -4458 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588382 600054
rect 588618 599818 588800 600054
rect -4876 599734 588800 599818
rect -4876 599498 -4694 599734
rect -4458 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588382 599734
rect 588618 599498 588800 599734
rect -4876 599476 588800 599498
rect -4876 599474 -4276 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588200 599474 588800 599476
rect -2956 596476 -2356 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586280 596476 586880 596478
rect -2956 596454 586880 596476
rect -2956 596218 -2774 596454
rect -2538 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586462 596454
rect 586698 596218 586880 596454
rect -2956 596134 586880 596218
rect -2956 595898 -2774 596134
rect -2538 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586462 596134
rect 586698 595898 586880 596134
rect -2956 595876 586880 595898
rect -2956 595874 -2356 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586280 595874 586880 595876
rect -3916 582076 -3316 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587240 582076 587840 582078
rect -4876 582054 588800 582076
rect -4876 581818 -3734 582054
rect -3498 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587422 582054
rect 587658 581818 588800 582054
rect -4876 581734 588800 581818
rect -4876 581498 -3734 581734
rect -3498 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587422 581734
rect 587658 581498 588800 581734
rect -4876 581476 588800 581498
rect -3916 581474 -3316 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587240 581474 587840 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2956 578454 586880 578476
rect -2956 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586880 578454
rect -2956 578134 586880 578218
rect -2956 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586880 578134
rect -2956 577876 586880 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -4876 564076 -4276 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588200 564076 588800 564078
rect -4876 564054 588800 564076
rect -4876 563818 -4694 564054
rect -4458 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588382 564054
rect 588618 563818 588800 564054
rect -4876 563734 588800 563818
rect -4876 563498 -4694 563734
rect -4458 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588382 563734
rect 588618 563498 588800 563734
rect -4876 563476 588800 563498
rect -4876 563474 -4276 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588200 563474 588800 563476
rect -2956 560476 -2356 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586280 560476 586880 560478
rect -2956 560454 586880 560476
rect -2956 560218 -2774 560454
rect -2538 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586462 560454
rect 586698 560218 586880 560454
rect -2956 560134 586880 560218
rect -2956 559898 -2774 560134
rect -2538 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586462 560134
rect 586698 559898 586880 560134
rect -2956 559876 586880 559898
rect -2956 559874 -2356 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586280 559874 586880 559876
rect -3916 546076 -3316 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587240 546076 587840 546078
rect -4876 546054 588800 546076
rect -4876 545818 -3734 546054
rect -3498 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587422 546054
rect 587658 545818 588800 546054
rect -4876 545734 588800 545818
rect -4876 545498 -3734 545734
rect -3498 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587422 545734
rect 587658 545498 588800 545734
rect -4876 545476 588800 545498
rect -3916 545474 -3316 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587240 545474 587840 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2956 542454 586880 542476
rect -2956 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586880 542454
rect -2956 542134 586880 542218
rect -2956 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586880 542134
rect -2956 541876 586880 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -4876 528076 -4276 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588200 528076 588800 528078
rect -4876 528054 588800 528076
rect -4876 527818 -4694 528054
rect -4458 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588382 528054
rect 588618 527818 588800 528054
rect -4876 527734 588800 527818
rect -4876 527498 -4694 527734
rect -4458 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588382 527734
rect 588618 527498 588800 527734
rect -4876 527476 588800 527498
rect -4876 527474 -4276 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588200 527474 588800 527476
rect -2956 524476 -2356 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586280 524476 586880 524478
rect -2956 524454 586880 524476
rect -2956 524218 -2774 524454
rect -2538 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586462 524454
rect 586698 524218 586880 524454
rect -2956 524134 586880 524218
rect -2956 523898 -2774 524134
rect -2538 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586462 524134
rect 586698 523898 586880 524134
rect -2956 523876 586880 523898
rect -2956 523874 -2356 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586280 523874 586880 523876
rect -3916 510076 -3316 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587240 510076 587840 510078
rect -4876 510054 588800 510076
rect -4876 509818 -3734 510054
rect -3498 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587422 510054
rect 587658 509818 588800 510054
rect -4876 509734 588800 509818
rect -4876 509498 -3734 509734
rect -3498 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587422 509734
rect 587658 509498 588800 509734
rect -4876 509476 588800 509498
rect -3916 509474 -3316 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587240 509474 587840 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2956 506454 586880 506476
rect -2956 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586880 506454
rect -2956 506134 586880 506218
rect -2956 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586880 506134
rect -2956 505876 586880 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -4876 492076 -4276 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588200 492076 588800 492078
rect -4876 492054 588800 492076
rect -4876 491818 -4694 492054
rect -4458 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588382 492054
rect 588618 491818 588800 492054
rect -4876 491734 588800 491818
rect -4876 491498 -4694 491734
rect -4458 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588382 491734
rect 588618 491498 588800 491734
rect -4876 491476 588800 491498
rect -4876 491474 -4276 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588200 491474 588800 491476
rect -2956 488476 -2356 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586280 488476 586880 488478
rect -2956 488454 586880 488476
rect -2956 488218 -2774 488454
rect -2538 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586462 488454
rect 586698 488218 586880 488454
rect -2956 488134 586880 488218
rect -2956 487898 -2774 488134
rect -2538 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586462 488134
rect 586698 487898 586880 488134
rect -2956 487876 586880 487898
rect -2956 487874 -2356 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586280 487874 586880 487876
rect -3916 474076 -3316 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587240 474076 587840 474078
rect -4876 474054 588800 474076
rect -4876 473818 -3734 474054
rect -3498 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587422 474054
rect 587658 473818 588800 474054
rect -4876 473734 588800 473818
rect -4876 473498 -3734 473734
rect -3498 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587422 473734
rect 587658 473498 588800 473734
rect -4876 473476 588800 473498
rect -3916 473474 -3316 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587240 473474 587840 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2956 470454 586880 470476
rect -2956 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586880 470454
rect -2956 470134 586880 470218
rect -2956 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586880 470134
rect -2956 469876 586880 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -4876 456076 -4276 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588200 456076 588800 456078
rect -4876 456054 588800 456076
rect -4876 455818 -4694 456054
rect -4458 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588382 456054
rect 588618 455818 588800 456054
rect -4876 455734 588800 455818
rect -4876 455498 -4694 455734
rect -4458 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588382 455734
rect 588618 455498 588800 455734
rect -4876 455476 588800 455498
rect -4876 455474 -4276 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588200 455474 588800 455476
rect -2956 452476 -2356 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586280 452476 586880 452478
rect -2956 452454 586880 452476
rect -2956 452218 -2774 452454
rect -2538 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586462 452454
rect 586698 452218 586880 452454
rect -2956 452134 586880 452218
rect -2956 451898 -2774 452134
rect -2538 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586462 452134
rect 586698 451898 586880 452134
rect -2956 451876 586880 451898
rect -2956 451874 -2356 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586280 451874 586880 451876
rect -3916 438076 -3316 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587240 438076 587840 438078
rect -4876 438054 588800 438076
rect -4876 437818 -3734 438054
rect -3498 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587422 438054
rect 587658 437818 588800 438054
rect -4876 437734 588800 437818
rect -4876 437498 -3734 437734
rect -3498 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587422 437734
rect 587658 437498 588800 437734
rect -4876 437476 588800 437498
rect -3916 437474 -3316 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587240 437474 587840 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2956 434454 586880 434476
rect -2956 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586880 434454
rect -2956 434134 586880 434218
rect -2956 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586880 434134
rect -2956 433876 586880 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -4876 420076 -4276 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 101568 420076 101888 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588200 420076 588800 420078
rect -4876 420054 588800 420076
rect -4876 419818 -4694 420054
rect -4458 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 101610 420054
rect 101846 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588382 420054
rect 588618 419818 588800 420054
rect -4876 419734 588800 419818
rect -4876 419498 -4694 419734
rect -4458 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 101610 419734
rect 101846 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588382 419734
rect 588618 419498 588800 419734
rect -4876 419476 588800 419498
rect -4876 419474 -4276 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 101568 419474 101888 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588200 419474 588800 419476
rect -2956 416476 -2356 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 101568 416476 101888 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586280 416476 586880 416478
rect -2956 416454 586880 416476
rect -2956 416218 -2774 416454
rect -2538 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 101610 416454
rect 101846 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586462 416454
rect 586698 416218 586880 416454
rect -2956 416134 586880 416218
rect -2956 415898 -2774 416134
rect -2538 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 101610 416134
rect 101846 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586462 416134
rect 586698 415898 586880 416134
rect -2956 415876 586880 415898
rect -2956 415874 -2356 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 101568 415874 101888 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586280 415874 586880 415876
rect -3916 402076 -3316 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 86208 402076 86528 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587240 402076 587840 402078
rect -4876 402054 588800 402076
rect -4876 401818 -3734 402054
rect -3498 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 86250 402054
rect 86486 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587422 402054
rect 587658 401818 588800 402054
rect -4876 401734 588800 401818
rect -4876 401498 -3734 401734
rect -3498 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 86250 401734
rect 86486 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587422 401734
rect 587658 401498 588800 401734
rect -4876 401476 588800 401498
rect -3916 401474 -3316 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 86208 401474 86528 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587240 401474 587840 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 86208 398476 86528 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2956 398454 586880 398476
rect -2956 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 86250 398454
rect 86486 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586880 398454
rect -2956 398134 586880 398218
rect -2956 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 86250 398134
rect 86486 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586880 398134
rect -2956 397876 586880 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 86208 397874 86528 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -4876 384076 -4276 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 101568 384076 101888 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588200 384076 588800 384078
rect -4876 384054 588800 384076
rect -4876 383818 -4694 384054
rect -4458 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 101610 384054
rect 101846 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588382 384054
rect 588618 383818 588800 384054
rect -4876 383734 588800 383818
rect -4876 383498 -4694 383734
rect -4458 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 101610 383734
rect 101846 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588382 383734
rect 588618 383498 588800 383734
rect -4876 383476 588800 383498
rect -4876 383474 -4276 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 101568 383474 101888 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588200 383474 588800 383476
rect -2956 380476 -2356 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 101568 380476 101888 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586280 380476 586880 380478
rect -2956 380454 586880 380476
rect -2956 380218 -2774 380454
rect -2538 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 101610 380454
rect 101846 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586462 380454
rect 586698 380218 586880 380454
rect -2956 380134 586880 380218
rect -2956 379898 -2774 380134
rect -2538 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 101610 380134
rect 101846 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586462 380134
rect 586698 379898 586880 380134
rect -2956 379876 586880 379898
rect -2956 379874 -2356 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 101568 379874 101888 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586280 379874 586880 379876
rect -3916 366076 -3316 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 86208 366076 86528 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587240 366076 587840 366078
rect -4876 366054 588800 366076
rect -4876 365818 -3734 366054
rect -3498 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 86250 366054
rect 86486 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587422 366054
rect 587658 365818 588800 366054
rect -4876 365734 588800 365818
rect -4876 365498 -3734 365734
rect -3498 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 86250 365734
rect 86486 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587422 365734
rect 587658 365498 588800 365734
rect -4876 365476 588800 365498
rect -3916 365474 -3316 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 86208 365474 86528 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587240 365474 587840 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 86208 362476 86528 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2956 362454 586880 362476
rect -2956 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 86250 362454
rect 86486 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586880 362454
rect -2956 362134 586880 362218
rect -2956 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 86250 362134
rect 86486 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586880 362134
rect -2956 361876 586880 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 86208 361874 86528 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -4876 348076 -4276 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 101568 348076 101888 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588200 348076 588800 348078
rect -4876 348054 588800 348076
rect -4876 347818 -4694 348054
rect -4458 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 101610 348054
rect 101846 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588382 348054
rect 588618 347818 588800 348054
rect -4876 347734 588800 347818
rect -4876 347498 -4694 347734
rect -4458 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 101610 347734
rect 101846 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588382 347734
rect 588618 347498 588800 347734
rect -4876 347476 588800 347498
rect -4876 347474 -4276 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 101568 347474 101888 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588200 347474 588800 347476
rect -2956 344476 -2356 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 101568 344476 101888 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586280 344476 586880 344478
rect -2956 344454 586880 344476
rect -2956 344218 -2774 344454
rect -2538 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 101610 344454
rect 101846 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586462 344454
rect 586698 344218 586880 344454
rect -2956 344134 586880 344218
rect -2956 343898 -2774 344134
rect -2538 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 101610 344134
rect 101846 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586462 344134
rect 586698 343898 586880 344134
rect -2956 343876 586880 343898
rect -2956 343874 -2356 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 101568 343874 101888 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586280 343874 586880 343876
rect -3916 330076 -3316 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 86208 330076 86528 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587240 330076 587840 330078
rect -4876 330054 588800 330076
rect -4876 329818 -3734 330054
rect -3498 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 86250 330054
rect 86486 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587422 330054
rect 587658 329818 588800 330054
rect -4876 329734 588800 329818
rect -4876 329498 -3734 329734
rect -3498 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 86250 329734
rect 86486 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587422 329734
rect 587658 329498 588800 329734
rect -4876 329476 588800 329498
rect -3916 329474 -3316 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 86208 329474 86528 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587240 329474 587840 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 86208 326476 86528 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2956 326454 586880 326476
rect -2956 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 86250 326454
rect 86486 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586880 326454
rect -2956 326134 586880 326218
rect -2956 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 86250 326134
rect 86486 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586880 326134
rect -2956 325876 586880 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 86208 325874 86528 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -4876 312076 -4276 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 101568 312076 101888 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588200 312076 588800 312078
rect -4876 312054 588800 312076
rect -4876 311818 -4694 312054
rect -4458 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 101610 312054
rect 101846 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588382 312054
rect 588618 311818 588800 312054
rect -4876 311734 588800 311818
rect -4876 311498 -4694 311734
rect -4458 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 101610 311734
rect 101846 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588382 311734
rect 588618 311498 588800 311734
rect -4876 311476 588800 311498
rect -4876 311474 -4276 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 101568 311474 101888 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588200 311474 588800 311476
rect -2956 308476 -2356 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 101568 308476 101888 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586280 308476 586880 308478
rect -2956 308454 586880 308476
rect -2956 308218 -2774 308454
rect -2538 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 101610 308454
rect 101846 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586462 308454
rect 586698 308218 586880 308454
rect -2956 308134 586880 308218
rect -2956 307898 -2774 308134
rect -2538 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 101610 308134
rect 101846 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586462 308134
rect 586698 307898 586880 308134
rect -2956 307876 586880 307898
rect -2956 307874 -2356 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 101568 307874 101888 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586280 307874 586880 307876
rect -3916 294076 -3316 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 86208 294076 86528 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587240 294076 587840 294078
rect -4876 294054 588800 294076
rect -4876 293818 -3734 294054
rect -3498 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 86250 294054
rect 86486 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587422 294054
rect 587658 293818 588800 294054
rect -4876 293734 588800 293818
rect -4876 293498 -3734 293734
rect -3498 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 86250 293734
rect 86486 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587422 293734
rect 587658 293498 588800 293734
rect -4876 293476 588800 293498
rect -3916 293474 -3316 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 86208 293474 86528 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587240 293474 587840 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 86208 290476 86528 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2956 290454 586880 290476
rect -2956 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 86250 290454
rect 86486 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586880 290454
rect -2956 290134 586880 290218
rect -2956 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 86250 290134
rect 86486 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586880 290134
rect -2956 289876 586880 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 86208 289874 86528 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -4876 276076 -4276 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 101568 276076 101888 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588200 276076 588800 276078
rect -4876 276054 588800 276076
rect -4876 275818 -4694 276054
rect -4458 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 101610 276054
rect 101846 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588382 276054
rect 588618 275818 588800 276054
rect -4876 275734 588800 275818
rect -4876 275498 -4694 275734
rect -4458 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 101610 275734
rect 101846 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588382 275734
rect 588618 275498 588800 275734
rect -4876 275476 588800 275498
rect -4876 275474 -4276 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 101568 275474 101888 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588200 275474 588800 275476
rect -2956 272476 -2356 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 101568 272476 101888 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586280 272476 586880 272478
rect -2956 272454 586880 272476
rect -2956 272218 -2774 272454
rect -2538 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 101610 272454
rect 101846 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586462 272454
rect 586698 272218 586880 272454
rect -2956 272134 586880 272218
rect -2956 271898 -2774 272134
rect -2538 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 101610 272134
rect 101846 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586462 272134
rect 586698 271898 586880 272134
rect -2956 271876 586880 271898
rect -2956 271874 -2356 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 101568 271874 101888 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586280 271874 586880 271876
rect -3916 258076 -3316 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 86208 258076 86528 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587240 258076 587840 258078
rect -4876 258054 588800 258076
rect -4876 257818 -3734 258054
rect -3498 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 86250 258054
rect 86486 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587422 258054
rect 587658 257818 588800 258054
rect -4876 257734 588800 257818
rect -4876 257498 -3734 257734
rect -3498 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 86250 257734
rect 86486 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587422 257734
rect 587658 257498 588800 257734
rect -4876 257476 588800 257498
rect -3916 257474 -3316 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 86208 257474 86528 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587240 257474 587840 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 86208 254476 86528 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2956 254454 586880 254476
rect -2956 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 86250 254454
rect 86486 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586880 254454
rect -2956 254134 586880 254218
rect -2956 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 86250 254134
rect 86486 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586880 254134
rect -2956 253876 586880 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 86208 253874 86528 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -4876 240076 -4276 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 101568 240076 101888 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588200 240076 588800 240078
rect -4876 240054 588800 240076
rect -4876 239818 -4694 240054
rect -4458 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 101610 240054
rect 101846 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588382 240054
rect 588618 239818 588800 240054
rect -4876 239734 588800 239818
rect -4876 239498 -4694 239734
rect -4458 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 101610 239734
rect 101846 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588382 239734
rect 588618 239498 588800 239734
rect -4876 239476 588800 239498
rect -4876 239474 -4276 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 101568 239474 101888 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588200 239474 588800 239476
rect -2956 236476 -2356 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 101568 236476 101888 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586280 236476 586880 236478
rect -2956 236454 586880 236476
rect -2956 236218 -2774 236454
rect -2538 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 101610 236454
rect 101846 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586462 236454
rect 586698 236218 586880 236454
rect -2956 236134 586880 236218
rect -2956 235898 -2774 236134
rect -2538 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 101610 236134
rect 101846 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586462 236134
rect 586698 235898 586880 236134
rect -2956 235876 586880 235898
rect -2956 235874 -2356 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 101568 235874 101888 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586280 235874 586880 235876
rect -3916 222076 -3316 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 86208 222076 86528 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587240 222076 587840 222078
rect -4876 222054 588800 222076
rect -4876 221818 -3734 222054
rect -3498 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 86250 222054
rect 86486 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587422 222054
rect 587658 221818 588800 222054
rect -4876 221734 588800 221818
rect -4876 221498 -3734 221734
rect -3498 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 86250 221734
rect 86486 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587422 221734
rect 587658 221498 588800 221734
rect -4876 221476 588800 221498
rect -3916 221474 -3316 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 86208 221474 86528 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587240 221474 587840 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 86208 218476 86528 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2956 218454 586880 218476
rect -2956 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 86250 218454
rect 86486 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586880 218454
rect -2956 218134 586880 218218
rect -2956 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 86250 218134
rect 86486 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586880 218134
rect -2956 217876 586880 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 86208 217874 86528 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -4876 204076 -4276 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 101568 204076 101888 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588200 204076 588800 204078
rect -4876 204054 588800 204076
rect -4876 203818 -4694 204054
rect -4458 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 101610 204054
rect 101846 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588382 204054
rect 588618 203818 588800 204054
rect -4876 203734 588800 203818
rect -4876 203498 -4694 203734
rect -4458 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 101610 203734
rect 101846 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588382 203734
rect 588618 203498 588800 203734
rect -4876 203476 588800 203498
rect -4876 203474 -4276 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 101568 203474 101888 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588200 203474 588800 203476
rect -2956 200476 -2356 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 101568 200476 101888 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586280 200476 586880 200478
rect -2956 200454 586880 200476
rect -2956 200218 -2774 200454
rect -2538 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 101610 200454
rect 101846 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586462 200454
rect 586698 200218 586880 200454
rect -2956 200134 586880 200218
rect -2956 199898 -2774 200134
rect -2538 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 101610 200134
rect 101846 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586462 200134
rect 586698 199898 586880 200134
rect -2956 199876 586880 199898
rect -2956 199874 -2356 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 101568 199874 101888 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586280 199874 586880 199876
rect -3916 186076 -3316 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 86208 186076 86528 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587240 186076 587840 186078
rect -4876 186054 588800 186076
rect -4876 185818 -3734 186054
rect -3498 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 86250 186054
rect 86486 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587422 186054
rect 587658 185818 588800 186054
rect -4876 185734 588800 185818
rect -4876 185498 -3734 185734
rect -3498 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 86250 185734
rect 86486 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587422 185734
rect 587658 185498 588800 185734
rect -4876 185476 588800 185498
rect -3916 185474 -3316 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 86208 185474 86528 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587240 185474 587840 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 86208 182476 86528 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2956 182454 586880 182476
rect -2956 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 86250 182454
rect 86486 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586880 182454
rect -2956 182134 586880 182218
rect -2956 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 86250 182134
rect 86486 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586880 182134
rect -2956 181876 586880 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 86208 181874 86528 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -4876 168076 -4276 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 101568 168076 101888 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588200 168076 588800 168078
rect -4876 168054 588800 168076
rect -4876 167818 -4694 168054
rect -4458 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 101610 168054
rect 101846 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588382 168054
rect 588618 167818 588800 168054
rect -4876 167734 588800 167818
rect -4876 167498 -4694 167734
rect -4458 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 101610 167734
rect 101846 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588382 167734
rect 588618 167498 588800 167734
rect -4876 167476 588800 167498
rect -4876 167474 -4276 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 101568 167474 101888 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588200 167474 588800 167476
rect -2956 164476 -2356 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 101568 164476 101888 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586280 164476 586880 164478
rect -2956 164454 586880 164476
rect -2956 164218 -2774 164454
rect -2538 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 101610 164454
rect 101846 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586462 164454
rect 586698 164218 586880 164454
rect -2956 164134 586880 164218
rect -2956 163898 -2774 164134
rect -2538 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 101610 164134
rect 101846 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586462 164134
rect 586698 163898 586880 164134
rect -2956 163876 586880 163898
rect -2956 163874 -2356 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 101568 163874 101888 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586280 163874 586880 163876
rect -3916 150076 -3316 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 86208 150076 86528 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587240 150076 587840 150078
rect -4876 150054 588800 150076
rect -4876 149818 -3734 150054
rect -3498 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 86250 150054
rect 86486 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587422 150054
rect 587658 149818 588800 150054
rect -4876 149734 588800 149818
rect -4876 149498 -3734 149734
rect -3498 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 86250 149734
rect 86486 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587422 149734
rect 587658 149498 588800 149734
rect -4876 149476 588800 149498
rect -3916 149474 -3316 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 86208 149474 86528 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587240 149474 587840 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 86208 146476 86528 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2956 146454 586880 146476
rect -2956 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 86250 146454
rect 86486 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586880 146454
rect -2956 146134 586880 146218
rect -2956 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 86250 146134
rect 86486 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586880 146134
rect -2956 145876 586880 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 86208 145874 86528 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -4876 132076 -4276 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 101568 132076 101888 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588200 132076 588800 132078
rect -4876 132054 588800 132076
rect -4876 131818 -4694 132054
rect -4458 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 101610 132054
rect 101846 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588382 132054
rect 588618 131818 588800 132054
rect -4876 131734 588800 131818
rect -4876 131498 -4694 131734
rect -4458 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 101610 131734
rect 101846 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588382 131734
rect 588618 131498 588800 131734
rect -4876 131476 588800 131498
rect -4876 131474 -4276 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 101568 131474 101888 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588200 131474 588800 131476
rect -2956 128476 -2356 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 101568 128476 101888 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586280 128476 586880 128478
rect -2956 128454 586880 128476
rect -2956 128218 -2774 128454
rect -2538 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 101610 128454
rect 101846 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586462 128454
rect 586698 128218 586880 128454
rect -2956 128134 586880 128218
rect -2956 127898 -2774 128134
rect -2538 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 101610 128134
rect 101846 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586462 128134
rect 586698 127898 586880 128134
rect -2956 127876 586880 127898
rect -2956 127874 -2356 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 101568 127874 101888 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586280 127874 586880 127876
rect -3916 114076 -3316 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 86208 114076 86528 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587240 114076 587840 114078
rect -4876 114054 588800 114076
rect -4876 113818 -3734 114054
rect -3498 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 86250 114054
rect 86486 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587422 114054
rect 587658 113818 588800 114054
rect -4876 113734 588800 113818
rect -4876 113498 -3734 113734
rect -3498 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 86250 113734
rect 86486 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587422 113734
rect 587658 113498 588800 113734
rect -4876 113476 588800 113498
rect -3916 113474 -3316 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 86208 113474 86528 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587240 113474 587840 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 86208 110476 86528 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2956 110454 586880 110476
rect -2956 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 86250 110454
rect 86486 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586880 110454
rect -2956 110134 586880 110218
rect -2956 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 86250 110134
rect 86486 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586880 110134
rect -2956 109876 586880 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 86208 109874 86528 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -4876 96076 -4276 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588200 96076 588800 96078
rect -4876 96054 588800 96076
rect -4876 95818 -4694 96054
rect -4458 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588382 96054
rect 588618 95818 588800 96054
rect -4876 95734 588800 95818
rect -4876 95498 -4694 95734
rect -4458 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588382 95734
rect 588618 95498 588800 95734
rect -4876 95476 588800 95498
rect -4876 95474 -4276 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588200 95474 588800 95476
rect -2956 92476 -2356 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586280 92476 586880 92478
rect -2956 92454 586880 92476
rect -2956 92218 -2774 92454
rect -2538 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586462 92454
rect 586698 92218 586880 92454
rect -2956 92134 586880 92218
rect -2956 91898 -2774 92134
rect -2538 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586462 92134
rect 586698 91898 586880 92134
rect -2956 91876 586880 91898
rect -2956 91874 -2356 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586280 91874 586880 91876
rect -3916 78076 -3316 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587240 78076 587840 78078
rect -4876 78054 588800 78076
rect -4876 77818 -3734 78054
rect -3498 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587422 78054
rect 587658 77818 588800 78054
rect -4876 77734 588800 77818
rect -4876 77498 -3734 77734
rect -3498 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587422 77734
rect 587658 77498 588800 77734
rect -4876 77476 588800 77498
rect -3916 77474 -3316 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587240 77474 587840 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2956 74454 586880 74476
rect -2956 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586880 74454
rect -2956 74134 586880 74218
rect -2956 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586880 74134
rect -2956 73876 586880 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -4876 60076 -4276 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588200 60076 588800 60078
rect -4876 60054 588800 60076
rect -4876 59818 -4694 60054
rect -4458 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588382 60054
rect 588618 59818 588800 60054
rect -4876 59734 588800 59818
rect -4876 59498 -4694 59734
rect -4458 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588382 59734
rect 588618 59498 588800 59734
rect -4876 59476 588800 59498
rect -4876 59474 -4276 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588200 59474 588800 59476
rect -2956 56476 -2356 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586280 56476 586880 56478
rect -2956 56454 586880 56476
rect -2956 56218 -2774 56454
rect -2538 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586462 56454
rect 586698 56218 586880 56454
rect -2956 56134 586880 56218
rect -2956 55898 -2774 56134
rect -2538 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586462 56134
rect 586698 55898 586880 56134
rect -2956 55876 586880 55898
rect -2956 55874 -2356 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586280 55874 586880 55876
rect -3916 42076 -3316 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587240 42076 587840 42078
rect -4876 42054 588800 42076
rect -4876 41818 -3734 42054
rect -3498 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587422 42054
rect 587658 41818 588800 42054
rect -4876 41734 588800 41818
rect -4876 41498 -3734 41734
rect -3498 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587422 41734
rect 587658 41498 588800 41734
rect -4876 41476 588800 41498
rect -3916 41474 -3316 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587240 41474 587840 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2956 38454 586880 38476
rect -2956 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586880 38454
rect -2956 38134 586880 38218
rect -2956 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586880 38134
rect -2956 37876 586880 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -4876 24076 -4276 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588200 24076 588800 24078
rect -4876 24054 588800 24076
rect -4876 23818 -4694 24054
rect -4458 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588382 24054
rect 588618 23818 588800 24054
rect -4876 23734 588800 23818
rect -4876 23498 -4694 23734
rect -4458 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588382 23734
rect 588618 23498 588800 23734
rect -4876 23476 588800 23498
rect -4876 23474 -4276 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588200 23474 588800 23476
rect -2956 20476 -2356 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586280 20476 586880 20478
rect -2956 20454 586880 20476
rect -2956 20218 -2774 20454
rect -2538 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586462 20454
rect 586698 20218 586880 20454
rect -2956 20134 586880 20218
rect -2956 19898 -2774 20134
rect -2538 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586462 20134
rect 586698 19898 586880 20134
rect -2956 19876 586880 19898
rect -2956 19874 -2356 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586280 19874 586880 19876
rect -3916 6076 -3316 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587240 6076 587840 6078
rect -4876 6054 588800 6076
rect -4876 5818 -3734 6054
rect -3498 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587422 6054
rect 587658 5818 588800 6054
rect -4876 5734 588800 5818
rect -4876 5498 -3734 5734
rect -3498 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587422 5734
rect 587658 5498 588800 5734
rect -4876 5476 588800 5498
rect -3916 5474 -3316 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587240 5474 587840 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2956 2454 586880 2476
rect -2956 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586880 2454
rect -2956 2134 586880 2218
rect -2956 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586880 2134
rect -2956 1876 586880 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2956 -1284 -2356 -1282
rect 18804 -1284 19404 -1282
rect 54804 -1284 55404 -1282
rect 90804 -1284 91404 -1282
rect 126804 -1284 127404 -1282
rect 162804 -1284 163404 -1282
rect 198804 -1284 199404 -1282
rect 234804 -1284 235404 -1282
rect 270804 -1284 271404 -1282
rect 306804 -1284 307404 -1282
rect 342804 -1284 343404 -1282
rect 378804 -1284 379404 -1282
rect 414804 -1284 415404 -1282
rect 450804 -1284 451404 -1282
rect 486804 -1284 487404 -1282
rect 522804 -1284 523404 -1282
rect 558804 -1284 559404 -1282
rect 586280 -1284 586880 -1282
rect -2956 -1306 586880 -1284
rect -2956 -1542 -2774 -1306
rect -2538 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586462 -1306
rect 586698 -1542 586880 -1306
rect -2956 -1626 586880 -1542
rect -2956 -1862 -2774 -1626
rect -2538 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586462 -1626
rect 586698 -1862 586880 -1626
rect -2956 -1884 586880 -1862
rect -2956 -1886 -2356 -1884
rect 18804 -1886 19404 -1884
rect 54804 -1886 55404 -1884
rect 90804 -1886 91404 -1884
rect 126804 -1886 127404 -1884
rect 162804 -1886 163404 -1884
rect 198804 -1886 199404 -1884
rect 234804 -1886 235404 -1884
rect 270804 -1886 271404 -1884
rect 306804 -1886 307404 -1884
rect 342804 -1886 343404 -1884
rect 378804 -1886 379404 -1884
rect 414804 -1886 415404 -1884
rect 450804 -1886 451404 -1884
rect 486804 -1886 487404 -1884
rect 522804 -1886 523404 -1884
rect 558804 -1886 559404 -1884
rect 586280 -1886 586880 -1884
rect -3916 -2244 -3316 -2242
rect 4404 -2244 5004 -2242
rect 40404 -2244 41004 -2242
rect 76404 -2244 77004 -2242
rect 112404 -2244 113004 -2242
rect 148404 -2244 149004 -2242
rect 184404 -2244 185004 -2242
rect 220404 -2244 221004 -2242
rect 256404 -2244 257004 -2242
rect 292404 -2244 293004 -2242
rect 328404 -2244 329004 -2242
rect 364404 -2244 365004 -2242
rect 400404 -2244 401004 -2242
rect 436404 -2244 437004 -2242
rect 472404 -2244 473004 -2242
rect 508404 -2244 509004 -2242
rect 544404 -2244 545004 -2242
rect 580404 -2244 581004 -2242
rect 587240 -2244 587840 -2242
rect -3916 -2266 587840 -2244
rect -3916 -2502 -3734 -2266
rect -3498 -2502 4586 -2266
rect 4822 -2502 40586 -2266
rect 40822 -2502 76586 -2266
rect 76822 -2502 112586 -2266
rect 112822 -2502 148586 -2266
rect 148822 -2502 184586 -2266
rect 184822 -2502 220586 -2266
rect 220822 -2502 256586 -2266
rect 256822 -2502 292586 -2266
rect 292822 -2502 328586 -2266
rect 328822 -2502 364586 -2266
rect 364822 -2502 400586 -2266
rect 400822 -2502 436586 -2266
rect 436822 -2502 472586 -2266
rect 472822 -2502 508586 -2266
rect 508822 -2502 544586 -2266
rect 544822 -2502 580586 -2266
rect 580822 -2502 587422 -2266
rect 587658 -2502 587840 -2266
rect -3916 -2586 587840 -2502
rect -3916 -2822 -3734 -2586
rect -3498 -2822 4586 -2586
rect 4822 -2822 40586 -2586
rect 40822 -2822 76586 -2586
rect 76822 -2822 112586 -2586
rect 112822 -2822 148586 -2586
rect 148822 -2822 184586 -2586
rect 184822 -2822 220586 -2586
rect 220822 -2822 256586 -2586
rect 256822 -2822 292586 -2586
rect 292822 -2822 328586 -2586
rect 328822 -2822 364586 -2586
rect 364822 -2822 400586 -2586
rect 400822 -2822 436586 -2586
rect 436822 -2822 472586 -2586
rect 472822 -2822 508586 -2586
rect 508822 -2822 544586 -2586
rect 544822 -2822 580586 -2586
rect 580822 -2822 587422 -2586
rect 587658 -2822 587840 -2586
rect -3916 -2844 587840 -2822
rect -3916 -2846 -3316 -2844
rect 4404 -2846 5004 -2844
rect 40404 -2846 41004 -2844
rect 76404 -2846 77004 -2844
rect 112404 -2846 113004 -2844
rect 148404 -2846 149004 -2844
rect 184404 -2846 185004 -2844
rect 220404 -2846 221004 -2844
rect 256404 -2846 257004 -2844
rect 292404 -2846 293004 -2844
rect 328404 -2846 329004 -2844
rect 364404 -2846 365004 -2844
rect 400404 -2846 401004 -2844
rect 436404 -2846 437004 -2844
rect 472404 -2846 473004 -2844
rect 508404 -2846 509004 -2844
rect 544404 -2846 545004 -2844
rect 580404 -2846 581004 -2844
rect 587240 -2846 587840 -2844
rect -4876 -3204 -4276 -3202
rect 22404 -3204 23004 -3202
rect 58404 -3204 59004 -3202
rect 94404 -3204 95004 -3202
rect 130404 -3204 131004 -3202
rect 166404 -3204 167004 -3202
rect 202404 -3204 203004 -3202
rect 238404 -3204 239004 -3202
rect 274404 -3204 275004 -3202
rect 310404 -3204 311004 -3202
rect 346404 -3204 347004 -3202
rect 382404 -3204 383004 -3202
rect 418404 -3204 419004 -3202
rect 454404 -3204 455004 -3202
rect 490404 -3204 491004 -3202
rect 526404 -3204 527004 -3202
rect 562404 -3204 563004 -3202
rect 588200 -3204 588800 -3202
rect -4876 -3226 588800 -3204
rect -4876 -3462 -4694 -3226
rect -4458 -3462 22586 -3226
rect 22822 -3462 58586 -3226
rect 58822 -3462 94586 -3226
rect 94822 -3462 130586 -3226
rect 130822 -3462 166586 -3226
rect 166822 -3462 202586 -3226
rect 202822 -3462 238586 -3226
rect 238822 -3462 274586 -3226
rect 274822 -3462 310586 -3226
rect 310822 -3462 346586 -3226
rect 346822 -3462 382586 -3226
rect 382822 -3462 418586 -3226
rect 418822 -3462 454586 -3226
rect 454822 -3462 490586 -3226
rect 490822 -3462 526586 -3226
rect 526822 -3462 562586 -3226
rect 562822 -3462 588382 -3226
rect 588618 -3462 588800 -3226
rect -4876 -3546 588800 -3462
rect -4876 -3782 -4694 -3546
rect -4458 -3782 22586 -3546
rect 22822 -3782 58586 -3546
rect 58822 -3782 94586 -3546
rect 94822 -3782 130586 -3546
rect 130822 -3782 166586 -3546
rect 166822 -3782 202586 -3546
rect 202822 -3782 238586 -3546
rect 238822 -3782 274586 -3546
rect 274822 -3782 310586 -3546
rect 310822 -3782 346586 -3546
rect 346822 -3782 382586 -3546
rect 382822 -3782 418586 -3546
rect 418822 -3782 454586 -3546
rect 454822 -3782 490586 -3546
rect 490822 -3782 526586 -3546
rect 526822 -3782 562586 -3546
rect 562822 -3782 588382 -3546
rect 588618 -3782 588800 -3546
rect -4876 -3804 588800 -3782
rect -4876 -3806 -4276 -3804
rect 22404 -3806 23004 -3804
rect 58404 -3806 59004 -3804
rect 94404 -3806 95004 -3804
rect 130404 -3806 131004 -3804
rect 166404 -3806 167004 -3804
rect 202404 -3806 203004 -3804
rect 238404 -3806 239004 -3804
rect 274404 -3806 275004 -3804
rect 310404 -3806 311004 -3804
rect 346404 -3806 347004 -3804
rect 382404 -3806 383004 -3804
rect 418404 -3806 419004 -3804
rect 454404 -3806 455004 -3804
rect 490404 -3806 491004 -3804
rect 526404 -3806 527004 -3804
rect 562404 -3806 563004 -3804
rect 588200 -3806 588800 -3804
use Ibtida_top_dffram_cv  mprj
timestamp 1607975982
transform 1 0 82000 0 1 102000
box 0 0 318293 320437
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2956 -1884 586880 -1284 8 vssd1
port 637 nsew default input
rlabel metal5 s -3916 -2844 587840 -2244 8 vccd2
port 638 nsew default input
rlabel metal5 s -4876 -3804 588800 -3204 8 vssd2
port 639 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
