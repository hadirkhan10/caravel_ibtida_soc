VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 972.980 2270.030 973.040 ;
        RECT 2418.290 972.980 2418.610 973.040 ;
        RECT 2269.710 972.840 2418.610 972.980 ;
        RECT 2269.710 972.780 2270.030 972.840 ;
        RECT 2418.290 972.780 2418.610 972.840 ;
        RECT 2418.290 89.660 2418.610 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2418.290 89.520 2899.310 89.660 ;
        RECT 2418.290 89.460 2418.610 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2269.740 972.780 2270.000 973.040 ;
        RECT 2418.320 972.780 2418.580 973.040 ;
        RECT 2418.320 89.460 2418.580 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2269.730 977.995 2270.010 978.365 ;
        RECT 2269.800 973.070 2269.940 977.995 ;
        RECT 2269.740 972.750 2270.000 973.070 ;
        RECT 2418.320 972.750 2418.580 973.070 ;
        RECT 2418.380 89.750 2418.520 972.750 ;
        RECT 2418.320 89.430 2418.580 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2269.730 978.040 2270.010 978.320 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2269.705 978.330 2270.035 978.345 ;
        RECT 2250.780 978.320 2270.035 978.330 ;
        RECT 2247.465 978.030 2270.035 978.320 ;
        RECT 2247.465 977.720 2251.465 978.030 ;
        RECT 2269.705 978.015 2270.035 978.030 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2280.290 2429.200 2280.610 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2280.290 2429.060 2901.150 2429.200 ;
        RECT 2280.290 2429.000 2280.610 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2266.950 2047.040 2267.270 2047.100 ;
        RECT 2280.290 2047.040 2280.610 2047.100 ;
        RECT 2266.950 2046.900 2280.610 2047.040 ;
        RECT 2266.950 2046.840 2267.270 2046.900 ;
        RECT 2280.290 2046.840 2280.610 2046.900 ;
      LAYER via ;
        RECT 2280.320 2429.000 2280.580 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2266.980 2046.840 2267.240 2047.100 ;
        RECT 2280.320 2046.840 2280.580 2047.100 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2280.320 2428.970 2280.580 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2280.380 2047.130 2280.520 2428.970 ;
        RECT 2266.980 2046.810 2267.240 2047.130 ;
        RECT 2280.320 2046.810 2280.580 2047.130 ;
        RECT 2267.040 2045.965 2267.180 2046.810 ;
        RECT 2266.970 2045.595 2267.250 2045.965 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2266.970 2045.640 2267.250 2045.920 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2266.945 2045.930 2267.275 2045.945 ;
        RECT 2250.780 2045.920 2267.275 2045.930 ;
        RECT 2247.465 2045.630 2267.275 2045.920 ;
        RECT 2247.465 2045.320 2251.465 2045.630 ;
        RECT 2266.945 2045.615 2267.275 2045.630 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2425.190 2663.800 2425.510 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2425.190 2663.660 2901.150 2663.800 ;
        RECT 2425.190 2663.600 2425.510 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2269.710 2152.780 2270.030 2152.840 ;
        RECT 2425.190 2152.780 2425.510 2152.840 ;
        RECT 2269.710 2152.640 2425.510 2152.780 ;
        RECT 2269.710 2152.580 2270.030 2152.640 ;
        RECT 2425.190 2152.580 2425.510 2152.640 ;
      LAYER via ;
        RECT 2425.220 2663.600 2425.480 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2269.740 2152.580 2270.000 2152.840 ;
        RECT 2425.220 2152.580 2425.480 2152.840 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2425.220 2663.570 2425.480 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2425.280 2152.870 2425.420 2663.570 ;
        RECT 2269.740 2152.725 2270.000 2152.870 ;
        RECT 2269.730 2152.355 2270.010 2152.725 ;
        RECT 2425.220 2152.550 2425.480 2152.870 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2269.730 2152.400 2270.010 2152.680 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2269.705 2152.690 2270.035 2152.705 ;
        RECT 2250.780 2152.680 2270.035 2152.690 ;
        RECT 2247.465 2152.390 2270.035 2152.680 ;
        RECT 2247.465 2152.080 2251.465 2152.390 ;
        RECT 2269.705 2152.375 2270.035 2152.390 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2445.890 2898.400 2446.210 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2445.890 2898.260 2901.150 2898.400 ;
        RECT 2445.890 2898.200 2446.210 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2269.710 2262.940 2270.030 2263.000 ;
        RECT 2445.890 2262.940 2446.210 2263.000 ;
        RECT 2269.710 2262.800 2446.210 2262.940 ;
        RECT 2269.710 2262.740 2270.030 2262.800 ;
        RECT 2445.890 2262.740 2446.210 2262.800 ;
      LAYER via ;
        RECT 2445.920 2898.200 2446.180 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2269.740 2262.740 2270.000 2263.000 ;
        RECT 2445.920 2262.740 2446.180 2263.000 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2445.920 2898.170 2446.180 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2445.980 2263.030 2446.120 2898.170 ;
        RECT 2269.740 2262.710 2270.000 2263.030 ;
        RECT 2445.920 2262.710 2446.180 2263.030 ;
        RECT 2269.800 2259.485 2269.940 2262.710 ;
        RECT 2269.730 2259.115 2270.010 2259.485 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2269.730 2259.160 2270.010 2259.440 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2269.705 2259.450 2270.035 2259.465 ;
        RECT 2250.780 2259.440 2270.035 2259.450 ;
        RECT 2247.465 2259.150 2270.035 2259.440 ;
        RECT 2247.465 2258.840 2251.465 2259.150 ;
        RECT 2269.705 2259.135 2270.035 2259.150 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2397.590 3133.000 2397.910 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2397.590 3132.860 2901.150 3133.000 ;
        RECT 2397.590 3132.800 2397.910 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2269.710 2366.640 2270.030 2366.700 ;
        RECT 2397.590 2366.640 2397.910 2366.700 ;
        RECT 2269.710 2366.500 2397.910 2366.640 ;
        RECT 2269.710 2366.440 2270.030 2366.500 ;
        RECT 2397.590 2366.440 2397.910 2366.500 ;
      LAYER via ;
        RECT 2397.620 3132.800 2397.880 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2269.740 2366.440 2270.000 2366.700 ;
        RECT 2397.620 2366.440 2397.880 2366.700 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2397.620 3132.770 2397.880 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2397.680 2366.730 2397.820 3132.770 ;
        RECT 2269.740 2366.410 2270.000 2366.730 ;
        RECT 2397.620 2366.410 2397.880 2366.730 ;
        RECT 2269.800 2366.245 2269.940 2366.410 ;
        RECT 2269.730 2365.875 2270.010 2366.245 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2269.730 2365.920 2270.010 2366.200 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2269.705 2366.210 2270.035 2366.225 ;
        RECT 2250.780 2366.200 2270.035 2366.210 ;
        RECT 2247.465 2365.910 2270.035 2366.200 ;
        RECT 2247.465 2365.600 2251.465 2365.910 ;
        RECT 2269.705 2365.895 2270.035 2365.910 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2418.290 3367.600 2418.610 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2418.290 3367.460 2901.150 3367.600 ;
        RECT 2418.290 3367.400 2418.610 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2269.710 2477.140 2270.030 2477.200 ;
        RECT 2418.290 2477.140 2418.610 2477.200 ;
        RECT 2269.710 2477.000 2418.610 2477.140 ;
        RECT 2269.710 2476.940 2270.030 2477.000 ;
        RECT 2418.290 2476.940 2418.610 2477.000 ;
      LAYER via ;
        RECT 2418.320 3367.400 2418.580 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2269.740 2476.940 2270.000 2477.200 ;
        RECT 2418.320 2476.940 2418.580 2477.200 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2418.320 3367.370 2418.580 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2418.380 2477.230 2418.520 3367.370 ;
        RECT 2269.740 2476.910 2270.000 2477.230 ;
        RECT 2418.320 2476.910 2418.580 2477.230 ;
        RECT 2269.800 2473.005 2269.940 2476.910 ;
        RECT 2269.730 2472.635 2270.010 2473.005 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2269.730 2472.680 2270.010 2472.960 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2269.705 2472.970 2270.035 2472.985 ;
        RECT 2250.780 2472.960 2270.035 2472.970 ;
        RECT 2247.465 2472.670 2270.035 2472.960 ;
        RECT 2247.465 2472.360 2251.465 2472.670 ;
        RECT 2269.705 2472.655 2270.035 2472.670 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3415.555 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
        RECT 2795.105 2753.065 2795.275 2801.175 ;
      LAYER mcon ;
        RECT 2796.485 3415.385 2796.655 3415.555 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
        RECT 2795.105 2801.005 2795.275 2801.175 ;
      LAYER met1 ;
        RECT 2794.570 3422.340 2794.890 3422.400 ;
        RECT 2798.250 3422.340 2798.570 3422.400 ;
        RECT 2794.570 3422.200 2798.570 3422.340 ;
        RECT 2794.570 3422.140 2794.890 3422.200 ;
        RECT 2798.250 3422.140 2798.570 3422.200 ;
        RECT 2794.570 3415.540 2794.890 3415.600 ;
        RECT 2796.425 3415.540 2796.715 3415.585 ;
        RECT 2794.570 3415.400 2796.715 3415.540 ;
        RECT 2794.570 3415.340 2794.890 3415.400 ;
        RECT 2796.425 3415.355 2796.715 3415.400 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2795.030 2801.160 2795.350 2801.220 ;
        RECT 2794.835 2801.020 2795.350 2801.160 ;
        RECT 2795.030 2800.960 2795.350 2801.020 ;
        RECT 2795.045 2753.220 2795.335 2753.265 ;
        RECT 2795.950 2753.220 2796.270 2753.280 ;
        RECT 2795.045 2753.080 2796.270 2753.220 ;
        RECT 2795.045 2753.035 2795.335 2753.080 ;
        RECT 2795.950 2753.020 2796.270 2753.080 ;
        RECT 2795.030 2718.200 2795.350 2718.260 ;
        RECT 2795.950 2718.200 2796.270 2718.260 ;
        RECT 2795.030 2718.060 2796.270 2718.200 ;
        RECT 2795.030 2718.000 2795.350 2718.060 ;
        RECT 2795.950 2718.000 2796.270 2718.060 ;
        RECT 2221.870 2577.100 2222.190 2577.160 ;
        RECT 2795.950 2577.100 2796.270 2577.160 ;
        RECT 2221.870 2576.960 2796.270 2577.100 ;
        RECT 2221.870 2576.900 2222.190 2576.960 ;
        RECT 2795.950 2576.900 2796.270 2576.960 ;
      LAYER via ;
        RECT 2794.600 3422.140 2794.860 3422.400 ;
        RECT 2798.280 3422.140 2798.540 3422.400 ;
        RECT 2794.600 3415.340 2794.860 3415.600 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2795.060 2800.960 2795.320 2801.220 ;
        RECT 2795.980 2753.020 2796.240 2753.280 ;
        RECT 2795.060 2718.000 2795.320 2718.260 ;
        RECT 2795.980 2718.000 2796.240 2718.260 ;
        RECT 2221.900 2576.900 2222.160 2577.160 ;
        RECT 2795.980 2576.900 2796.240 2577.160 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.430 2798.480 3517.600 ;
        RECT 2794.600 3422.110 2794.860 3422.430 ;
        RECT 2798.280 3422.110 2798.540 3422.430 ;
        RECT 2794.660 3415.630 2794.800 3422.110 ;
        RECT 2794.600 3415.310 2794.860 3415.630 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.250 2795.260 2814.870 ;
        RECT 2795.060 2800.930 2795.320 2801.250 ;
        RECT 2795.980 2752.990 2796.240 2753.310 ;
        RECT 2796.040 2718.290 2796.180 2752.990 ;
        RECT 2795.060 2717.970 2795.320 2718.290 ;
        RECT 2795.980 2717.970 2796.240 2718.290 ;
        RECT 2795.120 2670.090 2795.260 2717.970 ;
        RECT 2795.120 2669.950 2795.720 2670.090 ;
        RECT 2795.580 2622.490 2795.720 2669.950 ;
        RECT 2795.580 2622.350 2796.180 2622.490 ;
        RECT 2796.040 2577.190 2796.180 2622.350 ;
        RECT 2221.900 2576.870 2222.160 2577.190 ;
        RECT 2795.980 2576.870 2796.240 2577.190 ;
        RECT 2221.960 2562.185 2222.100 2576.870 ;
        RECT 2221.790 2561.900 2222.100 2562.185 ;
        RECT 2221.790 2558.185 2222.070 2561.900 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2470.805 2815.285 2470.975 2849.455 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2470.805 2849.285 2470.975 2849.455 ;
      LAYER met1 ;
        RECT 2471.190 3429.480 2471.510 3429.540 ;
        RECT 2474.410 3429.480 2474.730 3429.540 ;
        RECT 2471.190 3429.340 2474.730 3429.480 ;
        RECT 2471.190 3429.280 2471.510 3429.340 ;
        RECT 2474.410 3429.280 2474.730 3429.340 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2470.535 2849.300 2471.050 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2470.745 2815.440 2471.035 2815.485 ;
        RECT 2471.650 2815.440 2471.970 2815.500 ;
        RECT 2470.745 2815.300 2471.970 2815.440 ;
        RECT 2470.745 2815.255 2471.035 2815.300 ;
        RECT 2471.650 2815.240 2471.970 2815.300 ;
        RECT 2470.730 2753.220 2471.050 2753.280 ;
        RECT 2472.110 2753.220 2472.430 2753.280 ;
        RECT 2470.730 2753.080 2472.430 2753.220 ;
        RECT 2470.730 2753.020 2471.050 2753.080 ;
        RECT 2472.110 2753.020 2472.430 2753.080 ;
        RECT 2472.110 2719.220 2472.430 2719.280 ;
        RECT 2471.740 2719.080 2472.430 2719.220 ;
        RECT 2471.740 2718.600 2471.880 2719.080 ;
        RECT 2472.110 2719.020 2472.430 2719.080 ;
        RECT 2471.650 2718.340 2471.970 2718.600 ;
        RECT 2470.730 2656.660 2471.050 2656.720 ;
        RECT 2472.110 2656.660 2472.430 2656.720 ;
        RECT 2470.730 2656.520 2472.430 2656.660 ;
        RECT 2470.730 2656.460 2471.050 2656.520 ;
        RECT 2472.110 2656.460 2472.430 2656.520 ;
        RECT 2471.190 2608.380 2471.510 2608.440 ;
        RECT 2472.110 2608.380 2472.430 2608.440 ;
        RECT 2471.190 2608.240 2472.430 2608.380 ;
        RECT 2471.190 2608.180 2471.510 2608.240 ;
        RECT 2472.110 2608.180 2472.430 2608.240 ;
        RECT 2045.230 2578.120 2045.550 2578.180 ;
        RECT 2471.190 2578.120 2471.510 2578.180 ;
        RECT 2045.230 2577.980 2471.510 2578.120 ;
        RECT 2045.230 2577.920 2045.550 2577.980 ;
        RECT 2471.190 2577.920 2471.510 2577.980 ;
      LAYER via ;
        RECT 2471.220 3429.280 2471.480 3429.540 ;
        RECT 2474.440 3429.280 2474.700 3429.540 ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 2470.760 2753.020 2471.020 2753.280 ;
        RECT 2472.140 2753.020 2472.400 2753.280 ;
        RECT 2472.140 2719.020 2472.400 2719.280 ;
        RECT 2471.680 2718.340 2471.940 2718.600 ;
        RECT 2470.760 2656.460 2471.020 2656.720 ;
        RECT 2472.140 2656.460 2472.400 2656.720 ;
        RECT 2471.220 2608.180 2471.480 2608.440 ;
        RECT 2472.140 2608.180 2472.400 2608.440 ;
        RECT 2045.260 2577.920 2045.520 2578.180 ;
        RECT 2471.220 2577.920 2471.480 2578.180 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3429.570 2474.640 3517.230 ;
        RECT 2471.220 3429.250 2471.480 3429.570 ;
        RECT 2474.440 3429.250 2474.700 3429.570 ;
        RECT 2471.280 3394.970 2471.420 3429.250 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.685 2469.580 2946.110 ;
        RECT 2469.370 2898.315 2469.650 2898.685 ;
        RECT 2470.290 2898.315 2470.570 2898.685 ;
        RECT 2470.360 2863.210 2470.500 2898.315 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.445 2471.880 2815.210 ;
        RECT 2470.750 2801.075 2471.030 2801.445 ;
        RECT 2471.670 2801.075 2471.950 2801.445 ;
        RECT 2470.820 2753.310 2470.960 2801.075 ;
        RECT 2470.760 2752.990 2471.020 2753.310 ;
        RECT 2472.140 2752.990 2472.400 2753.310 ;
        RECT 2472.200 2719.310 2472.340 2752.990 ;
        RECT 2472.140 2718.990 2472.400 2719.310 ;
        RECT 2471.680 2718.310 2471.940 2718.630 ;
        RECT 2471.740 2704.885 2471.880 2718.310 ;
        RECT 2470.750 2704.515 2471.030 2704.885 ;
        RECT 2471.670 2704.515 2471.950 2704.885 ;
        RECT 2470.820 2656.750 2470.960 2704.515 ;
        RECT 2470.760 2656.430 2471.020 2656.750 ;
        RECT 2472.140 2656.430 2472.400 2656.750 ;
        RECT 2472.200 2608.470 2472.340 2656.430 ;
        RECT 2471.220 2608.150 2471.480 2608.470 ;
        RECT 2472.140 2608.150 2472.400 2608.470 ;
        RECT 2471.280 2578.210 2471.420 2608.150 ;
        RECT 2045.260 2577.890 2045.520 2578.210 ;
        RECT 2471.220 2577.890 2471.480 2578.210 ;
        RECT 2045.320 2562.185 2045.460 2577.890 ;
        RECT 2045.150 2561.900 2045.460 2562.185 ;
        RECT 2045.150 2558.185 2045.430 2561.900 ;
      LAYER via2 ;
        RECT 2469.370 2898.360 2469.650 2898.640 ;
        RECT 2470.290 2898.360 2470.570 2898.640 ;
        RECT 2470.750 2801.120 2471.030 2801.400 ;
        RECT 2471.670 2801.120 2471.950 2801.400 ;
        RECT 2470.750 2704.560 2471.030 2704.840 ;
        RECT 2471.670 2704.560 2471.950 2704.840 ;
      LAYER met3 ;
        RECT 2469.345 2898.650 2469.675 2898.665 ;
        RECT 2470.265 2898.650 2470.595 2898.665 ;
        RECT 2469.345 2898.350 2470.595 2898.650 ;
        RECT 2469.345 2898.335 2469.675 2898.350 ;
        RECT 2470.265 2898.335 2470.595 2898.350 ;
        RECT 2470.725 2801.410 2471.055 2801.425 ;
        RECT 2471.645 2801.410 2471.975 2801.425 ;
        RECT 2470.725 2801.110 2471.975 2801.410 ;
        RECT 2470.725 2801.095 2471.055 2801.110 ;
        RECT 2471.645 2801.095 2471.975 2801.110 ;
        RECT 2470.725 2704.850 2471.055 2704.865 ;
        RECT 2471.645 2704.850 2471.975 2704.865 ;
        RECT 2470.725 2704.550 2471.975 2704.850 ;
        RECT 2470.725 2704.535 2471.055 2704.550 ;
        RECT 2471.645 2704.535 2471.975 2704.550 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3415.555 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
        RECT 2146.505 2753.065 2146.675 2801.175 ;
      LAYER mcon ;
        RECT 2147.885 3415.385 2148.055 3415.555 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
        RECT 2146.505 2801.005 2146.675 2801.175 ;
      LAYER met1 ;
        RECT 2145.970 3422.340 2146.290 3422.400 ;
        RECT 2149.190 3422.340 2149.510 3422.400 ;
        RECT 2145.970 3422.200 2149.510 3422.340 ;
        RECT 2145.970 3422.140 2146.290 3422.200 ;
        RECT 2149.190 3422.140 2149.510 3422.200 ;
        RECT 2145.970 3415.540 2146.290 3415.600 ;
        RECT 2147.825 3415.540 2148.115 3415.585 ;
        RECT 2145.970 3415.400 2148.115 3415.540 ;
        RECT 2145.970 3415.340 2146.290 3415.400 ;
        RECT 2147.825 3415.355 2148.115 3415.400 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2146.235 2801.020 2146.750 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2146.445 2753.220 2146.735 2753.265 ;
        RECT 2147.350 2753.220 2147.670 2753.280 ;
        RECT 2146.445 2753.080 2147.670 2753.220 ;
        RECT 2146.445 2753.035 2146.735 2753.080 ;
        RECT 2147.350 2753.020 2147.670 2753.080 ;
        RECT 2146.430 2718.200 2146.750 2718.260 ;
        RECT 2147.350 2718.200 2147.670 2718.260 ;
        RECT 2146.430 2718.060 2147.670 2718.200 ;
        RECT 2146.430 2718.000 2146.750 2718.060 ;
        RECT 2147.350 2718.000 2147.670 2718.060 ;
        RECT 1868.130 2577.100 1868.450 2577.160 ;
        RECT 2147.350 2577.100 2147.670 2577.160 ;
        RECT 1868.130 2576.960 2147.670 2577.100 ;
        RECT 1868.130 2576.900 1868.450 2576.960 ;
        RECT 2147.350 2576.900 2147.670 2576.960 ;
      LAYER via ;
        RECT 2146.000 3422.140 2146.260 3422.400 ;
        RECT 2149.220 3422.140 2149.480 3422.400 ;
        RECT 2146.000 3415.340 2146.260 3415.600 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2753.020 2147.640 2753.280 ;
        RECT 2146.460 2718.000 2146.720 2718.260 ;
        RECT 2147.380 2718.000 2147.640 2718.260 ;
        RECT 1868.160 2576.900 1868.420 2577.160 ;
        RECT 2147.380 2576.900 2147.640 2577.160 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3422.430 2149.420 3517.600 ;
        RECT 2146.000 3422.110 2146.260 3422.430 ;
        RECT 2149.220 3422.110 2149.480 3422.430 ;
        RECT 2146.060 3415.630 2146.200 3422.110 ;
        RECT 2146.000 3415.310 2146.260 3415.630 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.250 2146.660 2814.870 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2752.990 2147.640 2753.310 ;
        RECT 2147.440 2718.290 2147.580 2752.990 ;
        RECT 2146.460 2717.970 2146.720 2718.290 ;
        RECT 2147.380 2717.970 2147.640 2718.290 ;
        RECT 2146.520 2670.090 2146.660 2717.970 ;
        RECT 2146.520 2669.950 2147.120 2670.090 ;
        RECT 2146.980 2622.490 2147.120 2669.950 ;
        RECT 2146.980 2622.350 2147.580 2622.490 ;
        RECT 2147.440 2577.190 2147.580 2622.350 ;
        RECT 1868.160 2576.870 1868.420 2577.190 ;
        RECT 2147.380 2576.870 2147.640 2577.190 ;
        RECT 1868.220 2562.185 1868.360 2576.870 ;
        RECT 1868.050 2561.900 1868.360 2562.185 ;
        RECT 1868.050 2558.185 1868.330 2561.900 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 2898.245 1821.915 2946.355 ;
        RECT 1822.205 2815.285 1822.375 2849.455 ;
      LAYER mcon ;
        RECT 1821.745 2946.185 1821.915 2946.355 ;
        RECT 1822.205 2849.285 1822.375 2849.455 ;
      LAYER met1 ;
        RECT 1821.670 3464.160 1821.990 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1821.670 3464.020 1825.670 3464.160 ;
        RECT 1821.670 3463.960 1821.990 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1821.670 3367.600 1821.990 3367.660 ;
        RECT 1822.590 3367.600 1822.910 3367.660 ;
        RECT 1821.670 3367.460 1822.910 3367.600 ;
        RECT 1821.670 3367.400 1821.990 3367.460 ;
        RECT 1822.590 3367.400 1822.910 3367.460 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1821.685 2946.340 1821.975 2946.385 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1821.685 2946.200 1822.450 2946.340 ;
        RECT 1821.685 2946.155 1821.975 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1821.670 2898.400 1821.990 2898.460 ;
        RECT 1821.475 2898.260 1821.990 2898.400 ;
        RECT 1821.670 2898.200 1821.990 2898.260 ;
        RECT 1822.130 2849.440 1822.450 2849.500 ;
        RECT 1821.935 2849.300 1822.450 2849.440 ;
        RECT 1822.130 2849.240 1822.450 2849.300 ;
        RECT 1822.145 2815.440 1822.435 2815.485 ;
        RECT 1823.050 2815.440 1823.370 2815.500 ;
        RECT 1822.145 2815.300 1823.370 2815.440 ;
        RECT 1822.145 2815.255 1822.435 2815.300 ;
        RECT 1823.050 2815.240 1823.370 2815.300 ;
        RECT 1822.130 2753.220 1822.450 2753.280 ;
        RECT 1823.510 2753.220 1823.830 2753.280 ;
        RECT 1822.130 2753.080 1823.830 2753.220 ;
        RECT 1822.130 2753.020 1822.450 2753.080 ;
        RECT 1823.510 2753.020 1823.830 2753.080 ;
        RECT 1823.510 2719.220 1823.830 2719.280 ;
        RECT 1823.140 2719.080 1823.830 2719.220 ;
        RECT 1823.140 2718.600 1823.280 2719.080 ;
        RECT 1823.510 2719.020 1823.830 2719.080 ;
        RECT 1823.050 2718.340 1823.370 2718.600 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1822.590 2608.380 1822.910 2608.440 ;
        RECT 1823.510 2608.380 1823.830 2608.440 ;
        RECT 1822.590 2608.240 1823.830 2608.380 ;
        RECT 1822.590 2608.180 1822.910 2608.240 ;
        RECT 1823.510 2608.180 1823.830 2608.240 ;
        RECT 1691.490 2577.100 1691.810 2577.160 ;
        RECT 1822.590 2577.100 1822.910 2577.160 ;
        RECT 1691.490 2576.960 1822.910 2577.100 ;
        RECT 1691.490 2576.900 1691.810 2576.960 ;
        RECT 1822.590 2576.900 1822.910 2576.960 ;
      LAYER via ;
        RECT 1821.700 3463.960 1821.960 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1821.700 3367.400 1821.960 3367.660 ;
        RECT 1822.620 3367.400 1822.880 3367.660 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1821.700 2898.200 1821.960 2898.460 ;
        RECT 1822.160 2849.240 1822.420 2849.500 ;
        RECT 1823.080 2815.240 1823.340 2815.500 ;
        RECT 1822.160 2753.020 1822.420 2753.280 ;
        RECT 1823.540 2753.020 1823.800 2753.280 ;
        RECT 1823.540 2719.020 1823.800 2719.280 ;
        RECT 1823.080 2718.340 1823.340 2718.600 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1822.620 2608.180 1822.880 2608.440 ;
        RECT 1823.540 2608.180 1823.800 2608.440 ;
        RECT 1691.520 2576.900 1691.780 2577.160 ;
        RECT 1822.620 2576.900 1822.880 2577.160 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1821.700 3463.930 1821.960 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1821.760 3415.370 1821.900 3463.930 ;
        RECT 1821.760 3415.230 1822.820 3415.370 ;
        RECT 1822.680 3367.690 1822.820 3415.230 ;
        RECT 1821.700 3367.370 1821.960 3367.690 ;
        RECT 1822.620 3367.370 1822.880 3367.690 ;
        RECT 1821.760 3318.810 1821.900 3367.370 ;
        RECT 1821.760 3318.670 1822.820 3318.810 ;
        RECT 1822.680 3270.790 1822.820 3318.670 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1821.700 2898.170 1821.960 2898.490 ;
        RECT 1821.760 2863.210 1821.900 2898.170 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2849.530 1822.360 2863.070 ;
        RECT 1822.160 2849.210 1822.420 2849.530 ;
        RECT 1823.080 2815.210 1823.340 2815.530 ;
        RECT 1823.140 2801.445 1823.280 2815.210 ;
        RECT 1822.150 2801.075 1822.430 2801.445 ;
        RECT 1823.070 2801.075 1823.350 2801.445 ;
        RECT 1822.220 2753.310 1822.360 2801.075 ;
        RECT 1822.160 2752.990 1822.420 2753.310 ;
        RECT 1823.540 2752.990 1823.800 2753.310 ;
        RECT 1823.600 2719.310 1823.740 2752.990 ;
        RECT 1823.540 2718.990 1823.800 2719.310 ;
        RECT 1823.080 2718.310 1823.340 2718.630 ;
        RECT 1823.140 2704.885 1823.280 2718.310 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2608.470 1823.740 2656.430 ;
        RECT 1822.620 2608.150 1822.880 2608.470 ;
        RECT 1823.540 2608.150 1823.800 2608.470 ;
        RECT 1822.680 2577.190 1822.820 2608.150 ;
        RECT 1691.520 2576.870 1691.780 2577.190 ;
        RECT 1822.620 2576.870 1822.880 2577.190 ;
        RECT 1691.580 2562.185 1691.720 2576.870 ;
        RECT 1691.410 2561.900 1691.720 2562.185 ;
        RECT 1691.410 2558.185 1691.690 2561.900 ;
      LAYER via2 ;
        RECT 1822.150 2801.120 1822.430 2801.400 ;
        RECT 1823.070 2801.120 1823.350 2801.400 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
      LAYER met3 ;
        RECT 1822.125 2801.410 1822.455 2801.425 ;
        RECT 1823.045 2801.410 1823.375 2801.425 ;
        RECT 1822.125 2801.110 1823.375 2801.410 ;
        RECT 1822.125 2801.095 1822.455 2801.110 ;
        RECT 1823.045 2801.095 1823.375 2801.110 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 2574.380 1504.130 2574.440 ;
        RECT 1514.850 2574.380 1515.170 2574.440 ;
        RECT 1503.810 2574.240 1515.170 2574.380 ;
        RECT 1503.810 2574.180 1504.130 2574.240 ;
        RECT 1514.850 2574.180 1515.170 2574.240 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 2574.180 1504.100 2574.440 ;
        RECT 1514.880 2574.180 1515.140 2574.440 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 2574.470 1504.040 3498.270 ;
        RECT 1503.840 2574.150 1504.100 2574.470 ;
        RECT 1514.880 2574.150 1515.140 2574.470 ;
        RECT 1514.940 2562.185 1515.080 2574.150 ;
        RECT 1514.770 2561.900 1515.080 2562.185 ;
        RECT 1514.770 2558.185 1515.050 2561.900 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2268.790 1084.160 2269.110 1084.220 ;
        RECT 2280.290 1084.160 2280.610 1084.220 ;
        RECT 2268.790 1084.020 2280.610 1084.160 ;
        RECT 2268.790 1083.960 2269.110 1084.020 ;
        RECT 2280.290 1083.960 2280.610 1084.020 ;
        RECT 2280.290 324.260 2280.610 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2280.290 324.120 2899.310 324.260 ;
        RECT 2280.290 324.060 2280.610 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2268.820 1083.960 2269.080 1084.220 ;
        RECT 2280.320 1083.960 2280.580 1084.220 ;
        RECT 2280.320 324.060 2280.580 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2268.810 1084.755 2269.090 1085.125 ;
        RECT 2268.880 1084.250 2269.020 1084.755 ;
        RECT 2268.820 1083.930 2269.080 1084.250 ;
        RECT 2280.320 1083.930 2280.580 1084.250 ;
        RECT 2280.380 324.350 2280.520 1083.930 ;
        RECT 2280.320 324.030 2280.580 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2268.810 1084.800 2269.090 1085.080 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2268.785 1085.090 2269.115 1085.105 ;
        RECT 2250.780 1085.080 2269.115 1085.090 ;
        RECT 2247.465 1084.790 2269.115 1085.080 ;
        RECT 2247.465 1084.480 2251.465 1084.790 ;
        RECT 2268.785 1084.775 2269.115 1084.790 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 2577.440 1179.830 2577.500 ;
        RECT 1337.750 2577.440 1338.070 2577.500 ;
        RECT 1179.510 2577.300 1338.070 2577.440 ;
        RECT 1179.510 2577.240 1179.830 2577.300 ;
        RECT 1337.750 2577.240 1338.070 2577.300 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 2577.240 1179.800 2577.500 ;
        RECT 1337.780 2577.240 1338.040 2577.500 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2577.530 1179.740 3498.270 ;
        RECT 1179.540 2577.210 1179.800 2577.530 ;
        RECT 1337.780 2577.210 1338.040 2577.530 ;
        RECT 1337.840 2562.185 1337.980 2577.210 ;
        RECT 1337.670 2561.900 1337.980 2562.185 ;
        RECT 1337.670 2558.185 1337.950 2561.900 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 855.210 3501.220 855.530 3501.280 ;
        RECT 851.530 3501.080 855.530 3501.220 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
        RECT 855.210 3501.020 855.530 3501.080 ;
        RECT 855.210 2577.780 855.530 2577.840 ;
        RECT 1161.110 2577.780 1161.430 2577.840 ;
        RECT 855.210 2577.640 1161.430 2577.780 ;
        RECT 855.210 2577.580 855.530 2577.640 ;
        RECT 1161.110 2577.580 1161.430 2577.640 ;
      LAYER via ;
        RECT 851.560 3501.020 851.820 3501.280 ;
        RECT 855.240 3501.020 855.500 3501.280 ;
        RECT 855.240 2577.580 855.500 2577.840 ;
        RECT 1161.140 2577.580 1161.400 2577.840 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 855.240 3500.990 855.500 3501.310 ;
        RECT 855.300 2577.870 855.440 3500.990 ;
        RECT 855.240 2577.550 855.500 2577.870 ;
        RECT 1161.140 2577.550 1161.400 2577.870 ;
        RECT 1161.200 2562.185 1161.340 2577.550 ;
        RECT 1161.030 2561.900 1161.340 2562.185 ;
        RECT 1161.030 2558.185 1161.310 2561.900 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 2578.800 531.230 2578.860 ;
        RECT 984.010 2578.800 984.330 2578.860 ;
        RECT 530.910 2578.660 984.330 2578.800 ;
        RECT 530.910 2578.600 531.230 2578.660 ;
        RECT 984.010 2578.600 984.330 2578.660 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 2578.600 531.200 2578.860 ;
        RECT 984.040 2578.600 984.300 2578.860 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2578.890 531.140 3498.270 ;
        RECT 530.940 2578.570 531.200 2578.890 ;
        RECT 984.040 2578.570 984.300 2578.890 ;
        RECT 984.100 2562.185 984.240 2578.570 ;
        RECT 983.930 2561.900 984.240 2562.185 ;
        RECT 983.930 2558.185 984.210 2561.900 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 2577.780 206.930 2577.840 ;
        RECT 807.370 2577.780 807.690 2577.840 ;
        RECT 206.610 2577.640 807.690 2577.780 ;
        RECT 206.610 2577.580 206.930 2577.640 ;
        RECT 807.370 2577.580 807.690 2577.640 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 2577.580 206.900 2577.840 ;
        RECT 807.400 2577.580 807.660 2577.840 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 2577.870 206.840 3501.670 ;
        RECT 206.640 2577.550 206.900 2577.870 ;
        RECT 807.400 2577.550 807.660 2577.870 ;
        RECT 807.460 2562.185 807.600 2577.550 ;
        RECT 807.290 2561.900 807.600 2562.185 ;
        RECT 807.290 2558.185 807.570 2561.900 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 3408.740 16.950 3408.800 ;
        RECT 30.890 3408.740 31.210 3408.800 ;
        RECT 16.630 3408.600 31.210 3408.740 ;
        RECT 16.630 3408.540 16.950 3408.600 ;
        RECT 30.890 3408.540 31.210 3408.600 ;
        RECT 30.890 2546.160 31.210 2546.220 ;
        RECT 641.770 2546.160 642.090 2546.220 ;
        RECT 30.890 2546.020 642.090 2546.160 ;
        RECT 30.890 2545.960 31.210 2546.020 ;
        RECT 641.770 2545.960 642.090 2546.020 ;
      LAYER via ;
        RECT 16.660 3408.540 16.920 3408.800 ;
        RECT 30.920 3408.540 31.180 3408.800 ;
        RECT 30.920 2545.960 31.180 2546.220 ;
        RECT 641.800 2545.960 642.060 2546.220 ;
      LAYER met2 ;
        RECT 16.650 3411.035 16.930 3411.405 ;
        RECT 16.720 3408.830 16.860 3411.035 ;
        RECT 16.660 3408.510 16.920 3408.830 ;
        RECT 30.920 3408.510 31.180 3408.830 ;
        RECT 30.980 2546.250 31.120 3408.510 ;
        RECT 30.920 2545.930 31.180 2546.250 ;
        RECT 641.800 2545.930 642.060 2546.250 ;
        RECT 641.860 2543.045 642.000 2545.930 ;
        RECT 641.790 2542.675 642.070 2543.045 ;
      LAYER via2 ;
        RECT 16.650 3411.080 16.930 3411.360 ;
        RECT 641.790 2542.720 642.070 2543.000 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 16.625 3411.370 16.955 3411.385 ;
        RECT -4.800 3411.070 16.955 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 16.625 3411.055 16.955 3411.070 ;
        RECT 641.765 2543.010 642.095 2543.025 ;
        RECT 641.765 2543.000 660.100 2543.010 ;
        RECT 641.765 2542.710 664.000 2543.000 ;
        RECT 641.765 2542.695 642.095 2542.710 ;
        RECT 660.000 2542.400 664.000 2542.710 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 44.690 3119.060 45.010 3119.120 ;
        RECT 16.170 3118.920 45.010 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 44.690 3118.860 45.010 3118.920 ;
        RECT 44.690 2428.860 45.010 2428.920 ;
        RECT 641.770 2428.860 642.090 2428.920 ;
        RECT 44.690 2428.720 642.090 2428.860 ;
        RECT 44.690 2428.660 45.010 2428.720 ;
        RECT 641.770 2428.660 642.090 2428.720 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 44.720 3118.860 44.980 3119.120 ;
        RECT 44.720 2428.660 44.980 2428.920 ;
        RECT 641.800 2428.660 642.060 2428.920 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 44.720 3118.830 44.980 3119.150 ;
        RECT 44.780 2428.950 44.920 3118.830 ;
        RECT 44.720 2428.630 44.980 2428.950 ;
        RECT 641.800 2428.805 642.060 2428.950 ;
        RECT 641.790 2428.435 642.070 2428.805 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
        RECT 641.790 2428.480 642.070 2428.760 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
        RECT 641.765 2428.770 642.095 2428.785 ;
        RECT 641.765 2428.760 660.100 2428.770 ;
        RECT 641.765 2428.470 664.000 2428.760 ;
        RECT 641.765 2428.455 642.095 2428.470 ;
        RECT 660.000 2428.160 664.000 2428.470 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2836.520 20.630 2836.580 ;
        RECT 51.590 2836.520 51.910 2836.580 ;
        RECT 20.310 2836.380 51.910 2836.520 ;
        RECT 20.310 2836.320 20.630 2836.380 ;
        RECT 51.590 2836.320 51.910 2836.380 ;
        RECT 51.590 2318.360 51.910 2318.420 ;
        RECT 641.770 2318.360 642.090 2318.420 ;
        RECT 51.590 2318.220 642.090 2318.360 ;
        RECT 51.590 2318.160 51.910 2318.220 ;
        RECT 641.770 2318.160 642.090 2318.220 ;
      LAYER via ;
        RECT 20.340 2836.320 20.600 2836.580 ;
        RECT 51.620 2836.320 51.880 2836.580 ;
        RECT 51.620 2318.160 51.880 2318.420 ;
        RECT 641.800 2318.160 642.060 2318.420 ;
      LAYER met2 ;
        RECT 20.330 2836.435 20.610 2836.805 ;
        RECT 20.340 2836.290 20.600 2836.435 ;
        RECT 51.620 2836.290 51.880 2836.610 ;
        RECT 51.680 2318.450 51.820 2836.290 ;
        RECT 51.620 2318.130 51.880 2318.450 ;
        RECT 641.800 2318.130 642.060 2318.450 ;
        RECT 641.860 2314.565 642.000 2318.130 ;
        RECT 641.790 2314.195 642.070 2314.565 ;
      LAYER via2 ;
        RECT 20.330 2836.480 20.610 2836.760 ;
        RECT 641.790 2314.240 642.070 2314.520 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 20.305 2836.770 20.635 2836.785 ;
        RECT -4.800 2836.470 20.635 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 20.305 2836.455 20.635 2836.470 ;
        RECT 641.765 2314.530 642.095 2314.545 ;
        RECT 641.765 2314.520 660.100 2314.530 ;
        RECT 641.765 2314.230 664.000 2314.520 ;
        RECT 641.765 2314.215 642.095 2314.230 ;
        RECT 660.000 2313.920 664.000 2314.230 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2546.500 16.490 2546.560 ;
        RECT 37.790 2546.500 38.110 2546.560 ;
        RECT 16.170 2546.360 38.110 2546.500 ;
        RECT 16.170 2546.300 16.490 2546.360 ;
        RECT 37.790 2546.300 38.110 2546.360 ;
        RECT 37.790 2201.060 38.110 2201.120 ;
        RECT 641.770 2201.060 642.090 2201.120 ;
        RECT 37.790 2200.920 642.090 2201.060 ;
        RECT 37.790 2200.860 38.110 2200.920 ;
        RECT 641.770 2200.860 642.090 2200.920 ;
      LAYER via ;
        RECT 16.200 2546.300 16.460 2546.560 ;
        RECT 37.820 2546.300 38.080 2546.560 ;
        RECT 37.820 2200.860 38.080 2201.120 ;
        RECT 641.800 2200.860 642.060 2201.120 ;
      LAYER met2 ;
        RECT 16.190 2549.475 16.470 2549.845 ;
        RECT 16.260 2546.590 16.400 2549.475 ;
        RECT 16.200 2546.270 16.460 2546.590 ;
        RECT 37.820 2546.270 38.080 2546.590 ;
        RECT 37.880 2201.150 38.020 2546.270 ;
        RECT 37.820 2200.830 38.080 2201.150 ;
        RECT 641.800 2200.830 642.060 2201.150 ;
        RECT 641.860 2200.325 642.000 2200.830 ;
        RECT 641.790 2199.955 642.070 2200.325 ;
      LAYER via2 ;
        RECT 16.190 2549.520 16.470 2549.800 ;
        RECT 641.790 2200.000 642.070 2200.280 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.165 2549.810 16.495 2549.825 ;
        RECT -4.800 2549.510 16.495 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.165 2549.495 16.495 2549.510 ;
        RECT 641.765 2200.290 642.095 2200.305 ;
        RECT 641.765 2200.280 660.100 2200.290 ;
        RECT 641.765 2199.990 664.000 2200.280 ;
        RECT 641.765 2199.975 642.095 2199.990 ;
        RECT 660.000 2199.680 664.000 2199.990 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2090.560 17.870 2090.620 ;
        RECT 641.770 2090.560 642.090 2090.620 ;
        RECT 17.550 2090.420 642.090 2090.560 ;
        RECT 17.550 2090.360 17.870 2090.420 ;
        RECT 641.770 2090.360 642.090 2090.420 ;
      LAYER via ;
        RECT 17.580 2090.360 17.840 2090.620 ;
        RECT 641.800 2090.360 642.060 2090.620 ;
      LAYER met2 ;
        RECT 17.570 2261.835 17.850 2262.205 ;
        RECT 17.640 2090.650 17.780 2261.835 ;
        RECT 17.580 2090.330 17.840 2090.650 ;
        RECT 641.800 2090.330 642.060 2090.650 ;
        RECT 641.860 2085.405 642.000 2090.330 ;
        RECT 641.790 2085.035 642.070 2085.405 ;
      LAYER via2 ;
        RECT 17.570 2261.880 17.850 2262.160 ;
        RECT 641.790 2085.080 642.070 2085.360 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.545 2262.170 17.875 2262.185 ;
        RECT -4.800 2261.870 17.875 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.545 2261.855 17.875 2261.870 ;
        RECT 641.765 2085.370 642.095 2085.385 ;
        RECT 641.765 2085.360 660.100 2085.370 ;
        RECT 641.765 2085.070 664.000 2085.360 ;
        RECT 641.765 2085.055 642.095 2085.070 ;
        RECT 660.000 2084.760 664.000 2085.070 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1973.260 17.410 1973.320 ;
        RECT 641.770 1973.260 642.090 1973.320 ;
        RECT 17.090 1973.120 642.090 1973.260 ;
        RECT 17.090 1973.060 17.410 1973.120 ;
        RECT 641.770 1973.060 642.090 1973.120 ;
      LAYER via ;
        RECT 17.120 1973.060 17.380 1973.320 ;
        RECT 641.800 1973.060 642.060 1973.320 ;
      LAYER met2 ;
        RECT 17.110 1974.875 17.390 1975.245 ;
        RECT 17.180 1973.350 17.320 1974.875 ;
        RECT 17.120 1973.030 17.380 1973.350 ;
        RECT 641.800 1973.030 642.060 1973.350 ;
        RECT 641.860 1971.165 642.000 1973.030 ;
        RECT 641.790 1970.795 642.070 1971.165 ;
      LAYER via2 ;
        RECT 17.110 1974.920 17.390 1975.200 ;
        RECT 641.790 1970.840 642.070 1971.120 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 17.085 1975.210 17.415 1975.225 ;
        RECT -4.800 1974.910 17.415 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 17.085 1974.895 17.415 1974.910 ;
        RECT 641.765 1971.130 642.095 1971.145 ;
        RECT 641.765 1971.120 660.100 1971.130 ;
        RECT 641.765 1970.830 664.000 1971.120 ;
        RECT 641.765 1970.815 642.095 1970.830 ;
        RECT 660.000 1970.520 664.000 1970.830 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1187.180 2270.030 1187.240 ;
        RECT 2349.290 1187.180 2349.610 1187.240 ;
        RECT 2269.710 1187.040 2349.610 1187.180 ;
        RECT 2269.710 1186.980 2270.030 1187.040 ;
        RECT 2349.290 1186.980 2349.610 1187.040 ;
        RECT 2349.290 558.860 2349.610 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2349.290 558.720 2899.310 558.860 ;
        RECT 2349.290 558.660 2349.610 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2269.740 1186.980 2270.000 1187.240 ;
        RECT 2349.320 1186.980 2349.580 1187.240 ;
        RECT 2349.320 558.660 2349.580 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2269.730 1191.515 2270.010 1191.885 ;
        RECT 2269.800 1187.270 2269.940 1191.515 ;
        RECT 2269.740 1186.950 2270.000 1187.270 ;
        RECT 2349.320 1186.950 2349.580 1187.270 ;
        RECT 2349.380 558.950 2349.520 1186.950 ;
        RECT 2349.320 558.630 2349.580 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2269.730 1191.560 2270.010 1191.840 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2269.705 1191.850 2270.035 1191.865 ;
        RECT 2250.780 1191.840 2270.035 1191.850 ;
        RECT 2247.465 1191.550 2270.035 1191.840 ;
        RECT 2247.465 1191.240 2251.465 1191.550 ;
        RECT 2269.705 1191.535 2270.035 1191.550 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 1690.380 17.870 1690.440 ;
        RECT 646.370 1690.380 646.690 1690.440 ;
        RECT 17.550 1690.240 646.690 1690.380 ;
        RECT 17.550 1690.180 17.870 1690.240 ;
        RECT 646.370 1690.180 646.690 1690.240 ;
      LAYER via ;
        RECT 17.580 1690.180 17.840 1690.440 ;
        RECT 646.400 1690.180 646.660 1690.440 ;
      LAYER met2 ;
        RECT 646.390 1856.555 646.670 1856.925 ;
        RECT 646.460 1690.470 646.600 1856.555 ;
        RECT 17.580 1690.150 17.840 1690.470 ;
        RECT 646.400 1690.150 646.660 1690.470 ;
        RECT 17.640 1687.605 17.780 1690.150 ;
        RECT 17.570 1687.235 17.850 1687.605 ;
      LAYER via2 ;
        RECT 646.390 1856.600 646.670 1856.880 ;
        RECT 17.570 1687.280 17.850 1687.560 ;
      LAYER met3 ;
        RECT 646.365 1856.890 646.695 1856.905 ;
        RECT 646.365 1856.880 660.100 1856.890 ;
        RECT 646.365 1856.590 664.000 1856.880 ;
        RECT 646.365 1856.575 646.695 1856.590 ;
        RECT 660.000 1856.280 664.000 1856.590 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.545 1687.570 17.875 1687.585 ;
        RECT -4.800 1687.270 17.875 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.545 1687.255 17.875 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1739.000 17.410 1739.060 ;
        RECT 641.770 1739.000 642.090 1739.060 ;
        RECT 17.090 1738.860 642.090 1739.000 ;
        RECT 17.090 1738.800 17.410 1738.860 ;
        RECT 641.770 1738.800 642.090 1738.860 ;
      LAYER via ;
        RECT 17.120 1738.800 17.380 1739.060 ;
        RECT 641.800 1738.800 642.060 1739.060 ;
      LAYER met2 ;
        RECT 641.790 1741.635 642.070 1742.005 ;
        RECT 641.860 1739.090 642.000 1741.635 ;
        RECT 17.120 1738.770 17.380 1739.090 ;
        RECT 641.800 1738.770 642.060 1739.090 ;
        RECT 17.180 1472.045 17.320 1738.770 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 641.790 1741.680 642.070 1741.960 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 641.765 1741.970 642.095 1741.985 ;
        RECT 641.765 1741.960 660.100 1741.970 ;
        RECT 641.765 1741.670 664.000 1741.960 ;
        RECT 641.765 1741.655 642.095 1741.670 ;
        RECT 660.000 1741.360 664.000 1741.670 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 1621.700 38.110 1621.760 ;
        RECT 641.770 1621.700 642.090 1621.760 ;
        RECT 37.790 1621.560 642.090 1621.700 ;
        RECT 37.790 1621.500 38.110 1621.560 ;
        RECT 641.770 1621.500 642.090 1621.560 ;
        RECT 17.550 1258.240 17.870 1258.300 ;
        RECT 37.790 1258.240 38.110 1258.300 ;
        RECT 17.550 1258.100 38.110 1258.240 ;
        RECT 17.550 1258.040 17.870 1258.100 ;
        RECT 37.790 1258.040 38.110 1258.100 ;
      LAYER via ;
        RECT 37.820 1621.500 38.080 1621.760 ;
        RECT 641.800 1621.500 642.060 1621.760 ;
        RECT 17.580 1258.040 17.840 1258.300 ;
        RECT 37.820 1258.040 38.080 1258.300 ;
      LAYER met2 ;
        RECT 641.790 1627.395 642.070 1627.765 ;
        RECT 641.860 1621.790 642.000 1627.395 ;
        RECT 37.820 1621.470 38.080 1621.790 ;
        RECT 641.800 1621.470 642.060 1621.790 ;
        RECT 37.880 1258.330 38.020 1621.470 ;
        RECT 17.580 1258.010 17.840 1258.330 ;
        RECT 37.820 1258.010 38.080 1258.330 ;
        RECT 17.640 1256.485 17.780 1258.010 ;
        RECT 17.570 1256.115 17.850 1256.485 ;
      LAYER via2 ;
        RECT 641.790 1627.440 642.070 1627.720 ;
        RECT 17.570 1256.160 17.850 1256.440 ;
      LAYER met3 ;
        RECT 641.765 1627.730 642.095 1627.745 ;
        RECT 641.765 1627.720 660.100 1627.730 ;
        RECT 641.765 1627.430 664.000 1627.720 ;
        RECT 641.765 1627.415 642.095 1627.430 ;
        RECT 660.000 1627.120 664.000 1627.430 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.545 1256.450 17.875 1256.465 ;
        RECT -4.800 1256.150 17.875 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.545 1256.135 17.875 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 30.890 1511.200 31.210 1511.260 ;
        RECT 641.770 1511.200 642.090 1511.260 ;
        RECT 30.890 1511.060 642.090 1511.200 ;
        RECT 30.890 1511.000 31.210 1511.060 ;
        RECT 641.770 1511.000 642.090 1511.060 ;
        RECT 15.710 1040.980 16.030 1041.040 ;
        RECT 30.890 1040.980 31.210 1041.040 ;
        RECT 15.710 1040.840 31.210 1040.980 ;
        RECT 15.710 1040.780 16.030 1040.840 ;
        RECT 30.890 1040.780 31.210 1040.840 ;
      LAYER via ;
        RECT 30.920 1511.000 31.180 1511.260 ;
        RECT 641.800 1511.000 642.060 1511.260 ;
        RECT 15.740 1040.780 16.000 1041.040 ;
        RECT 30.920 1040.780 31.180 1041.040 ;
      LAYER met2 ;
        RECT 641.790 1513.155 642.070 1513.525 ;
        RECT 641.860 1511.290 642.000 1513.155 ;
        RECT 30.920 1510.970 31.180 1511.290 ;
        RECT 641.800 1510.970 642.060 1511.290 ;
        RECT 30.980 1041.070 31.120 1510.970 ;
        RECT 15.740 1040.925 16.000 1041.070 ;
        RECT 15.730 1040.555 16.010 1040.925 ;
        RECT 30.920 1040.750 31.180 1041.070 ;
      LAYER via2 ;
        RECT 641.790 1513.200 642.070 1513.480 ;
        RECT 15.730 1040.600 16.010 1040.880 ;
      LAYER met3 ;
        RECT 641.765 1513.490 642.095 1513.505 ;
        RECT 641.765 1513.480 660.100 1513.490 ;
        RECT 641.765 1513.190 664.000 1513.480 ;
        RECT 641.765 1513.175 642.095 1513.190 ;
        RECT 660.000 1512.880 664.000 1513.190 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 15.705 1040.890 16.035 1040.905 ;
        RECT -4.800 1040.590 16.035 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 15.705 1040.575 16.035 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1390.160 17.410 1390.220 ;
        RECT 641.310 1390.160 641.630 1390.220 ;
        RECT 17.090 1390.020 641.630 1390.160 ;
        RECT 17.090 1389.960 17.410 1390.020 ;
        RECT 641.310 1389.960 641.630 1390.020 ;
      LAYER via ;
        RECT 17.120 1389.960 17.380 1390.220 ;
        RECT 641.340 1389.960 641.600 1390.220 ;
      LAYER met2 ;
        RECT 641.330 1398.915 641.610 1399.285 ;
        RECT 641.400 1390.250 641.540 1398.915 ;
        RECT 17.120 1389.930 17.380 1390.250 ;
        RECT 641.340 1389.930 641.600 1390.250 ;
        RECT 17.180 825.365 17.320 1389.930 ;
        RECT 17.110 824.995 17.390 825.365 ;
      LAYER via2 ;
        RECT 641.330 1398.960 641.610 1399.240 ;
        RECT 17.110 825.040 17.390 825.320 ;
      LAYER met3 ;
        RECT 641.305 1399.250 641.635 1399.265 ;
        RECT 641.305 1399.240 660.100 1399.250 ;
        RECT 641.305 1398.950 664.000 1399.240 ;
        RECT 641.305 1398.935 641.635 1398.950 ;
        RECT 660.000 1398.640 664.000 1398.950 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.085 825.330 17.415 825.345 ;
        RECT -4.800 825.030 17.415 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.085 825.015 17.415 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 1283.740 51.910 1283.800 ;
        RECT 641.770 1283.740 642.090 1283.800 ;
        RECT 51.590 1283.600 642.090 1283.740 ;
        RECT 51.590 1283.540 51.910 1283.600 ;
        RECT 641.770 1283.540 642.090 1283.600 ;
        RECT 17.090 613.940 17.410 614.000 ;
        RECT 51.590 613.940 51.910 614.000 ;
        RECT 17.090 613.800 51.910 613.940 ;
        RECT 17.090 613.740 17.410 613.800 ;
        RECT 51.590 613.740 51.910 613.800 ;
      LAYER via ;
        RECT 51.620 1283.540 51.880 1283.800 ;
        RECT 641.800 1283.540 642.060 1283.800 ;
        RECT 17.120 613.740 17.380 614.000 ;
        RECT 51.620 613.740 51.880 614.000 ;
      LAYER met2 ;
        RECT 641.790 1283.995 642.070 1284.365 ;
        RECT 641.860 1283.830 642.000 1283.995 ;
        RECT 51.620 1283.510 51.880 1283.830 ;
        RECT 641.800 1283.510 642.060 1283.830 ;
        RECT 51.680 614.030 51.820 1283.510 ;
        RECT 17.120 613.710 17.380 614.030 ;
        RECT 51.620 613.710 51.880 614.030 ;
        RECT 17.180 610.485 17.320 613.710 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 641.790 1284.040 642.070 1284.320 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 641.765 1284.330 642.095 1284.345 ;
        RECT 641.765 1284.320 660.100 1284.330 ;
        RECT 641.765 1284.030 664.000 1284.320 ;
        RECT 641.765 1284.015 642.095 1284.030 ;
        RECT 660.000 1283.720 664.000 1284.030 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 72.290 1166.440 72.610 1166.500 ;
        RECT 641.770 1166.440 642.090 1166.500 ;
        RECT 72.290 1166.300 642.090 1166.440 ;
        RECT 72.290 1166.240 72.610 1166.300 ;
        RECT 641.770 1166.240 642.090 1166.300 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 72.290 400.080 72.610 400.140 ;
        RECT 17.090 399.940 72.610 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 72.290 399.880 72.610 399.940 ;
      LAYER via ;
        RECT 72.320 1166.240 72.580 1166.500 ;
        RECT 641.800 1166.240 642.060 1166.500 ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 72.320 399.880 72.580 400.140 ;
      LAYER met2 ;
        RECT 641.790 1169.755 642.070 1170.125 ;
        RECT 641.860 1166.530 642.000 1169.755 ;
        RECT 72.320 1166.210 72.580 1166.530 ;
        RECT 641.800 1166.210 642.060 1166.530 ;
        RECT 72.380 400.170 72.520 1166.210 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 72.320 399.850 72.580 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 641.790 1169.800 642.070 1170.080 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 641.765 1170.090 642.095 1170.105 ;
        RECT 641.765 1170.080 660.100 1170.090 ;
        RECT 641.765 1169.790 664.000 1170.080 ;
        RECT 641.765 1169.775 642.095 1169.790 ;
        RECT 660.000 1169.480 664.000 1169.790 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 1055.940 38.110 1056.000 ;
        RECT 641.770 1055.940 642.090 1056.000 ;
        RECT 37.790 1055.800 642.090 1055.940 ;
        RECT 37.790 1055.740 38.110 1055.800 ;
        RECT 641.770 1055.740 642.090 1055.800 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 37.790 179.420 38.110 179.480 ;
        RECT 17.090 179.280 38.110 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 37.790 179.220 38.110 179.280 ;
      LAYER via ;
        RECT 37.820 1055.740 38.080 1056.000 ;
        RECT 641.800 1055.740 642.060 1056.000 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 37.820 179.220 38.080 179.480 ;
      LAYER met2 ;
        RECT 37.820 1055.710 38.080 1056.030 ;
        RECT 641.800 1055.885 642.060 1056.030 ;
        RECT 37.880 179.510 38.020 1055.710 ;
        RECT 641.790 1055.515 642.070 1055.885 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 37.820 179.190 38.080 179.510 ;
      LAYER via2 ;
        RECT 641.790 1055.560 642.070 1055.840 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 641.765 1055.850 642.095 1055.865 ;
        RECT 641.765 1055.840 660.100 1055.850 ;
        RECT 641.765 1055.550 664.000 1055.840 ;
        RECT 641.765 1055.535 642.095 1055.550 ;
        RECT 660.000 1055.240 664.000 1055.550 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1297.340 2270.030 1297.400 ;
        RECT 2356.190 1297.340 2356.510 1297.400 ;
        RECT 2269.710 1297.200 2356.510 1297.340 ;
        RECT 2269.710 1297.140 2270.030 1297.200 ;
        RECT 2356.190 1297.140 2356.510 1297.200 ;
        RECT 2356.190 793.460 2356.510 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2356.190 793.320 2899.310 793.460 ;
        RECT 2356.190 793.260 2356.510 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2269.740 1297.140 2270.000 1297.400 ;
        RECT 2356.220 1297.140 2356.480 1297.400 ;
        RECT 2356.220 793.260 2356.480 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2269.730 1298.275 2270.010 1298.645 ;
        RECT 2269.800 1297.430 2269.940 1298.275 ;
        RECT 2269.740 1297.110 2270.000 1297.430 ;
        RECT 2356.220 1297.110 2356.480 1297.430 ;
        RECT 2356.280 793.550 2356.420 1297.110 ;
        RECT 2356.220 793.230 2356.480 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2269.730 1298.320 2270.010 1298.600 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2269.705 1298.610 2270.035 1298.625 ;
        RECT 2250.780 1298.600 2270.035 1298.610 ;
        RECT 2247.465 1298.310 2270.035 1298.600 ;
        RECT 2247.465 1298.000 2251.465 1298.310 ;
        RECT 2269.705 1298.295 2270.035 1298.310 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1401.040 2270.030 1401.100 ;
        RECT 2307.890 1401.040 2308.210 1401.100 ;
        RECT 2269.710 1400.900 2308.210 1401.040 ;
        RECT 2269.710 1400.840 2270.030 1400.900 ;
        RECT 2307.890 1400.840 2308.210 1400.900 ;
        RECT 2307.890 1028.060 2308.210 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2307.890 1027.920 2899.310 1028.060 ;
        RECT 2307.890 1027.860 2308.210 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2269.740 1400.840 2270.000 1401.100 ;
        RECT 2307.920 1400.840 2308.180 1401.100 ;
        RECT 2307.920 1027.860 2308.180 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2269.730 1405.035 2270.010 1405.405 ;
        RECT 2269.800 1401.130 2269.940 1405.035 ;
        RECT 2269.740 1400.810 2270.000 1401.130 ;
        RECT 2307.920 1400.810 2308.180 1401.130 ;
        RECT 2307.980 1028.150 2308.120 1400.810 ;
        RECT 2307.920 1027.830 2308.180 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2269.730 1405.080 2270.010 1405.360 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2269.705 1405.370 2270.035 1405.385 ;
        RECT 2250.780 1405.360 2270.035 1405.370 ;
        RECT 2247.465 1405.070 2270.035 1405.360 ;
        RECT 2247.465 1404.760 2251.465 1405.070 ;
        RECT 2269.705 1405.055 2270.035 1405.070 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2268.330 1511.880 2268.650 1511.940 ;
        RECT 2280.290 1511.880 2280.610 1511.940 ;
        RECT 2268.330 1511.740 2280.610 1511.880 ;
        RECT 2268.330 1511.680 2268.650 1511.740 ;
        RECT 2280.290 1511.680 2280.610 1511.740 ;
        RECT 2280.290 1262.660 2280.610 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2280.290 1262.520 2899.310 1262.660 ;
        RECT 2280.290 1262.460 2280.610 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2268.360 1511.680 2268.620 1511.940 ;
        RECT 2280.320 1511.680 2280.580 1511.940 ;
        RECT 2280.320 1262.460 2280.580 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2268.350 1511.795 2268.630 1512.165 ;
        RECT 2268.360 1511.650 2268.620 1511.795 ;
        RECT 2280.320 1511.650 2280.580 1511.970 ;
        RECT 2280.380 1262.750 2280.520 1511.650 ;
        RECT 2280.320 1262.430 2280.580 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2268.350 1511.840 2268.630 1512.120 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2268.325 1512.130 2268.655 1512.145 ;
        RECT 2250.780 1512.120 2268.655 1512.130 ;
        RECT 2247.465 1511.830 2268.655 1512.120 ;
        RECT 2247.465 1511.520 2251.465 1511.830 ;
        RECT 2268.325 1511.815 2268.655 1511.830 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.490 1497.260 2266.810 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 2266.490 1497.120 2899.310 1497.260 ;
        RECT 2266.490 1497.060 2266.810 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 2266.520 1497.060 2266.780 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 2266.510 1618.555 2266.790 1618.925 ;
        RECT 2266.580 1497.350 2266.720 1618.555 ;
        RECT 2266.520 1497.030 2266.780 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2266.510 1618.600 2266.790 1618.880 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2266.485 1618.890 2266.815 1618.905 ;
        RECT 2250.780 1618.880 2266.815 1618.890 ;
        RECT 2247.465 1618.590 2266.815 1618.880 ;
        RECT 2247.465 1618.280 2251.465 1618.590 ;
        RECT 2266.485 1618.575 2266.815 1618.590 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1728.460 2270.030 1728.520 ;
        RECT 2900.830 1728.460 2901.150 1728.520 ;
        RECT 2269.710 1728.320 2901.150 1728.460 ;
        RECT 2269.710 1728.260 2270.030 1728.320 ;
        RECT 2900.830 1728.260 2901.150 1728.320 ;
      LAYER via ;
        RECT 2269.740 1728.260 2270.000 1728.520 ;
        RECT 2900.860 1728.260 2901.120 1728.520 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1728.550 2901.060 1730.075 ;
        RECT 2269.740 1728.230 2270.000 1728.550 ;
        RECT 2900.860 1728.230 2901.120 1728.550 ;
        RECT 2269.800 1725.685 2269.940 1728.230 ;
        RECT 2269.730 1725.315 2270.010 1725.685 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 2269.730 1725.360 2270.010 1725.640 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2269.705 1725.650 2270.035 1725.665 ;
        RECT 2250.780 1725.640 2270.035 1725.650 ;
        RECT 2247.465 1725.350 2270.035 1725.640 ;
        RECT 2247.465 1725.040 2251.465 1725.350 ;
        RECT 2269.705 1725.335 2270.035 1725.350 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2300.990 1960.000 2301.310 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2300.990 1959.860 2901.150 1960.000 ;
        RECT 2300.990 1959.800 2301.310 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
        RECT 2269.710 1833.520 2270.030 1833.580 ;
        RECT 2300.990 1833.520 2301.310 1833.580 ;
        RECT 2269.710 1833.380 2301.310 1833.520 ;
        RECT 2269.710 1833.320 2270.030 1833.380 ;
        RECT 2300.990 1833.320 2301.310 1833.380 ;
      LAYER via ;
        RECT 2301.020 1959.800 2301.280 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
        RECT 2269.740 1833.320 2270.000 1833.580 ;
        RECT 2301.020 1833.320 2301.280 1833.580 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2301.020 1959.770 2301.280 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2301.080 1833.610 2301.220 1959.770 ;
        RECT 2269.740 1833.290 2270.000 1833.610 ;
        RECT 2301.020 1833.290 2301.280 1833.610 ;
        RECT 2269.800 1832.445 2269.940 1833.290 ;
        RECT 2269.730 1832.075 2270.010 1832.445 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2269.730 1832.120 2270.010 1832.400 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2269.705 1832.410 2270.035 1832.425 ;
        RECT 2250.780 1832.400 2270.035 1832.410 ;
        RECT 2247.465 1832.110 2270.035 1832.400 ;
        RECT 2247.465 1831.800 2251.465 1832.110 ;
        RECT 2269.705 1832.095 2270.035 1832.110 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.490 2194.600 2266.810 2194.660 ;
        RECT 2899.450 2194.600 2899.770 2194.660 ;
        RECT 2266.490 2194.460 2899.770 2194.600 ;
        RECT 2266.490 2194.400 2266.810 2194.460 ;
        RECT 2899.450 2194.400 2899.770 2194.460 ;
      LAYER via ;
        RECT 2266.520 2194.400 2266.780 2194.660 ;
        RECT 2899.480 2194.400 2899.740 2194.660 ;
      LAYER met2 ;
        RECT 2899.470 2199.275 2899.750 2199.645 ;
        RECT 2899.540 2194.690 2899.680 2199.275 ;
        RECT 2266.520 2194.370 2266.780 2194.690 ;
        RECT 2899.480 2194.370 2899.740 2194.690 ;
        RECT 2266.580 1939.205 2266.720 2194.370 ;
        RECT 2266.510 1938.835 2266.790 1939.205 ;
      LAYER via2 ;
        RECT 2899.470 2199.320 2899.750 2199.600 ;
        RECT 2266.510 1938.880 2266.790 1939.160 ;
      LAYER met3 ;
        RECT 2899.445 2199.610 2899.775 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2899.445 2199.310 2924.800 2199.610 ;
        RECT 2899.445 2199.295 2899.775 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2266.485 1939.170 2266.815 1939.185 ;
        RECT 2250.780 1939.160 2266.815 1939.170 ;
        RECT 2247.465 1938.870 2266.815 1939.160 ;
        RECT 2247.465 1938.560 2251.465 1938.870 ;
        RECT 2266.485 1938.855 2266.815 1938.870 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1049.140 2270.030 1049.200 ;
        RECT 2390.690 1049.140 2391.010 1049.200 ;
        RECT 2269.710 1049.000 2391.010 1049.140 ;
        RECT 2269.710 1048.940 2270.030 1049.000 ;
        RECT 2390.690 1048.940 2391.010 1049.000 ;
        RECT 2390.690 206.960 2391.010 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2390.690 206.820 2901.150 206.960 ;
        RECT 2390.690 206.760 2391.010 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2269.740 1048.940 2270.000 1049.200 ;
        RECT 2390.720 1048.940 2390.980 1049.200 ;
        RECT 2390.720 206.760 2390.980 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2269.740 1049.085 2270.000 1049.230 ;
        RECT 2269.730 1048.715 2270.010 1049.085 ;
        RECT 2390.720 1048.910 2390.980 1049.230 ;
        RECT 2390.780 207.050 2390.920 1048.910 ;
        RECT 2390.720 206.730 2390.980 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2269.730 1048.760 2270.010 1049.040 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2269.705 1049.050 2270.035 1049.065 ;
        RECT 2250.780 1049.040 2270.035 1049.050 ;
        RECT 2247.465 1048.750 2270.035 1049.040 ;
        RECT 2247.465 1048.440 2251.465 1048.750 ;
        RECT 2269.705 1048.735 2270.035 1048.750 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2314.790 2546.500 2315.110 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2314.790 2546.360 2901.150 2546.500 ;
        RECT 2314.790 2546.300 2315.110 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
        RECT 2269.710 2118.100 2270.030 2118.160 ;
        RECT 2314.790 2118.100 2315.110 2118.160 ;
        RECT 2269.710 2117.960 2315.110 2118.100 ;
        RECT 2269.710 2117.900 2270.030 2117.960 ;
        RECT 2314.790 2117.900 2315.110 2117.960 ;
      LAYER via ;
        RECT 2314.820 2546.300 2315.080 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
        RECT 2269.740 2117.900 2270.000 2118.160 ;
        RECT 2314.820 2117.900 2315.080 2118.160 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2314.820 2546.270 2315.080 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2314.880 2118.190 2315.020 2546.270 ;
        RECT 2269.740 2117.870 2270.000 2118.190 ;
        RECT 2314.820 2117.870 2315.080 2118.190 ;
        RECT 2269.800 2117.365 2269.940 2117.870 ;
        RECT 2269.730 2116.995 2270.010 2117.365 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2269.730 2117.040 2270.010 2117.320 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2269.705 2117.330 2270.035 2117.345 ;
        RECT 2250.780 2117.320 2270.035 2117.330 ;
        RECT 2247.465 2117.030 2270.035 2117.320 ;
        RECT 2247.465 2116.720 2251.465 2117.030 ;
        RECT 2269.705 2117.015 2270.035 2117.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2335.490 2781.100 2335.810 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2335.490 2780.960 2901.150 2781.100 ;
        RECT 2335.490 2780.900 2335.810 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2268.330 2228.600 2268.650 2228.660 ;
        RECT 2335.490 2228.600 2335.810 2228.660 ;
        RECT 2268.330 2228.460 2335.810 2228.600 ;
        RECT 2268.330 2228.400 2268.650 2228.460 ;
        RECT 2335.490 2228.400 2335.810 2228.460 ;
      LAYER via ;
        RECT 2335.520 2780.900 2335.780 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2268.360 2228.400 2268.620 2228.660 ;
        RECT 2335.520 2228.400 2335.780 2228.660 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2335.520 2780.870 2335.780 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2335.580 2228.690 2335.720 2780.870 ;
        RECT 2268.360 2228.370 2268.620 2228.690 ;
        RECT 2335.520 2228.370 2335.780 2228.690 ;
        RECT 2268.420 2224.125 2268.560 2228.370 ;
        RECT 2268.350 2223.755 2268.630 2224.125 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2268.350 2223.800 2268.630 2224.080 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2268.325 2224.090 2268.655 2224.105 ;
        RECT 2250.780 2224.080 2268.655 2224.090 ;
        RECT 2247.465 2223.790 2268.655 2224.080 ;
        RECT 2247.465 2223.480 2251.465 2223.790 ;
        RECT 2268.325 2223.775 2268.655 2223.790 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2356.190 3015.700 2356.510 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2356.190 3015.560 2901.150 3015.700 ;
        RECT 2356.190 3015.500 2356.510 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2263.730 2331.960 2264.050 2332.020 ;
        RECT 2356.190 2331.960 2356.510 2332.020 ;
        RECT 2263.730 2331.820 2356.510 2331.960 ;
        RECT 2263.730 2331.760 2264.050 2331.820 ;
        RECT 2356.190 2331.760 2356.510 2331.820 ;
      LAYER via ;
        RECT 2356.220 3015.500 2356.480 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2263.760 2331.760 2264.020 2332.020 ;
        RECT 2356.220 2331.760 2356.480 2332.020 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2356.220 3015.470 2356.480 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2356.280 2332.050 2356.420 3015.470 ;
        RECT 2263.760 2331.730 2264.020 2332.050 ;
        RECT 2356.220 2331.730 2356.480 2332.050 ;
        RECT 2263.820 2330.885 2263.960 2331.730 ;
        RECT 2263.750 2330.515 2264.030 2330.885 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2263.750 2330.560 2264.030 2330.840 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2263.725 2330.850 2264.055 2330.865 ;
        RECT 2250.780 2330.840 2264.055 2330.850 ;
        RECT 2247.465 2330.550 2264.055 2330.840 ;
        RECT 2247.465 2330.240 2251.465 2330.550 ;
        RECT 2263.725 2330.535 2264.055 2330.550 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2376.890 3250.300 2377.210 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2376.890 3250.160 2901.150 3250.300 ;
        RECT 2376.890 3250.100 2377.210 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2268.790 2442.460 2269.110 2442.520 ;
        RECT 2376.890 2442.460 2377.210 2442.520 ;
        RECT 2268.790 2442.320 2377.210 2442.460 ;
        RECT 2268.790 2442.260 2269.110 2442.320 ;
        RECT 2376.890 2442.260 2377.210 2442.320 ;
      LAYER via ;
        RECT 2376.920 3250.100 2377.180 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2268.820 2442.260 2269.080 2442.520 ;
        RECT 2376.920 2442.260 2377.180 2442.520 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2376.920 3250.070 2377.180 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2376.980 2442.550 2377.120 3250.070 ;
        RECT 2268.820 2442.230 2269.080 2442.550 ;
        RECT 2376.920 2442.230 2377.180 2442.550 ;
        RECT 2268.880 2437.645 2269.020 2442.230 ;
        RECT 2268.810 2437.275 2269.090 2437.645 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2268.810 2437.320 2269.090 2437.600 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2268.785 2437.610 2269.115 2437.625 ;
        RECT 2250.780 2437.600 2269.115 2437.610 ;
        RECT 2247.465 2437.310 2269.115 2437.600 ;
        RECT 2247.465 2437.000 2251.465 2437.310 ;
        RECT 2268.785 2437.295 2269.115 2437.310 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2383.790 3484.900 2384.110 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2383.790 3484.760 2901.150 3484.900 ;
        RECT 2383.790 3484.700 2384.110 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2266.030 2546.160 2266.350 2546.220 ;
        RECT 2383.790 2546.160 2384.110 2546.220 ;
        RECT 2266.030 2546.020 2384.110 2546.160 ;
        RECT 2266.030 2545.960 2266.350 2546.020 ;
        RECT 2383.790 2545.960 2384.110 2546.020 ;
      LAYER via ;
        RECT 2383.820 3484.700 2384.080 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2266.060 2545.960 2266.320 2546.220 ;
        RECT 2383.820 2545.960 2384.080 2546.220 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2383.820 3484.670 2384.080 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2383.880 2546.250 2384.020 3484.670 ;
        RECT 2266.060 2545.930 2266.320 2546.250 ;
        RECT 2383.820 2545.930 2384.080 2546.250 ;
        RECT 2266.120 2544.405 2266.260 2545.930 ;
        RECT 2266.050 2544.035 2266.330 2544.405 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2266.050 2544.080 2266.330 2544.360 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2266.025 2544.370 2266.355 2544.385 ;
        RECT 2250.780 2544.360 2266.355 2544.370 ;
        RECT 2247.465 2544.070 2266.355 2544.360 ;
        RECT 2247.465 2543.760 2251.465 2544.070 ;
        RECT 2266.025 2544.055 2266.355 2544.070 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.110 2577.780 2104.430 2577.840 ;
        RECT 2635.870 2577.780 2636.190 2577.840 ;
        RECT 2104.110 2577.640 2636.190 2577.780 ;
        RECT 2104.110 2577.580 2104.430 2577.640 ;
        RECT 2635.870 2577.580 2636.190 2577.640 ;
      LAYER via ;
        RECT 2104.140 2577.580 2104.400 2577.840 ;
        RECT 2635.900 2577.580 2636.160 2577.840 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 2577.870 2636.100 3517.600 ;
        RECT 2104.140 2577.550 2104.400 2577.870 ;
        RECT 2635.900 2577.550 2636.160 2577.870 ;
        RECT 2104.200 2562.185 2104.340 2577.550 ;
        RECT 2104.030 2561.900 2104.340 2562.185 ;
        RECT 2104.030 2558.185 2104.310 2561.900 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1927.470 2578.800 1927.790 2578.860 ;
        RECT 2311.570 2578.800 2311.890 2578.860 ;
        RECT 1927.470 2578.660 2311.890 2578.800 ;
        RECT 1927.470 2578.600 1927.790 2578.660 ;
        RECT 2311.570 2578.600 2311.890 2578.660 ;
      LAYER via ;
        RECT 1927.500 2578.600 1927.760 2578.860 ;
        RECT 2311.600 2578.600 2311.860 2578.860 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 2578.890 2311.800 3517.600 ;
        RECT 1927.500 2578.570 1927.760 2578.890 ;
        RECT 2311.600 2578.570 2311.860 2578.890 ;
        RECT 1927.560 2562.185 1927.700 2578.570 ;
        RECT 1927.390 2561.900 1927.700 2562.185 ;
        RECT 1927.390 2558.185 1927.670 2561.900 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1750.370 2577.780 1750.690 2577.840 ;
        RECT 1987.270 2577.780 1987.590 2577.840 ;
        RECT 1750.370 2577.640 1987.590 2577.780 ;
        RECT 1750.370 2577.580 1750.690 2577.640 ;
        RECT 1987.270 2577.580 1987.590 2577.640 ;
      LAYER via ;
        RECT 1750.400 2577.580 1750.660 2577.840 ;
        RECT 1987.300 2577.580 1987.560 2577.840 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 2577.870 1987.500 3517.600 ;
        RECT 1750.400 2577.550 1750.660 2577.870 ;
        RECT 1987.300 2577.550 1987.560 2577.870 ;
        RECT 1750.460 2562.185 1750.600 2577.550 ;
        RECT 1750.290 2561.900 1750.600 2562.185 ;
        RECT 1750.290 2558.185 1750.570 2561.900 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.070 3487.960 1656.390 3488.020 ;
        RECT 1662.510 3487.960 1662.830 3488.020 ;
        RECT 1656.070 3487.820 1662.830 3487.960 ;
        RECT 1656.070 3487.760 1656.390 3487.820 ;
        RECT 1662.510 3487.760 1662.830 3487.820 ;
        RECT 1573.730 2577.100 1574.050 2577.160 ;
        RECT 1656.070 2577.100 1656.390 2577.160 ;
        RECT 1573.730 2576.960 1656.390 2577.100 ;
        RECT 1573.730 2576.900 1574.050 2576.960 ;
        RECT 1656.070 2576.900 1656.390 2576.960 ;
      LAYER via ;
        RECT 1656.100 3487.760 1656.360 3488.020 ;
        RECT 1662.540 3487.760 1662.800 3488.020 ;
        RECT 1573.760 2576.900 1574.020 2577.160 ;
        RECT 1656.100 2576.900 1656.360 2577.160 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3488.050 1662.740 3517.600 ;
        RECT 1656.100 3487.730 1656.360 3488.050 ;
        RECT 1662.540 3487.730 1662.800 3488.050 ;
        RECT 1656.160 2577.190 1656.300 3487.730 ;
        RECT 1573.760 2576.870 1574.020 2577.190 ;
        RECT 1656.100 2576.870 1656.360 2577.190 ;
        RECT 1573.820 2562.185 1573.960 2576.870 ;
        RECT 1573.650 2561.900 1573.960 2562.185 ;
        RECT 1573.650 2558.185 1573.930 2561.900 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 2577.100 1338.530 2577.160 ;
        RECT 1396.630 2577.100 1396.950 2577.160 ;
        RECT 1338.210 2576.960 1396.950 2577.100 ;
        RECT 1338.210 2576.900 1338.530 2576.960 ;
        RECT 1396.630 2576.900 1396.950 2576.960 ;
      LAYER via ;
        RECT 1338.240 2576.900 1338.500 2577.160 ;
        RECT 1396.660 2576.900 1396.920 2577.160 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 2577.190 1338.440 3517.600 ;
        RECT 1338.240 2576.870 1338.500 2577.190 ;
        RECT 1396.660 2576.870 1396.920 2577.190 ;
        RECT 1396.720 2562.185 1396.860 2576.870 ;
        RECT 1396.550 2561.900 1396.860 2562.185 ;
        RECT 1396.550 2558.185 1396.830 2561.900 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2265.570 1152.500 2265.890 1152.560 ;
        RECT 2369.990 1152.500 2370.310 1152.560 ;
        RECT 2265.570 1152.360 2370.310 1152.500 ;
        RECT 2265.570 1152.300 2265.890 1152.360 ;
        RECT 2369.990 1152.300 2370.310 1152.360 ;
        RECT 2369.990 441.560 2370.310 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2369.990 441.420 2901.150 441.560 ;
        RECT 2369.990 441.360 2370.310 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2265.600 1152.300 2265.860 1152.560 ;
        RECT 2370.020 1152.300 2370.280 1152.560 ;
        RECT 2370.020 441.360 2370.280 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2265.590 1155.475 2265.870 1155.845 ;
        RECT 2265.660 1152.590 2265.800 1155.475 ;
        RECT 2265.600 1152.270 2265.860 1152.590 ;
        RECT 2370.020 1152.270 2370.280 1152.590 ;
        RECT 2370.080 441.650 2370.220 1152.270 ;
        RECT 2370.020 441.330 2370.280 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2265.590 1155.520 2265.870 1155.800 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2265.565 1155.810 2265.895 1155.825 ;
        RECT 2250.780 1155.800 2265.895 1155.810 ;
        RECT 2247.465 1155.510 2265.895 1155.800 ;
        RECT 2247.465 1155.200 2251.465 1155.510 ;
        RECT 2265.565 1155.495 2265.895 1155.510 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 2578.120 1014.230 2578.180 ;
        RECT 1219.990 2578.120 1220.310 2578.180 ;
        RECT 1013.910 2577.980 1220.310 2578.120 ;
        RECT 1013.910 2577.920 1014.230 2577.980 ;
        RECT 1219.990 2577.920 1220.310 2577.980 ;
      LAYER via ;
        RECT 1013.940 2577.920 1014.200 2578.180 ;
        RECT 1220.020 2577.920 1220.280 2578.180 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 2578.210 1014.140 3517.600 ;
        RECT 1013.940 2577.890 1014.200 2578.210 ;
        RECT 1220.020 2577.890 1220.280 2578.210 ;
        RECT 1220.080 2562.185 1220.220 2577.890 ;
        RECT 1219.910 2561.900 1220.220 2562.185 ;
        RECT 1219.910 2558.185 1220.190 2561.900 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 689.225 3429.325 689.395 3477.435 ;
        RECT 688.765 2898.585 688.935 2946.355 ;
        RECT 687.845 2849.625 688.015 2898.075 ;
        RECT 688.305 2753.065 688.475 2801.175 ;
        RECT 688.765 2608.225 688.935 2622.335 ;
      LAYER mcon ;
        RECT 689.225 3477.265 689.395 3477.435 ;
        RECT 688.765 2946.185 688.935 2946.355 ;
        RECT 687.845 2897.905 688.015 2898.075 ;
        RECT 688.305 2801.005 688.475 2801.175 ;
        RECT 688.765 2622.165 688.935 2622.335 ;
      LAYER met1 ;
        RECT 688.690 3491.360 689.010 3491.420 ;
        RECT 689.610 3491.360 689.930 3491.420 ;
        RECT 688.690 3491.220 689.930 3491.360 ;
        RECT 688.690 3491.160 689.010 3491.220 ;
        RECT 689.610 3491.160 689.930 3491.220 ;
        RECT 689.165 3477.420 689.455 3477.465 ;
        RECT 689.610 3477.420 689.930 3477.480 ;
        RECT 689.165 3477.280 689.930 3477.420 ;
        RECT 689.165 3477.235 689.455 3477.280 ;
        RECT 689.610 3477.220 689.930 3477.280 ;
        RECT 689.150 3429.480 689.470 3429.540 ;
        RECT 688.955 3429.340 689.470 3429.480 ;
        RECT 689.150 3429.280 689.470 3429.340 ;
        RECT 689.150 3395.140 689.470 3395.200 ;
        RECT 688.780 3395.000 689.470 3395.140 ;
        RECT 688.780 3394.860 688.920 3395.000 ;
        RECT 689.150 3394.940 689.470 3395.000 ;
        RECT 688.690 3394.600 689.010 3394.860 ;
        RECT 688.690 3367.600 689.010 3367.660 ;
        RECT 689.610 3367.600 689.930 3367.660 ;
        RECT 688.690 3367.460 689.930 3367.600 ;
        RECT 688.690 3367.400 689.010 3367.460 ;
        RECT 689.610 3367.400 689.930 3367.460 ;
        RECT 688.690 3270.700 689.010 3270.760 ;
        RECT 689.610 3270.700 689.930 3270.760 ;
        RECT 688.690 3270.560 689.930 3270.700 ;
        RECT 688.690 3270.500 689.010 3270.560 ;
        RECT 689.610 3270.500 689.930 3270.560 ;
        RECT 688.690 3174.140 689.010 3174.200 ;
        RECT 689.610 3174.140 689.930 3174.200 ;
        RECT 688.690 3174.000 689.930 3174.140 ;
        RECT 688.690 3173.940 689.010 3174.000 ;
        RECT 689.610 3173.940 689.930 3174.000 ;
        RECT 688.690 3077.580 689.010 3077.640 ;
        RECT 689.610 3077.580 689.930 3077.640 ;
        RECT 688.690 3077.440 689.930 3077.580 ;
        RECT 688.690 3077.380 689.010 3077.440 ;
        RECT 689.610 3077.380 689.930 3077.440 ;
        RECT 688.690 2981.020 689.010 2981.080 ;
        RECT 689.610 2981.020 689.930 2981.080 ;
        RECT 688.690 2980.880 689.930 2981.020 ;
        RECT 688.690 2980.820 689.010 2980.880 ;
        RECT 689.610 2980.820 689.930 2980.880 ;
        RECT 688.690 2946.340 689.010 2946.400 ;
        RECT 688.495 2946.200 689.010 2946.340 ;
        RECT 688.690 2946.140 689.010 2946.200 ;
        RECT 688.690 2898.740 689.010 2898.800 ;
        RECT 688.495 2898.600 689.010 2898.740 ;
        RECT 688.690 2898.540 689.010 2898.600 ;
        RECT 687.785 2898.060 688.075 2898.105 ;
        RECT 688.230 2898.060 688.550 2898.120 ;
        RECT 687.785 2897.920 688.550 2898.060 ;
        RECT 687.785 2897.875 688.075 2897.920 ;
        RECT 688.230 2897.860 688.550 2897.920 ;
        RECT 687.770 2849.780 688.090 2849.840 ;
        RECT 687.575 2849.640 688.090 2849.780 ;
        RECT 687.770 2849.580 688.090 2849.640 ;
        RECT 687.770 2815.240 688.090 2815.500 ;
        RECT 687.860 2814.760 688.000 2815.240 ;
        RECT 688.230 2814.760 688.550 2814.820 ;
        RECT 687.860 2814.620 688.550 2814.760 ;
        RECT 688.230 2814.560 688.550 2814.620 ;
        RECT 688.230 2801.160 688.550 2801.220 ;
        RECT 688.035 2801.020 688.550 2801.160 ;
        RECT 688.230 2800.960 688.550 2801.020 ;
        RECT 688.245 2753.220 688.535 2753.265 ;
        RECT 689.150 2753.220 689.470 2753.280 ;
        RECT 688.245 2753.080 689.470 2753.220 ;
        RECT 688.245 2753.035 688.535 2753.080 ;
        RECT 689.150 2753.020 689.470 2753.080 ;
        RECT 688.230 2718.200 688.550 2718.260 ;
        RECT 689.150 2718.200 689.470 2718.260 ;
        RECT 688.230 2718.060 689.470 2718.200 ;
        RECT 688.230 2718.000 688.550 2718.060 ;
        RECT 689.150 2718.000 689.470 2718.060 ;
        RECT 688.230 2670.260 688.550 2670.320 ;
        RECT 689.150 2670.260 689.470 2670.320 ;
        RECT 688.230 2670.120 689.470 2670.260 ;
        RECT 688.230 2670.060 688.550 2670.120 ;
        RECT 689.150 2670.060 689.470 2670.120 ;
        RECT 688.690 2622.320 689.010 2622.380 ;
        RECT 688.495 2622.180 689.010 2622.320 ;
        RECT 688.690 2622.120 689.010 2622.180 ;
        RECT 688.690 2608.380 689.010 2608.440 ;
        RECT 688.495 2608.240 689.010 2608.380 ;
        RECT 688.690 2608.180 689.010 2608.240 ;
        RECT 690.070 2577.100 690.390 2577.160 ;
        RECT 1042.890 2577.100 1043.210 2577.160 ;
        RECT 690.070 2576.960 1043.210 2577.100 ;
        RECT 690.070 2576.900 690.390 2576.960 ;
        RECT 1042.890 2576.900 1043.210 2576.960 ;
      LAYER via ;
        RECT 688.720 3491.160 688.980 3491.420 ;
        RECT 689.640 3491.160 689.900 3491.420 ;
        RECT 689.640 3477.220 689.900 3477.480 ;
        RECT 689.180 3429.280 689.440 3429.540 ;
        RECT 689.180 3394.940 689.440 3395.200 ;
        RECT 688.720 3394.600 688.980 3394.860 ;
        RECT 688.720 3367.400 688.980 3367.660 ;
        RECT 689.640 3367.400 689.900 3367.660 ;
        RECT 688.720 3270.500 688.980 3270.760 ;
        RECT 689.640 3270.500 689.900 3270.760 ;
        RECT 688.720 3173.940 688.980 3174.200 ;
        RECT 689.640 3173.940 689.900 3174.200 ;
        RECT 688.720 3077.380 688.980 3077.640 ;
        RECT 689.640 3077.380 689.900 3077.640 ;
        RECT 688.720 2980.820 688.980 2981.080 ;
        RECT 689.640 2980.820 689.900 2981.080 ;
        RECT 688.720 2946.140 688.980 2946.400 ;
        RECT 688.720 2898.540 688.980 2898.800 ;
        RECT 688.260 2897.860 688.520 2898.120 ;
        RECT 687.800 2849.580 688.060 2849.840 ;
        RECT 687.800 2815.240 688.060 2815.500 ;
        RECT 688.260 2814.560 688.520 2814.820 ;
        RECT 688.260 2800.960 688.520 2801.220 ;
        RECT 689.180 2753.020 689.440 2753.280 ;
        RECT 688.260 2718.000 688.520 2718.260 ;
        RECT 689.180 2718.000 689.440 2718.260 ;
        RECT 688.260 2670.060 688.520 2670.320 ;
        RECT 689.180 2670.060 689.440 2670.320 ;
        RECT 688.720 2622.120 688.980 2622.380 ;
        RECT 688.720 2608.180 688.980 2608.440 ;
        RECT 690.100 2576.900 690.360 2577.160 ;
        RECT 1042.920 2576.900 1043.180 2577.160 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.780 3517.230 689.380 3517.370 ;
        RECT 688.780 3491.450 688.920 3517.230 ;
        RECT 688.720 3491.130 688.980 3491.450 ;
        RECT 689.640 3491.130 689.900 3491.450 ;
        RECT 689.700 3477.510 689.840 3491.130 ;
        RECT 689.640 3477.190 689.900 3477.510 ;
        RECT 689.180 3429.250 689.440 3429.570 ;
        RECT 689.240 3395.230 689.380 3429.250 ;
        RECT 689.180 3394.910 689.440 3395.230 ;
        RECT 688.720 3394.570 688.980 3394.890 ;
        RECT 688.780 3367.690 688.920 3394.570 ;
        RECT 688.720 3367.370 688.980 3367.690 ;
        RECT 689.640 3367.370 689.900 3367.690 ;
        RECT 689.700 3318.810 689.840 3367.370 ;
        RECT 688.780 3318.670 689.840 3318.810 ;
        RECT 688.780 3270.790 688.920 3318.670 ;
        RECT 688.720 3270.470 688.980 3270.790 ;
        RECT 689.640 3270.470 689.900 3270.790 ;
        RECT 689.700 3222.250 689.840 3270.470 ;
        RECT 688.780 3222.110 689.840 3222.250 ;
        RECT 688.780 3174.230 688.920 3222.110 ;
        RECT 688.720 3173.910 688.980 3174.230 ;
        RECT 689.640 3173.910 689.900 3174.230 ;
        RECT 689.700 3125.690 689.840 3173.910 ;
        RECT 688.780 3125.550 689.840 3125.690 ;
        RECT 688.780 3077.670 688.920 3125.550 ;
        RECT 688.720 3077.350 688.980 3077.670 ;
        RECT 689.640 3077.350 689.900 3077.670 ;
        RECT 689.700 3029.130 689.840 3077.350 ;
        RECT 688.780 3028.990 689.840 3029.130 ;
        RECT 688.780 2981.110 688.920 3028.990 ;
        RECT 688.720 2980.790 688.980 2981.110 ;
        RECT 689.640 2980.850 689.900 2981.110 ;
        RECT 689.240 2980.790 689.900 2980.850 ;
        RECT 689.240 2980.710 689.840 2980.790 ;
        RECT 689.240 2959.770 689.380 2980.710 ;
        RECT 688.780 2959.630 689.380 2959.770 ;
        RECT 688.780 2946.430 688.920 2959.630 ;
        RECT 688.720 2946.110 688.980 2946.430 ;
        RECT 688.720 2898.570 688.980 2898.830 ;
        RECT 688.320 2898.510 688.980 2898.570 ;
        RECT 688.320 2898.430 688.920 2898.510 ;
        RECT 688.320 2898.150 688.460 2898.430 ;
        RECT 688.260 2897.830 688.520 2898.150 ;
        RECT 687.800 2849.550 688.060 2849.870 ;
        RECT 687.860 2815.530 688.000 2849.550 ;
        RECT 687.800 2815.210 688.060 2815.530 ;
        RECT 688.260 2814.530 688.520 2814.850 ;
        RECT 688.320 2801.250 688.460 2814.530 ;
        RECT 688.260 2800.930 688.520 2801.250 ;
        RECT 689.180 2752.990 689.440 2753.310 ;
        RECT 689.240 2718.290 689.380 2752.990 ;
        RECT 688.260 2717.970 688.520 2718.290 ;
        RECT 689.180 2717.970 689.440 2718.290 ;
        RECT 688.320 2670.350 688.460 2717.970 ;
        RECT 688.260 2670.030 688.520 2670.350 ;
        RECT 689.180 2670.030 689.440 2670.350 ;
        RECT 689.240 2656.490 689.380 2670.030 ;
        RECT 688.780 2656.350 689.380 2656.490 ;
        RECT 688.780 2622.410 688.920 2656.350 ;
        RECT 688.720 2622.090 688.980 2622.410 ;
        RECT 688.720 2608.150 688.980 2608.470 ;
        RECT 688.780 2594.610 688.920 2608.150 ;
        RECT 688.780 2594.470 689.840 2594.610 ;
        RECT 689.700 2577.610 689.840 2594.470 ;
        RECT 689.700 2577.470 690.300 2577.610 ;
        RECT 690.160 2577.190 690.300 2577.470 ;
        RECT 690.100 2576.870 690.360 2577.190 ;
        RECT 1042.920 2576.870 1043.180 2577.190 ;
        RECT 1042.980 2562.185 1043.120 2576.870 ;
        RECT 1042.810 2561.900 1043.120 2562.185 ;
        RECT 1042.810 2558.185 1043.090 2561.900 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
        RECT 364.925 3236.205 365.095 3284.315 ;
        RECT 365.385 3084.225 365.555 3132.675 ;
        RECT 364.465 2946.525 364.635 2994.635 ;
        RECT 363.085 2849.625 363.255 2898.075 ;
        RECT 363.545 2753.065 363.715 2801.175 ;
        RECT 364.005 2608.225 364.175 2622.335 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
        RECT 364.925 3284.145 365.095 3284.315 ;
        RECT 365.385 3132.505 365.555 3132.675 ;
        RECT 364.465 2994.465 364.635 2994.635 ;
        RECT 363.085 2897.905 363.255 2898.075 ;
        RECT 363.545 2801.005 363.715 2801.175 ;
        RECT 364.005 2622.165 364.175 2622.335 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 364.390 3298.240 364.710 3298.300 ;
        RECT 365.310 3298.240 365.630 3298.300 ;
        RECT 364.390 3298.100 365.630 3298.240 ;
        RECT 364.390 3298.040 364.710 3298.100 ;
        RECT 365.310 3298.040 365.630 3298.100 ;
        RECT 364.865 3284.300 365.155 3284.345 ;
        RECT 365.310 3284.300 365.630 3284.360 ;
        RECT 364.865 3284.160 365.630 3284.300 ;
        RECT 364.865 3284.115 365.155 3284.160 ;
        RECT 365.310 3284.100 365.630 3284.160 ;
        RECT 364.850 3236.360 365.170 3236.420 ;
        RECT 364.655 3236.220 365.170 3236.360 ;
        RECT 364.850 3236.160 365.170 3236.220 ;
        RECT 364.850 3202.020 365.170 3202.080 ;
        RECT 364.020 3201.880 365.170 3202.020 ;
        RECT 364.020 3201.400 364.160 3201.880 ;
        RECT 364.850 3201.820 365.170 3201.880 ;
        RECT 363.930 3201.140 364.250 3201.400 ;
        RECT 363.930 3187.740 364.250 3187.800 ;
        RECT 364.390 3187.740 364.710 3187.800 ;
        RECT 363.930 3187.600 364.710 3187.740 ;
        RECT 363.930 3187.540 364.250 3187.600 ;
        RECT 364.390 3187.540 364.710 3187.600 ;
        RECT 365.310 3132.660 365.630 3132.720 ;
        RECT 365.115 3132.520 365.630 3132.660 ;
        RECT 365.310 3132.460 365.630 3132.520 ;
        RECT 365.310 3084.380 365.630 3084.440 ;
        RECT 365.115 3084.240 365.630 3084.380 ;
        RECT 365.310 3084.180 365.630 3084.240 ;
        RECT 365.310 3057.180 365.630 3057.240 ;
        RECT 364.480 3057.040 365.630 3057.180 ;
        RECT 364.480 3056.560 364.620 3057.040 ;
        RECT 365.310 3056.980 365.630 3057.040 ;
        RECT 364.390 3056.300 364.710 3056.560 ;
        RECT 364.850 3007.880 365.170 3007.940 ;
        RECT 365.770 3007.880 366.090 3007.940 ;
        RECT 364.850 3007.740 366.090 3007.880 ;
        RECT 364.850 3007.680 365.170 3007.740 ;
        RECT 365.770 3007.680 366.090 3007.740 ;
        RECT 364.405 2994.620 364.695 2994.665 ;
        RECT 364.850 2994.620 365.170 2994.680 ;
        RECT 364.405 2994.480 365.170 2994.620 ;
        RECT 364.405 2994.435 364.695 2994.480 ;
        RECT 364.850 2994.420 365.170 2994.480 ;
        RECT 364.390 2946.680 364.710 2946.740 ;
        RECT 364.195 2946.540 364.710 2946.680 ;
        RECT 364.390 2946.480 364.710 2946.540 ;
        RECT 363.470 2912.000 363.790 2912.060 ;
        RECT 364.390 2912.000 364.710 2912.060 ;
        RECT 363.470 2911.860 364.710 2912.000 ;
        RECT 363.470 2911.800 363.790 2911.860 ;
        RECT 364.390 2911.800 364.710 2911.860 ;
        RECT 363.025 2898.060 363.315 2898.105 ;
        RECT 363.470 2898.060 363.790 2898.120 ;
        RECT 363.025 2897.920 363.790 2898.060 ;
        RECT 363.025 2897.875 363.315 2897.920 ;
        RECT 363.470 2897.860 363.790 2897.920 ;
        RECT 363.010 2849.780 363.330 2849.840 ;
        RECT 362.815 2849.640 363.330 2849.780 ;
        RECT 363.010 2849.580 363.330 2849.640 ;
        RECT 363.010 2815.240 363.330 2815.500 ;
        RECT 363.100 2814.760 363.240 2815.240 ;
        RECT 363.470 2814.760 363.790 2814.820 ;
        RECT 363.100 2814.620 363.790 2814.760 ;
        RECT 363.470 2814.560 363.790 2814.620 ;
        RECT 363.470 2801.160 363.790 2801.220 ;
        RECT 363.275 2801.020 363.790 2801.160 ;
        RECT 363.470 2800.960 363.790 2801.020 ;
        RECT 363.485 2753.220 363.775 2753.265 ;
        RECT 364.390 2753.220 364.710 2753.280 ;
        RECT 363.485 2753.080 364.710 2753.220 ;
        RECT 363.485 2753.035 363.775 2753.080 ;
        RECT 364.390 2753.020 364.710 2753.080 ;
        RECT 363.470 2718.200 363.790 2718.260 ;
        RECT 364.390 2718.200 364.710 2718.260 ;
        RECT 363.470 2718.060 364.710 2718.200 ;
        RECT 363.470 2718.000 363.790 2718.060 ;
        RECT 364.390 2718.000 364.710 2718.060 ;
        RECT 363.470 2670.260 363.790 2670.320 ;
        RECT 364.390 2670.260 364.710 2670.320 ;
        RECT 363.470 2670.120 364.710 2670.260 ;
        RECT 363.470 2670.060 363.790 2670.120 ;
        RECT 364.390 2670.060 364.710 2670.120 ;
        RECT 363.930 2622.320 364.250 2622.380 ;
        RECT 363.735 2622.180 364.250 2622.320 ;
        RECT 363.930 2622.120 364.250 2622.180 ;
        RECT 363.930 2608.380 364.250 2608.440 ;
        RECT 363.735 2608.240 364.250 2608.380 ;
        RECT 363.930 2608.180 364.250 2608.240 ;
        RECT 363.930 2578.120 364.250 2578.180 ;
        RECT 866.250 2578.120 866.570 2578.180 ;
        RECT 363.930 2577.980 866.570 2578.120 ;
        RECT 363.930 2577.920 364.250 2577.980 ;
        RECT 866.250 2577.920 866.570 2577.980 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 364.420 3298.040 364.680 3298.300 ;
        RECT 365.340 3298.040 365.600 3298.300 ;
        RECT 365.340 3284.100 365.600 3284.360 ;
        RECT 364.880 3236.160 365.140 3236.420 ;
        RECT 364.880 3201.820 365.140 3202.080 ;
        RECT 363.960 3201.140 364.220 3201.400 ;
        RECT 363.960 3187.540 364.220 3187.800 ;
        RECT 364.420 3187.540 364.680 3187.800 ;
        RECT 365.340 3132.460 365.600 3132.720 ;
        RECT 365.340 3084.180 365.600 3084.440 ;
        RECT 365.340 3056.980 365.600 3057.240 ;
        RECT 364.420 3056.300 364.680 3056.560 ;
        RECT 364.880 3007.680 365.140 3007.940 ;
        RECT 365.800 3007.680 366.060 3007.940 ;
        RECT 364.880 2994.420 365.140 2994.680 ;
        RECT 364.420 2946.480 364.680 2946.740 ;
        RECT 363.500 2911.800 363.760 2912.060 ;
        RECT 364.420 2911.800 364.680 2912.060 ;
        RECT 363.500 2897.860 363.760 2898.120 ;
        RECT 363.040 2849.580 363.300 2849.840 ;
        RECT 363.040 2815.240 363.300 2815.500 ;
        RECT 363.500 2814.560 363.760 2814.820 ;
        RECT 363.500 2800.960 363.760 2801.220 ;
        RECT 364.420 2753.020 364.680 2753.280 ;
        RECT 363.500 2718.000 363.760 2718.260 ;
        RECT 364.420 2718.000 364.680 2718.260 ;
        RECT 363.500 2670.060 363.760 2670.320 ;
        RECT 364.420 2670.060 364.680 2670.320 ;
        RECT 363.960 2622.120 364.220 2622.380 ;
        RECT 363.960 2608.180 364.220 2608.440 ;
        RECT 363.960 2577.920 364.220 2578.180 ;
        RECT 866.280 2577.920 866.540 2578.180 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.330 364.620 3298.410 ;
        RECT 364.020 3298.270 364.680 3298.330 ;
        RECT 364.420 3298.010 364.680 3298.270 ;
        RECT 365.340 3298.010 365.600 3298.330 ;
        RECT 365.400 3284.390 365.540 3298.010 ;
        RECT 365.340 3284.070 365.600 3284.390 ;
        RECT 364.880 3236.130 365.140 3236.450 ;
        RECT 364.940 3202.110 365.080 3236.130 ;
        RECT 364.880 3201.790 365.140 3202.110 ;
        RECT 363.960 3201.110 364.220 3201.430 ;
        RECT 364.020 3187.830 364.160 3201.110 ;
        RECT 363.960 3187.510 364.220 3187.830 ;
        RECT 364.420 3187.510 364.680 3187.830 ;
        RECT 364.480 3152.890 364.620 3187.510 ;
        RECT 364.480 3152.750 365.540 3152.890 ;
        RECT 365.400 3132.750 365.540 3152.750 ;
        RECT 365.340 3132.430 365.600 3132.750 ;
        RECT 365.340 3084.150 365.600 3084.470 ;
        RECT 365.400 3057.270 365.540 3084.150 ;
        RECT 365.340 3056.950 365.600 3057.270 ;
        RECT 364.420 3056.270 364.680 3056.590 ;
        RECT 364.480 3042.730 364.620 3056.270 ;
        RECT 364.870 3042.730 365.150 3042.845 ;
        RECT 364.480 3042.590 365.150 3042.730 ;
        RECT 364.870 3042.475 365.150 3042.590 ;
        RECT 365.790 3042.475 366.070 3042.845 ;
        RECT 365.860 3007.970 366.000 3042.475 ;
        RECT 364.880 3007.650 365.140 3007.970 ;
        RECT 365.800 3007.650 366.060 3007.970 ;
        RECT 364.940 2994.710 365.080 3007.650 ;
        RECT 364.880 2994.390 365.140 2994.710 ;
        RECT 364.420 2946.450 364.680 2946.770 ;
        RECT 364.480 2912.090 364.620 2946.450 ;
        RECT 363.500 2911.770 363.760 2912.090 ;
        RECT 364.420 2911.770 364.680 2912.090 ;
        RECT 363.560 2898.150 363.700 2911.770 ;
        RECT 363.500 2897.830 363.760 2898.150 ;
        RECT 363.040 2849.550 363.300 2849.870 ;
        RECT 363.100 2815.530 363.240 2849.550 ;
        RECT 363.040 2815.210 363.300 2815.530 ;
        RECT 363.500 2814.530 363.760 2814.850 ;
        RECT 363.560 2801.250 363.700 2814.530 ;
        RECT 363.500 2800.930 363.760 2801.250 ;
        RECT 364.420 2752.990 364.680 2753.310 ;
        RECT 364.480 2718.290 364.620 2752.990 ;
        RECT 363.500 2717.970 363.760 2718.290 ;
        RECT 364.420 2717.970 364.680 2718.290 ;
        RECT 363.560 2670.350 363.700 2717.970 ;
        RECT 363.500 2670.030 363.760 2670.350 ;
        RECT 364.420 2670.030 364.680 2670.350 ;
        RECT 364.480 2656.490 364.620 2670.030 ;
        RECT 364.020 2656.350 364.620 2656.490 ;
        RECT 364.020 2622.410 364.160 2656.350 ;
        RECT 363.960 2622.090 364.220 2622.410 ;
        RECT 363.960 2608.150 364.220 2608.470 ;
        RECT 364.020 2578.210 364.160 2608.150 ;
        RECT 363.960 2577.890 364.220 2578.210 ;
        RECT 866.280 2577.890 866.540 2578.210 ;
        RECT 866.340 2562.185 866.480 2577.890 ;
        RECT 866.170 2561.900 866.480 2562.185 ;
        RECT 866.170 2558.185 866.450 2561.900 ;
      LAYER via2 ;
        RECT 364.870 3042.520 365.150 3042.800 ;
        RECT 365.790 3042.520 366.070 3042.800 ;
      LAYER met3 ;
        RECT 364.845 3042.810 365.175 3042.825 ;
        RECT 365.765 3042.810 366.095 3042.825 ;
        RECT 364.845 3042.510 366.095 3042.810 ;
        RECT 364.845 3042.495 365.175 3042.510 ;
        RECT 365.765 3042.495 366.095 3042.510 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
        RECT 40.165 2898.585 40.335 2946.355 ;
        RECT 40.165 2718.725 40.335 2752.895 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
        RECT 40.165 2946.185 40.335 2946.355 ;
        RECT 40.165 2752.725 40.335 2752.895 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 40.090 2946.340 40.410 2946.400 ;
        RECT 39.895 2946.200 40.410 2946.340 ;
        RECT 40.090 2946.140 40.410 2946.200 ;
        RECT 40.090 2898.740 40.410 2898.800 ;
        RECT 39.895 2898.600 40.410 2898.740 ;
        RECT 40.090 2898.540 40.410 2898.600 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 40.550 2898.060 40.870 2898.120 ;
        RECT 39.630 2897.920 40.870 2898.060 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 40.550 2897.860 40.870 2897.920 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 40.550 2814.760 40.870 2814.820 ;
        RECT 39.630 2814.620 40.870 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.550 2814.560 40.870 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 39.895 2752.740 40.410 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.105 2718.880 40.395 2718.925 ;
        RECT 41.010 2718.880 41.330 2718.940 ;
        RECT 40.105 2718.740 41.330 2718.880 ;
        RECT 40.105 2718.695 40.395 2718.740 ;
        RECT 41.010 2718.680 41.330 2718.740 ;
        RECT 40.550 2621.640 40.870 2621.700 ;
        RECT 41.470 2621.640 41.790 2621.700 ;
        RECT 40.550 2621.500 41.790 2621.640 ;
        RECT 40.550 2621.440 40.870 2621.500 ;
        RECT 41.470 2621.440 41.790 2621.500 ;
        RECT 40.550 2577.100 40.870 2577.160 ;
        RECT 689.610 2577.100 689.930 2577.160 ;
        RECT 40.550 2576.960 689.930 2577.100 ;
        RECT 40.550 2576.900 40.870 2576.960 ;
        RECT 689.610 2576.900 689.930 2576.960 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 40.120 2946.140 40.380 2946.400 ;
        RECT 40.120 2898.540 40.380 2898.800 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 40.580 2897.860 40.840 2898.120 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.580 2814.560 40.840 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 41.040 2718.680 41.300 2718.940 ;
        RECT 40.580 2621.440 40.840 2621.700 ;
        RECT 41.500 2621.440 41.760 2621.700 ;
        RECT 40.580 2576.900 40.840 2577.160 ;
        RECT 689.640 2576.900 689.900 2577.160 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2946.430 40.320 2959.630 ;
        RECT 40.120 2946.110 40.380 2946.430 ;
        RECT 40.120 2898.570 40.380 2898.830 ;
        RECT 39.720 2898.510 40.380 2898.570 ;
        RECT 39.720 2898.430 40.320 2898.510 ;
        RECT 39.720 2898.150 39.860 2898.430 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 40.580 2897.830 40.840 2898.150 ;
        RECT 40.640 2814.850 40.780 2897.830 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 40.580 2814.530 40.840 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 41.040 2718.650 41.300 2718.970 ;
        RECT 41.100 2704.885 41.240 2718.650 ;
        RECT 41.030 2704.515 41.310 2704.885 ;
        RECT 41.950 2704.515 42.230 2704.885 ;
        RECT 42.020 2669.410 42.160 2704.515 ;
        RECT 40.640 2669.270 42.160 2669.410 ;
        RECT 40.640 2656.605 40.780 2669.270 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.490 2656.235 41.770 2656.605 ;
        RECT 41.560 2621.730 41.700 2656.235 ;
        RECT 40.580 2621.410 40.840 2621.730 ;
        RECT 41.500 2621.410 41.760 2621.730 ;
        RECT 40.640 2577.190 40.780 2621.410 ;
        RECT 40.580 2576.870 40.840 2577.190 ;
        RECT 689.640 2576.870 689.900 2577.190 ;
        RECT 689.700 2562.185 689.840 2576.870 ;
        RECT 689.530 2561.900 689.840 2562.185 ;
        RECT 689.530 2558.185 689.810 2561.900 ;
      LAYER via2 ;
        RECT 41.030 2704.560 41.310 2704.840 ;
        RECT 41.950 2704.560 42.230 2704.840 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.490 2656.280 41.770 2656.560 ;
      LAYER met3 ;
        RECT 41.005 2704.850 41.335 2704.865 ;
        RECT 41.925 2704.850 42.255 2704.865 ;
        RECT 41.005 2704.550 42.255 2704.850 ;
        RECT 41.005 2704.535 41.335 2704.550 ;
        RECT 41.925 2704.535 42.255 2704.550 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.465 2656.570 41.795 2656.585 ;
        RECT 40.545 2656.270 41.795 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.465 2656.255 41.795 2656.270 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 45.150 3263.900 45.470 3263.960 ;
        RECT 15.250 3263.760 45.470 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 45.150 3263.700 45.470 3263.760 ;
        RECT 45.150 3122.120 45.470 3122.180 ;
        RECT 644.990 3122.120 645.310 3122.180 ;
        RECT 45.150 3121.980 645.310 3122.120 ;
        RECT 45.150 3121.920 45.470 3121.980 ;
        RECT 644.990 3121.920 645.310 3121.980 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 45.180 3263.700 45.440 3263.960 ;
        RECT 45.180 3121.920 45.440 3122.180 ;
        RECT 645.020 3121.920 645.280 3122.180 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 45.180 3263.670 45.440 3263.990 ;
        RECT 45.240 3122.210 45.380 3263.670 ;
        RECT 45.180 3121.890 45.440 3122.210 ;
        RECT 645.020 3121.890 645.280 3122.210 ;
        RECT 645.080 2466.885 645.220 3121.890 ;
        RECT 645.010 2466.515 645.290 2466.885 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 645.010 2466.560 645.290 2466.840 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 644.985 2466.850 645.315 2466.865 ;
        RECT 644.985 2466.840 660.100 2466.850 ;
        RECT 644.985 2466.550 664.000 2466.840 ;
        RECT 644.985 2466.535 645.315 2466.550 ;
        RECT 660.000 2466.240 664.000 2466.550 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 58.490 2974.220 58.810 2974.280 ;
        RECT 16.630 2974.080 58.810 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 58.490 2974.020 58.810 2974.080 ;
        RECT 58.490 2352.700 58.810 2352.760 ;
        RECT 641.770 2352.700 642.090 2352.760 ;
        RECT 58.490 2352.560 642.090 2352.700 ;
        RECT 58.490 2352.500 58.810 2352.560 ;
        RECT 641.770 2352.500 642.090 2352.560 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 58.520 2974.020 58.780 2974.280 ;
        RECT 58.520 2352.500 58.780 2352.760 ;
        RECT 641.800 2352.500 642.060 2352.760 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 58.520 2973.990 58.780 2974.310 ;
        RECT 58.580 2352.790 58.720 2973.990 ;
        RECT 58.520 2352.470 58.780 2352.790 ;
        RECT 641.800 2352.645 642.060 2352.790 ;
        RECT 641.790 2352.275 642.070 2352.645 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
        RECT 641.790 2352.320 642.070 2352.600 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
        RECT 641.765 2352.610 642.095 2352.625 ;
        RECT 641.765 2352.600 660.100 2352.610 ;
        RECT 641.765 2352.310 664.000 2352.600 ;
        RECT 641.765 2352.295 642.095 2352.310 ;
        RECT 660.000 2352.000 664.000 2352.310 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2242.540 18.790 2242.600 ;
        RECT 641.770 2242.540 642.090 2242.600 ;
        RECT 18.470 2242.400 642.090 2242.540 ;
        RECT 18.470 2242.340 18.790 2242.400 ;
        RECT 641.770 2242.340 642.090 2242.400 ;
      LAYER via ;
        RECT 18.500 2242.340 18.760 2242.600 ;
        RECT 641.800 2242.340 642.060 2242.600 ;
      LAYER met2 ;
        RECT 18.490 2692.955 18.770 2693.325 ;
        RECT 18.560 2242.630 18.700 2692.955 ;
        RECT 18.500 2242.310 18.760 2242.630 ;
        RECT 641.800 2242.310 642.060 2242.630 ;
        RECT 641.860 2238.405 642.000 2242.310 ;
        RECT 641.790 2238.035 642.070 2238.405 ;
      LAYER via2 ;
        RECT 18.490 2693.000 18.770 2693.280 ;
        RECT 641.790 2238.080 642.070 2238.360 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 18.465 2693.290 18.795 2693.305 ;
        RECT -4.800 2692.990 18.795 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 18.465 2692.975 18.795 2692.990 ;
        RECT 641.765 2238.370 642.095 2238.385 ;
        RECT 641.765 2238.360 660.100 2238.370 ;
        RECT 641.765 2238.070 664.000 2238.360 ;
        RECT 641.765 2238.055 642.095 2238.070 ;
        RECT 660.000 2237.760 664.000 2238.070 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2125.240 19.250 2125.300 ;
        RECT 641.770 2125.240 642.090 2125.300 ;
        RECT 18.930 2125.100 642.090 2125.240 ;
        RECT 18.930 2125.040 19.250 2125.100 ;
        RECT 641.770 2125.040 642.090 2125.100 ;
      LAYER via ;
        RECT 18.960 2125.040 19.220 2125.300 ;
        RECT 641.800 2125.040 642.060 2125.300 ;
      LAYER met2 ;
        RECT 18.950 2405.315 19.230 2405.685 ;
        RECT 19.020 2125.330 19.160 2405.315 ;
        RECT 18.960 2125.010 19.220 2125.330 ;
        RECT 641.800 2125.010 642.060 2125.330 ;
        RECT 641.860 2123.485 642.000 2125.010 ;
        RECT 641.790 2123.115 642.070 2123.485 ;
      LAYER via2 ;
        RECT 18.950 2405.360 19.230 2405.640 ;
        RECT 641.790 2123.160 642.070 2123.440 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 18.925 2405.650 19.255 2405.665 ;
        RECT -4.800 2405.350 19.255 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 18.925 2405.335 19.255 2405.350 ;
        RECT 641.765 2123.450 642.095 2123.465 ;
        RECT 641.765 2123.440 660.100 2123.450 ;
        RECT 641.765 2123.150 664.000 2123.440 ;
        RECT 641.765 2123.135 642.095 2123.150 ;
        RECT 660.000 2122.840 664.000 2123.150 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2014.740 17.410 2014.800 ;
        RECT 641.770 2014.740 642.090 2014.800 ;
        RECT 17.090 2014.600 642.090 2014.740 ;
        RECT 17.090 2014.540 17.410 2014.600 ;
        RECT 641.770 2014.540 642.090 2014.600 ;
      LAYER via ;
        RECT 17.120 2014.540 17.380 2014.800 ;
        RECT 641.800 2014.540 642.060 2014.800 ;
      LAYER met2 ;
        RECT 17.110 2118.355 17.390 2118.725 ;
        RECT 17.180 2014.830 17.320 2118.355 ;
        RECT 17.120 2014.510 17.380 2014.830 ;
        RECT 641.800 2014.510 642.060 2014.830 ;
        RECT 641.860 2009.245 642.000 2014.510 ;
        RECT 641.790 2008.875 642.070 2009.245 ;
      LAYER via2 ;
        RECT 17.110 2118.400 17.390 2118.680 ;
        RECT 641.790 2008.920 642.070 2009.200 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 17.085 2118.690 17.415 2118.705 ;
        RECT -4.800 2118.390 17.415 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 17.085 2118.375 17.415 2118.390 ;
        RECT 641.765 2009.210 642.095 2009.225 ;
        RECT 641.765 2009.200 660.100 2009.210 ;
        RECT 641.765 2008.910 664.000 2009.200 ;
        RECT 641.765 2008.895 642.095 2008.910 ;
        RECT 660.000 2008.600 664.000 2008.910 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 644.990 1835.220 645.310 1835.280 ;
        RECT 15.710 1835.080 645.310 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 644.990 1835.020 645.310 1835.080 ;
      LAYER via ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 645.020 1835.020 645.280 1835.280 ;
      LAYER met2 ;
        RECT 645.010 1894.635 645.290 1895.005 ;
        RECT 645.080 1835.310 645.220 1894.635 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 645.020 1834.990 645.280 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 645.010 1894.680 645.290 1894.960 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 644.985 1894.970 645.315 1894.985 ;
        RECT 644.985 1894.960 660.100 1894.970 ;
        RECT 644.985 1894.670 664.000 1894.960 ;
        RECT 644.985 1894.655 645.315 1894.670 ;
        RECT 660.000 1894.360 664.000 1894.670 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2265.110 1256.200 2265.430 1256.260 ;
        RECT 2287.190 1256.200 2287.510 1256.260 ;
        RECT 2265.110 1256.060 2287.510 1256.200 ;
        RECT 2265.110 1256.000 2265.430 1256.060 ;
        RECT 2287.190 1256.000 2287.510 1256.060 ;
        RECT 2287.190 676.160 2287.510 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2287.190 676.020 2901.150 676.160 ;
        RECT 2287.190 675.960 2287.510 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2265.140 1256.000 2265.400 1256.260 ;
        RECT 2287.220 1256.000 2287.480 1256.260 ;
        RECT 2287.220 675.960 2287.480 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2265.130 1262.235 2265.410 1262.605 ;
        RECT 2265.200 1256.290 2265.340 1262.235 ;
        RECT 2265.140 1255.970 2265.400 1256.290 ;
        RECT 2287.220 1255.970 2287.480 1256.290 ;
        RECT 2287.280 676.250 2287.420 1255.970 ;
        RECT 2287.220 675.930 2287.480 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2265.130 1262.280 2265.410 1262.560 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2265.105 1262.570 2265.435 1262.585 ;
        RECT 2250.780 1262.560 2265.435 1262.570 ;
        RECT 2247.465 1262.270 2265.435 1262.560 ;
        RECT 2247.465 1261.960 2251.465 1262.270 ;
        RECT 2265.105 1262.255 2265.435 1262.270 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 645.910 1545.540 646.230 1545.600 ;
        RECT 16.630 1545.400 646.230 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 645.910 1545.340 646.230 1545.400 ;
      LAYER via ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 645.940 1545.340 646.200 1545.600 ;
      LAYER met2 ;
        RECT 645.930 1780.395 646.210 1780.765 ;
        RECT 646.000 1545.630 646.140 1780.395 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 645.940 1545.310 646.200 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 645.930 1780.440 646.210 1780.720 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 645.905 1780.730 646.235 1780.745 ;
        RECT 645.905 1780.720 660.100 1780.730 ;
        RECT 645.905 1780.430 664.000 1780.720 ;
        RECT 645.905 1780.415 646.235 1780.430 ;
        RECT 660.000 1780.120 664.000 1780.430 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 44.690 1663.180 45.010 1663.240 ;
        RECT 641.770 1663.180 642.090 1663.240 ;
        RECT 44.690 1663.040 642.090 1663.180 ;
        RECT 44.690 1662.980 45.010 1663.040 ;
        RECT 641.770 1662.980 642.090 1663.040 ;
        RECT 17.550 1330.320 17.870 1330.380 ;
        RECT 44.690 1330.320 45.010 1330.380 ;
        RECT 17.550 1330.180 45.010 1330.320 ;
        RECT 17.550 1330.120 17.870 1330.180 ;
        RECT 44.690 1330.120 45.010 1330.180 ;
      LAYER via ;
        RECT 44.720 1662.980 44.980 1663.240 ;
        RECT 641.800 1662.980 642.060 1663.240 ;
        RECT 17.580 1330.120 17.840 1330.380 ;
        RECT 44.720 1330.120 44.980 1330.380 ;
      LAYER met2 ;
        RECT 641.790 1665.475 642.070 1665.845 ;
        RECT 641.860 1663.270 642.000 1665.475 ;
        RECT 44.720 1662.950 44.980 1663.270 ;
        RECT 641.800 1662.950 642.060 1663.270 ;
        RECT 44.780 1330.410 44.920 1662.950 ;
        RECT 17.580 1330.090 17.840 1330.410 ;
        RECT 44.720 1330.090 44.980 1330.410 ;
        RECT 17.640 1328.565 17.780 1330.090 ;
        RECT 17.570 1328.195 17.850 1328.565 ;
      LAYER via2 ;
        RECT 641.790 1665.520 642.070 1665.800 ;
        RECT 17.570 1328.240 17.850 1328.520 ;
      LAYER met3 ;
        RECT 641.765 1665.810 642.095 1665.825 ;
        RECT 641.765 1665.800 660.100 1665.810 ;
        RECT 641.765 1665.510 664.000 1665.800 ;
        RECT 641.765 1665.495 642.095 1665.510 ;
        RECT 660.000 1665.200 664.000 1665.510 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 17.545 1328.530 17.875 1328.545 ;
        RECT -4.800 1328.230 17.875 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 17.545 1328.215 17.875 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 58.490 1545.880 58.810 1545.940 ;
        RECT 641.770 1545.880 642.090 1545.940 ;
        RECT 58.490 1545.740 642.090 1545.880 ;
        RECT 58.490 1545.680 58.810 1545.740 ;
        RECT 641.770 1545.680 642.090 1545.740 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 58.490 1117.820 58.810 1117.880 ;
        RECT 15.710 1117.680 58.810 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 58.490 1117.620 58.810 1117.680 ;
      LAYER via ;
        RECT 58.520 1545.680 58.780 1545.940 ;
        RECT 641.800 1545.680 642.060 1545.940 ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 58.520 1117.620 58.780 1117.880 ;
      LAYER met2 ;
        RECT 641.790 1551.235 642.070 1551.605 ;
        RECT 641.860 1545.970 642.000 1551.235 ;
        RECT 58.520 1545.650 58.780 1545.970 ;
        RECT 641.800 1545.650 642.060 1545.970 ;
        RECT 58.580 1117.910 58.720 1545.650 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 58.520 1117.590 58.780 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 641.790 1551.280 642.070 1551.560 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 641.765 1551.570 642.095 1551.585 ;
        RECT 641.765 1551.560 660.100 1551.570 ;
        RECT 641.765 1551.270 664.000 1551.560 ;
        RECT 641.765 1551.255 642.095 1551.270 ;
        RECT 660.000 1550.960 664.000 1551.270 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 1435.380 65.710 1435.440 ;
        RECT 641.770 1435.380 642.090 1435.440 ;
        RECT 65.390 1435.240 642.090 1435.380 ;
        RECT 65.390 1435.180 65.710 1435.240 ;
        RECT 641.770 1435.180 642.090 1435.240 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 65.390 903.960 65.710 904.020 ;
        RECT 16.170 903.820 65.710 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 65.390 903.760 65.710 903.820 ;
      LAYER via ;
        RECT 65.420 1435.180 65.680 1435.440 ;
        RECT 641.800 1435.180 642.060 1435.440 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 65.420 903.760 65.680 904.020 ;
      LAYER met2 ;
        RECT 641.790 1436.995 642.070 1437.365 ;
        RECT 641.860 1435.470 642.000 1436.995 ;
        RECT 65.420 1435.150 65.680 1435.470 ;
        RECT 641.800 1435.150 642.060 1435.470 ;
        RECT 65.480 904.050 65.620 1435.150 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 65.420 903.730 65.680 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 641.790 1437.040 642.070 1437.320 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 641.765 1437.330 642.095 1437.345 ;
        RECT 641.765 1437.320 660.100 1437.330 ;
        RECT 641.765 1437.030 664.000 1437.320 ;
        RECT 641.765 1437.015 642.095 1437.030 ;
        RECT 660.000 1436.720 664.000 1437.030 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 44.690 1318.080 45.010 1318.140 ;
        RECT 641.770 1318.080 642.090 1318.140 ;
        RECT 44.690 1317.940 642.090 1318.080 ;
        RECT 44.690 1317.880 45.010 1317.940 ;
        RECT 641.770 1317.880 642.090 1317.940 ;
        RECT 17.090 682.620 17.410 682.680 ;
        RECT 44.690 682.620 45.010 682.680 ;
        RECT 17.090 682.480 45.010 682.620 ;
        RECT 17.090 682.420 17.410 682.480 ;
        RECT 44.690 682.420 45.010 682.480 ;
      LAYER via ;
        RECT 44.720 1317.880 44.980 1318.140 ;
        RECT 641.800 1317.880 642.060 1318.140 ;
        RECT 17.120 682.420 17.380 682.680 ;
        RECT 44.720 682.420 44.980 682.680 ;
      LAYER met2 ;
        RECT 641.790 1322.075 642.070 1322.445 ;
        RECT 641.860 1318.170 642.000 1322.075 ;
        RECT 44.720 1317.850 44.980 1318.170 ;
        RECT 641.800 1317.850 642.060 1318.170 ;
        RECT 44.780 682.710 44.920 1317.850 ;
        RECT 17.120 682.390 17.380 682.710 ;
        RECT 44.720 682.390 44.980 682.710 ;
        RECT 17.180 681.885 17.320 682.390 ;
        RECT 17.110 681.515 17.390 681.885 ;
      LAYER via2 ;
        RECT 641.790 1322.120 642.070 1322.400 ;
        RECT 17.110 681.560 17.390 681.840 ;
      LAYER met3 ;
        RECT 641.765 1322.410 642.095 1322.425 ;
        RECT 641.765 1322.400 660.100 1322.410 ;
        RECT 641.765 1322.110 664.000 1322.400 ;
        RECT 641.765 1322.095 642.095 1322.110 ;
        RECT 660.000 1321.800 664.000 1322.110 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.085 681.850 17.415 681.865 ;
        RECT -4.800 681.550 17.415 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 17.085 681.535 17.415 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 1207.580 79.510 1207.640 ;
        RECT 641.770 1207.580 642.090 1207.640 ;
        RECT 79.190 1207.440 642.090 1207.580 ;
        RECT 79.190 1207.380 79.510 1207.440 ;
        RECT 641.770 1207.380 642.090 1207.440 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 79.190 469.100 79.510 469.160 ;
        RECT 17.090 468.960 79.510 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 79.190 468.900 79.510 468.960 ;
      LAYER via ;
        RECT 79.220 1207.380 79.480 1207.640 ;
        RECT 641.800 1207.380 642.060 1207.640 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 79.220 468.900 79.480 469.160 ;
      LAYER met2 ;
        RECT 641.790 1207.835 642.070 1208.205 ;
        RECT 641.860 1207.670 642.000 1207.835 ;
        RECT 79.220 1207.350 79.480 1207.670 ;
        RECT 641.800 1207.350 642.060 1207.670 ;
        RECT 79.280 469.190 79.420 1207.350 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 79.220 468.870 79.480 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 641.790 1207.880 642.070 1208.160 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 641.765 1208.170 642.095 1208.185 ;
        RECT 641.765 1208.160 660.100 1208.170 ;
        RECT 641.765 1207.870 664.000 1208.160 ;
        RECT 641.765 1207.855 642.095 1207.870 ;
        RECT 660.000 1207.560 664.000 1207.870 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 58.490 1090.280 58.810 1090.340 ;
        RECT 641.770 1090.280 642.090 1090.340 ;
        RECT 58.490 1090.140 642.090 1090.280 ;
        RECT 58.490 1090.080 58.810 1090.140 ;
        RECT 641.770 1090.080 642.090 1090.140 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 58.490 255.240 58.810 255.300 ;
        RECT 17.090 255.100 58.810 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 58.490 255.040 58.810 255.100 ;
      LAYER via ;
        RECT 58.520 1090.080 58.780 1090.340 ;
        RECT 641.800 1090.080 642.060 1090.340 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 58.520 255.040 58.780 255.300 ;
      LAYER met2 ;
        RECT 641.790 1093.595 642.070 1093.965 ;
        RECT 641.860 1090.370 642.000 1093.595 ;
        RECT 58.520 1090.050 58.780 1090.370 ;
        RECT 641.800 1090.050 642.060 1090.370 ;
        RECT 58.580 255.330 58.720 1090.050 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 58.520 255.010 58.780 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 641.790 1093.640 642.070 1093.920 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 641.765 1093.930 642.095 1093.945 ;
        RECT 641.765 1093.920 660.100 1093.930 ;
        RECT 641.765 1093.630 664.000 1093.920 ;
        RECT 641.765 1093.615 642.095 1093.630 ;
        RECT 660.000 1093.320 664.000 1093.630 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 30.890 972.980 31.210 973.040 ;
        RECT 643.150 972.980 643.470 973.040 ;
        RECT 30.890 972.840 643.470 972.980 ;
        RECT 30.890 972.780 31.210 972.840 ;
        RECT 643.150 972.780 643.470 972.840 ;
        RECT 13.870 40.700 14.190 40.760 ;
        RECT 30.890 40.700 31.210 40.760 ;
        RECT 13.870 40.560 31.210 40.700 ;
        RECT 13.870 40.500 14.190 40.560 ;
        RECT 30.890 40.500 31.210 40.560 ;
      LAYER via ;
        RECT 30.920 972.780 31.180 973.040 ;
        RECT 643.180 972.780 643.440 973.040 ;
        RECT 13.900 40.500 14.160 40.760 ;
        RECT 30.920 40.500 31.180 40.760 ;
      LAYER met2 ;
        RECT 643.170 979.355 643.450 979.725 ;
        RECT 643.240 973.070 643.380 979.355 ;
        RECT 30.920 972.750 31.180 973.070 ;
        RECT 643.180 972.750 643.440 973.070 ;
        RECT 30.980 40.790 31.120 972.750 ;
        RECT 13.900 40.470 14.160 40.790 ;
        RECT 30.920 40.470 31.180 40.790 ;
        RECT 13.960 35.885 14.100 40.470 ;
        RECT 13.890 35.515 14.170 35.885 ;
      LAYER via2 ;
        RECT 643.170 979.400 643.450 979.680 ;
        RECT 13.890 35.560 14.170 35.840 ;
      LAYER met3 ;
        RECT 643.145 979.690 643.475 979.705 ;
        RECT 643.145 979.680 660.100 979.690 ;
        RECT 643.145 979.390 664.000 979.680 ;
        RECT 643.145 979.375 643.475 979.390 ;
        RECT 660.000 979.080 664.000 979.390 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 13.865 35.850 14.195 35.865 ;
        RECT -4.800 35.550 14.195 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 13.865 35.535 14.195 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2268.330 910.760 2268.650 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2268.330 910.620 2901.150 910.760 ;
        RECT 2268.330 910.560 2268.650 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2268.360 910.560 2268.620 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2268.350 1368.995 2268.630 1369.365 ;
        RECT 2268.420 910.850 2268.560 1368.995 ;
        RECT 2268.360 910.530 2268.620 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2268.350 1369.040 2268.630 1369.320 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2268.325 1369.330 2268.655 1369.345 ;
        RECT 2250.780 1369.320 2268.655 1369.330 ;
        RECT 2247.465 1369.030 2268.655 1369.320 ;
        RECT 2247.465 1368.720 2251.465 1369.030 ;
        RECT 2268.325 1369.015 2268.655 1369.030 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 1145.360 2267.270 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2266.950 1145.220 2901.150 1145.360 ;
        RECT 2266.950 1145.160 2267.270 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2266.980 1145.160 2267.240 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2266.970 1475.755 2267.250 1476.125 ;
        RECT 2267.040 1145.450 2267.180 1475.755 ;
        RECT 2266.980 1145.130 2267.240 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2266.970 1475.800 2267.250 1476.080 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2266.945 1476.090 2267.275 1476.105 ;
        RECT 2250.780 1476.080 2267.275 1476.090 ;
        RECT 2247.465 1475.790 2267.275 1476.080 ;
        RECT 2247.465 1475.480 2251.465 1475.790 ;
        RECT 2266.945 1475.775 2267.275 1475.790 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.870 1379.960 2268.190 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2267.870 1379.820 2901.150 1379.960 ;
        RECT 2267.870 1379.760 2268.190 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2267.900 1379.760 2268.160 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2267.890 1583.195 2268.170 1583.565 ;
        RECT 2267.960 1380.050 2268.100 1583.195 ;
        RECT 2267.900 1379.730 2268.160 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2267.890 1583.240 2268.170 1583.520 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2267.865 1583.530 2268.195 1583.545 ;
        RECT 2250.780 1583.520 2268.195 1583.530 ;
        RECT 2247.465 1583.230 2268.195 1583.520 ;
        RECT 2247.465 1582.920 2251.465 1583.230 ;
        RECT 2267.865 1583.215 2268.195 1583.230 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.410 1614.560 2267.730 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2267.410 1614.420 2901.150 1614.560 ;
        RECT 2267.410 1614.360 2267.730 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2267.440 1614.360 2267.700 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2267.430 1689.955 2267.710 1690.325 ;
        RECT 2267.500 1614.650 2267.640 1689.955 ;
        RECT 2267.440 1614.330 2267.700 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2267.430 1690.000 2267.710 1690.280 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2267.405 1690.290 2267.735 1690.305 ;
        RECT 2250.780 1690.280 2267.735 1690.290 ;
        RECT 2247.465 1689.990 2267.735 1690.280 ;
        RECT 2247.465 1689.680 2251.465 1689.990 ;
        RECT 2267.405 1689.975 2267.735 1689.990 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1800.880 2270.030 1800.940 ;
        RECT 2901.290 1800.880 2901.610 1800.940 ;
        RECT 2269.710 1800.740 2901.610 1800.880 ;
        RECT 2269.710 1800.680 2270.030 1800.740 ;
        RECT 2901.290 1800.680 2901.610 1800.740 ;
      LAYER via ;
        RECT 2269.740 1800.680 2270.000 1800.940 ;
        RECT 2901.320 1800.680 2901.580 1800.940 ;
      LAYER met2 ;
        RECT 2901.310 1847.715 2901.590 1848.085 ;
        RECT 2901.380 1800.970 2901.520 1847.715 ;
        RECT 2269.740 1800.650 2270.000 1800.970 ;
        RECT 2901.320 1800.650 2901.580 1800.970 ;
        RECT 2269.800 1797.085 2269.940 1800.650 ;
        RECT 2269.730 1796.715 2270.010 1797.085 ;
      LAYER via2 ;
        RECT 2901.310 1847.760 2901.590 1848.040 ;
        RECT 2269.730 1796.760 2270.010 1797.040 ;
      LAYER met3 ;
        RECT 2901.285 1848.050 2901.615 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.285 1847.750 2924.800 1848.050 ;
        RECT 2901.285 1847.735 2901.615 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2269.705 1797.050 2270.035 1797.065 ;
        RECT 2250.780 1797.040 2270.035 1797.050 ;
        RECT 2247.465 1796.750 2270.035 1797.040 ;
        RECT 2247.465 1796.440 2251.465 1796.750 ;
        RECT 2269.705 1796.735 2270.035 1796.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1904.240 2270.030 1904.300 ;
        RECT 2894.390 1904.240 2894.710 1904.300 ;
        RECT 2269.710 1904.100 2894.710 1904.240 ;
        RECT 2269.710 1904.040 2270.030 1904.100 ;
        RECT 2894.390 1904.040 2894.710 1904.100 ;
      LAYER via ;
        RECT 2269.740 1904.040 2270.000 1904.300 ;
        RECT 2894.420 1904.040 2894.680 1904.300 ;
      LAYER met2 ;
        RECT 2894.410 2082.315 2894.690 2082.685 ;
        RECT 2894.480 1904.330 2894.620 2082.315 ;
        RECT 2269.740 1904.010 2270.000 1904.330 ;
        RECT 2894.420 1904.010 2894.680 1904.330 ;
        RECT 2269.800 1903.845 2269.940 1904.010 ;
        RECT 2269.730 1903.475 2270.010 1903.845 ;
      LAYER via2 ;
        RECT 2894.410 2082.360 2894.690 2082.640 ;
        RECT 2269.730 1903.520 2270.010 1903.800 ;
      LAYER met3 ;
        RECT 2894.385 2082.650 2894.715 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2894.385 2082.350 2924.800 2082.650 ;
        RECT 2894.385 2082.335 2894.715 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2269.705 1903.810 2270.035 1903.825 ;
        RECT 2250.780 1903.800 2270.035 1903.810 ;
        RECT 2247.465 1903.510 2270.035 1903.800 ;
        RECT 2247.465 1903.200 2251.465 1903.510 ;
        RECT 2269.705 1903.495 2270.035 1903.510 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2714.990 2311.900 2715.310 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2714.990 2311.760 2901.150 2311.900 ;
        RECT 2714.990 2311.700 2715.310 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 2269.710 2014.740 2270.030 2014.800 ;
        RECT 2714.990 2014.740 2715.310 2014.800 ;
        RECT 2269.710 2014.600 2715.310 2014.740 ;
        RECT 2269.710 2014.540 2270.030 2014.600 ;
        RECT 2714.990 2014.540 2715.310 2014.600 ;
      LAYER via ;
        RECT 2715.020 2311.700 2715.280 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 2269.740 2014.540 2270.000 2014.800 ;
        RECT 2715.020 2014.540 2715.280 2014.800 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2715.020 2311.670 2715.280 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2715.080 2014.830 2715.220 2311.670 ;
        RECT 2269.740 2014.510 2270.000 2014.830 ;
        RECT 2715.020 2014.510 2715.280 2014.830 ;
        RECT 2269.800 2010.605 2269.940 2014.510 ;
        RECT 2269.730 2010.235 2270.010 2010.605 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2269.730 2010.280 2270.010 2010.560 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2269.705 2010.570 2270.035 2010.585 ;
        RECT 2250.780 2010.560 2270.035 2010.570 ;
        RECT 2247.465 2010.270 2270.035 2010.560 ;
        RECT 2247.465 2009.960 2251.465 2010.270 ;
        RECT 2269.705 2010.255 2270.035 2010.270 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.490 151.540 2266.810 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2266.490 151.400 2901.150 151.540 ;
        RECT 2266.490 151.340 2266.810 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2266.520 151.340 2266.780 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2266.510 1013.355 2266.790 1013.725 ;
        RECT 2266.580 151.630 2266.720 1013.355 ;
        RECT 2266.520 151.310 2266.780 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2266.510 1013.400 2266.790 1013.680 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2266.485 1013.690 2266.815 1013.705 ;
        RECT 2250.780 1013.680 2266.815 1013.690 ;
        RECT 2247.465 1013.390 2266.815 1013.680 ;
        RECT 2247.465 1013.080 2251.465 1013.390 ;
        RECT 2266.485 1013.375 2266.815 1013.390 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2300.990 2491.080 2301.310 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2300.990 2490.940 2901.150 2491.080 ;
        RECT 2300.990 2490.880 2301.310 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 2269.710 2082.060 2270.030 2082.120 ;
        RECT 2300.990 2082.060 2301.310 2082.120 ;
        RECT 2269.710 2081.920 2301.310 2082.060 ;
        RECT 2269.710 2081.860 2270.030 2081.920 ;
        RECT 2300.990 2081.860 2301.310 2081.920 ;
      LAYER via ;
        RECT 2301.020 2490.880 2301.280 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 2269.740 2081.860 2270.000 2082.120 ;
        RECT 2301.020 2081.860 2301.280 2082.120 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2301.020 2490.850 2301.280 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2301.080 2082.150 2301.220 2490.850 ;
        RECT 2269.740 2082.005 2270.000 2082.150 ;
        RECT 2269.730 2081.635 2270.010 2082.005 ;
        RECT 2301.020 2081.830 2301.280 2082.150 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2269.730 2081.680 2270.010 2081.960 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2269.705 2081.970 2270.035 2081.985 ;
        RECT 2250.780 2081.960 2270.035 2081.970 ;
        RECT 2247.465 2081.670 2270.035 2081.960 ;
        RECT 2247.465 2081.360 2251.465 2081.670 ;
        RECT 2269.705 2081.655 2270.035 2081.670 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.490 2725.680 2404.810 2725.740 ;
        RECT 2899.450 2725.680 2899.770 2725.740 ;
        RECT 2404.490 2725.540 2899.770 2725.680 ;
        RECT 2404.490 2725.480 2404.810 2725.540 ;
        RECT 2899.450 2725.480 2899.770 2725.540 ;
        RECT 2268.790 2194.260 2269.110 2194.320 ;
        RECT 2404.490 2194.260 2404.810 2194.320 ;
        RECT 2268.790 2194.120 2404.810 2194.260 ;
        RECT 2268.790 2194.060 2269.110 2194.120 ;
        RECT 2404.490 2194.060 2404.810 2194.120 ;
      LAYER via ;
        RECT 2404.520 2725.480 2404.780 2725.740 ;
        RECT 2899.480 2725.480 2899.740 2725.740 ;
        RECT 2268.820 2194.060 2269.080 2194.320 ;
        RECT 2404.520 2194.060 2404.780 2194.320 ;
      LAYER met2 ;
        RECT 2899.470 2727.635 2899.750 2728.005 ;
        RECT 2899.540 2725.770 2899.680 2727.635 ;
        RECT 2404.520 2725.450 2404.780 2725.770 ;
        RECT 2899.480 2725.450 2899.740 2725.770 ;
        RECT 2404.580 2194.350 2404.720 2725.450 ;
        RECT 2268.820 2194.030 2269.080 2194.350 ;
        RECT 2404.520 2194.030 2404.780 2194.350 ;
        RECT 2268.880 2188.765 2269.020 2194.030 ;
        RECT 2268.810 2188.395 2269.090 2188.765 ;
      LAYER via2 ;
        RECT 2899.470 2727.680 2899.750 2727.960 ;
        RECT 2268.810 2188.440 2269.090 2188.720 ;
      LAYER met3 ;
        RECT 2899.445 2727.970 2899.775 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2899.445 2727.670 2924.800 2727.970 ;
        RECT 2899.445 2727.655 2899.775 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2268.785 2188.730 2269.115 2188.745 ;
        RECT 2250.780 2188.720 2269.115 2188.730 ;
        RECT 2247.465 2188.430 2269.115 2188.720 ;
        RECT 2247.465 2188.120 2251.465 2188.430 ;
        RECT 2268.785 2188.415 2269.115 2188.430 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2411.390 2960.280 2411.710 2960.340 ;
        RECT 2899.450 2960.280 2899.770 2960.340 ;
        RECT 2411.390 2960.140 2899.770 2960.280 ;
        RECT 2411.390 2960.080 2411.710 2960.140 ;
        RECT 2899.450 2960.080 2899.770 2960.140 ;
        RECT 2266.950 2297.620 2267.270 2297.680 ;
        RECT 2411.390 2297.620 2411.710 2297.680 ;
        RECT 2266.950 2297.480 2411.710 2297.620 ;
        RECT 2266.950 2297.420 2267.270 2297.480 ;
        RECT 2411.390 2297.420 2411.710 2297.480 ;
      LAYER via ;
        RECT 2411.420 2960.080 2411.680 2960.340 ;
        RECT 2899.480 2960.080 2899.740 2960.340 ;
        RECT 2266.980 2297.420 2267.240 2297.680 ;
        RECT 2411.420 2297.420 2411.680 2297.680 ;
      LAYER met2 ;
        RECT 2899.470 2962.235 2899.750 2962.605 ;
        RECT 2899.540 2960.370 2899.680 2962.235 ;
        RECT 2411.420 2960.050 2411.680 2960.370 ;
        RECT 2899.480 2960.050 2899.740 2960.370 ;
        RECT 2411.480 2297.710 2411.620 2960.050 ;
        RECT 2266.980 2297.390 2267.240 2297.710 ;
        RECT 2411.420 2297.390 2411.680 2297.710 ;
        RECT 2267.040 2295.525 2267.180 2297.390 ;
        RECT 2266.970 2295.155 2267.250 2295.525 ;
      LAYER via2 ;
        RECT 2899.470 2962.280 2899.750 2962.560 ;
        RECT 2266.970 2295.200 2267.250 2295.480 ;
      LAYER met3 ;
        RECT 2899.445 2962.570 2899.775 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2899.445 2962.270 2924.800 2962.570 ;
        RECT 2899.445 2962.255 2899.775 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2266.945 2295.490 2267.275 2295.505 ;
        RECT 2250.780 2295.480 2267.275 2295.490 ;
        RECT 2247.465 2295.190 2267.275 2295.480 ;
        RECT 2247.465 2294.880 2251.465 2295.190 ;
        RECT 2266.945 2295.175 2267.275 2295.190 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2268.790 2408.120 2269.110 2408.180 ;
        RECT 2901.750 2408.120 2902.070 2408.180 ;
        RECT 2268.790 2407.980 2902.070 2408.120 ;
        RECT 2268.790 2407.920 2269.110 2407.980 ;
        RECT 2901.750 2407.920 2902.070 2407.980 ;
      LAYER via ;
        RECT 2268.820 2407.920 2269.080 2408.180 ;
        RECT 2901.780 2407.920 2902.040 2408.180 ;
      LAYER met2 ;
        RECT 2901.770 3196.835 2902.050 3197.205 ;
        RECT 2901.840 2408.210 2901.980 3196.835 ;
        RECT 2268.820 2407.890 2269.080 2408.210 ;
        RECT 2901.780 2407.890 2902.040 2408.210 ;
        RECT 2268.880 2402.285 2269.020 2407.890 ;
        RECT 2268.810 2401.915 2269.090 2402.285 ;
      LAYER via2 ;
        RECT 2901.770 3196.880 2902.050 3197.160 ;
        RECT 2268.810 2401.960 2269.090 2402.240 ;
      LAYER met3 ;
        RECT 2901.745 3197.170 2902.075 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.745 3196.870 2924.800 3197.170 ;
        RECT 2901.745 3196.855 2902.075 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2268.785 2402.250 2269.115 2402.265 ;
        RECT 2250.780 2402.240 2269.115 2402.250 ;
        RECT 2247.465 2401.950 2269.115 2402.240 ;
        RECT 2247.465 2401.640 2251.465 2401.950 ;
        RECT 2268.785 2401.935 2269.115 2401.950 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 2511.480 2267.270 2511.540 ;
        RECT 2901.290 2511.480 2901.610 2511.540 ;
        RECT 2266.950 2511.340 2901.610 2511.480 ;
        RECT 2266.950 2511.280 2267.270 2511.340 ;
        RECT 2901.290 2511.280 2901.610 2511.340 ;
      LAYER via ;
        RECT 2266.980 2511.280 2267.240 2511.540 ;
        RECT 2901.320 2511.280 2901.580 2511.540 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 2901.380 2511.570 2901.520 3431.435 ;
        RECT 2266.980 2511.250 2267.240 2511.570 ;
        RECT 2901.320 2511.250 2901.580 2511.570 ;
        RECT 2267.040 2509.045 2267.180 2511.250 ;
        RECT 2266.970 2508.675 2267.250 2509.045 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
        RECT 2266.970 2508.720 2267.250 2509.000 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2266.945 2509.010 2267.275 2509.025 ;
        RECT 2250.780 2509.000 2267.275 2509.010 ;
        RECT 2247.465 2508.710 2267.275 2509.000 ;
        RECT 2247.465 2508.400 2251.465 2508.710 ;
        RECT 2266.945 2508.695 2267.275 2508.710 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3415.555 ;
        RECT 2712.765 3008.405 2712.935 3042.915 ;
        RECT 2713.685 2946.525 2713.855 2994.635 ;
        RECT 2712.305 2753.065 2712.475 2801.175 ;
      LAYER mcon ;
        RECT 2713.685 3415.385 2713.855 3415.555 ;
        RECT 2712.765 3042.745 2712.935 3042.915 ;
        RECT 2713.685 2994.465 2713.855 2994.635 ;
        RECT 2712.305 2801.005 2712.475 2801.175 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2712.690 3470.620 2713.010 3470.680 ;
        RECT 2713.610 3470.620 2713.930 3470.680 ;
        RECT 2712.690 3470.480 2713.930 3470.620 ;
        RECT 2712.690 3470.420 2713.010 3470.480 ;
        RECT 2713.610 3470.420 2713.930 3470.480 ;
        RECT 2712.690 3463.820 2713.010 3463.880 ;
        RECT 2713.610 3463.820 2713.930 3463.880 ;
        RECT 2712.690 3463.680 2713.930 3463.820 ;
        RECT 2712.690 3463.620 2713.010 3463.680 ;
        RECT 2713.610 3463.620 2713.930 3463.680 ;
        RECT 2711.770 3415.540 2712.090 3415.600 ;
        RECT 2713.625 3415.540 2713.915 3415.585 ;
        RECT 2711.770 3415.400 2713.915 3415.540 ;
        RECT 2711.770 3415.340 2712.090 3415.400 ;
        RECT 2713.625 3415.355 2713.915 3415.400 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2712.690 3042.900 2713.010 3042.960 ;
        RECT 2712.495 3042.760 2713.010 3042.900 ;
        RECT 2712.690 3042.700 2713.010 3042.760 ;
        RECT 2712.705 3008.560 2712.995 3008.605 ;
        RECT 2713.610 3008.560 2713.930 3008.620 ;
        RECT 2712.705 3008.420 2713.930 3008.560 ;
        RECT 2712.705 3008.375 2712.995 3008.420 ;
        RECT 2713.610 3008.360 2713.930 3008.420 ;
        RECT 2713.610 2994.620 2713.930 2994.680 ;
        RECT 2713.415 2994.480 2713.930 2994.620 ;
        RECT 2713.610 2994.420 2713.930 2994.480 ;
        RECT 2713.625 2946.680 2713.915 2946.725 ;
        RECT 2714.070 2946.680 2714.390 2946.740 ;
        RECT 2713.625 2946.540 2714.390 2946.680 ;
        RECT 2713.625 2946.495 2713.915 2946.540 ;
        RECT 2714.070 2946.480 2714.390 2946.540 ;
        RECT 2714.070 2912.340 2714.390 2912.400 ;
        RECT 2713.700 2912.200 2714.390 2912.340 ;
        RECT 2713.700 2911.720 2713.840 2912.200 ;
        RECT 2714.070 2912.140 2714.390 2912.200 ;
        RECT 2713.610 2911.460 2713.930 2911.720 ;
        RECT 2712.230 2815.580 2712.550 2815.840 ;
        RECT 2712.320 2815.160 2712.460 2815.580 ;
        RECT 2712.230 2814.900 2712.550 2815.160 ;
        RECT 2712.230 2801.160 2712.550 2801.220 ;
        RECT 2712.035 2801.020 2712.550 2801.160 ;
        RECT 2712.230 2800.960 2712.550 2801.020 ;
        RECT 2712.245 2753.220 2712.535 2753.265 ;
        RECT 2713.150 2753.220 2713.470 2753.280 ;
        RECT 2712.245 2753.080 2713.470 2753.220 ;
        RECT 2712.245 2753.035 2712.535 2753.080 ;
        RECT 2713.150 2753.020 2713.470 2753.080 ;
        RECT 2712.230 2718.200 2712.550 2718.260 ;
        RECT 2713.150 2718.200 2713.470 2718.260 ;
        RECT 2712.230 2718.060 2713.470 2718.200 ;
        RECT 2712.230 2718.000 2712.550 2718.060 ;
        RECT 2713.150 2718.000 2713.470 2718.060 ;
        RECT 2162.990 2577.440 2163.310 2577.500 ;
        RECT 2713.150 2577.440 2713.470 2577.500 ;
        RECT 2162.990 2577.300 2713.470 2577.440 ;
        RECT 2162.990 2577.240 2163.310 2577.300 ;
        RECT 2713.150 2577.240 2713.470 2577.300 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2712.720 3470.420 2712.980 3470.680 ;
        RECT 2713.640 3470.420 2713.900 3470.680 ;
        RECT 2712.720 3463.620 2712.980 3463.880 ;
        RECT 2713.640 3463.620 2713.900 3463.880 ;
        RECT 2711.800 3415.340 2712.060 3415.600 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2712.720 3042.700 2712.980 3042.960 ;
        RECT 2713.640 3008.360 2713.900 3008.620 ;
        RECT 2713.640 2994.420 2713.900 2994.680 ;
        RECT 2714.100 2946.480 2714.360 2946.740 ;
        RECT 2714.100 2912.140 2714.360 2912.400 ;
        RECT 2713.640 2911.460 2713.900 2911.720 ;
        RECT 2712.260 2815.580 2712.520 2815.840 ;
        RECT 2712.260 2814.900 2712.520 2815.160 ;
        RECT 2712.260 2800.960 2712.520 2801.220 ;
        RECT 2713.180 2753.020 2713.440 2753.280 ;
        RECT 2712.260 2718.000 2712.520 2718.260 ;
        RECT 2713.180 2718.000 2713.440 2718.260 ;
        RECT 2163.020 2577.240 2163.280 2577.500 ;
        RECT 2713.180 2577.240 2713.440 2577.500 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3470.710 2713.840 3491.130 ;
        RECT 2712.720 3470.390 2712.980 3470.710 ;
        RECT 2713.640 3470.390 2713.900 3470.710 ;
        RECT 2712.780 3463.910 2712.920 3470.390 ;
        RECT 2712.720 3463.590 2712.980 3463.910 ;
        RECT 2713.640 3463.590 2713.900 3463.910 ;
        RECT 2713.700 3416.165 2713.840 3463.590 ;
        RECT 2711.790 3415.795 2712.070 3416.165 ;
        RECT 2713.630 3415.795 2713.910 3416.165 ;
        RECT 2711.860 3415.630 2712.000 3415.795 ;
        RECT 2711.800 3415.310 2712.060 3415.630 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3056.330 2712.460 3056.610 ;
        RECT 2712.320 3056.190 2712.920 3056.330 ;
        RECT 2712.780 3042.990 2712.920 3056.190 ;
        RECT 2712.720 3042.670 2712.980 3042.990 ;
        RECT 2713.640 3008.330 2713.900 3008.650 ;
        RECT 2713.700 2994.710 2713.840 3008.330 ;
        RECT 2713.640 2994.390 2713.900 2994.710 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.250 2712.460 2814.870 ;
        RECT 2712.260 2800.930 2712.520 2801.250 ;
        RECT 2713.180 2752.990 2713.440 2753.310 ;
        RECT 2713.240 2718.290 2713.380 2752.990 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2713.180 2717.970 2713.440 2718.290 ;
        RECT 2712.320 2670.090 2712.460 2717.970 ;
        RECT 2712.320 2669.950 2712.920 2670.090 ;
        RECT 2712.780 2622.490 2712.920 2669.950 ;
        RECT 2712.780 2622.350 2713.380 2622.490 ;
        RECT 2713.240 2577.530 2713.380 2622.350 ;
        RECT 2163.020 2577.210 2163.280 2577.530 ;
        RECT 2713.180 2577.210 2713.440 2577.530 ;
        RECT 2163.080 2562.185 2163.220 2577.210 ;
        RECT 2162.910 2561.900 2163.220 2562.185 ;
        RECT 2162.910 2558.185 2163.190 2561.900 ;
      LAYER via2 ;
        RECT 2711.790 3415.840 2712.070 3416.120 ;
        RECT 2713.630 3415.840 2713.910 3416.120 ;
      LAYER met3 ;
        RECT 2711.765 3416.130 2712.095 3416.145 ;
        RECT 2713.605 3416.130 2713.935 3416.145 ;
        RECT 2711.765 3415.830 2713.935 3416.130 ;
        RECT 2711.765 3415.815 2712.095 3415.830 ;
        RECT 2713.605 3415.815 2713.935 3415.830 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2387.545 2898.245 2387.715 2946.355 ;
        RECT 2388.005 2815.285 2388.175 2849.455 ;
      LAYER mcon ;
        RECT 2387.545 2946.185 2387.715 2946.355 ;
        RECT 2388.005 2849.285 2388.175 2849.455 ;
      LAYER met1 ;
        RECT 2387.470 3464.160 2387.790 3464.220 ;
        RECT 2392.990 3464.160 2393.310 3464.220 ;
        RECT 2387.470 3464.020 2393.310 3464.160 ;
        RECT 2387.470 3463.960 2387.790 3464.020 ;
        RECT 2392.990 3463.960 2393.310 3464.020 ;
        RECT 2387.470 3367.600 2387.790 3367.660 ;
        RECT 2388.390 3367.600 2388.710 3367.660 ;
        RECT 2387.470 3367.460 2388.710 3367.600 ;
        RECT 2387.470 3367.400 2387.790 3367.460 ;
        RECT 2388.390 3367.400 2388.710 3367.460 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 2387.470 3077.580 2387.790 3077.640 ;
        RECT 2388.390 3077.580 2388.710 3077.640 ;
        RECT 2387.470 3077.440 2388.710 3077.580 ;
        RECT 2387.470 3077.380 2387.790 3077.440 ;
        RECT 2388.390 3077.380 2388.710 3077.440 ;
        RECT 2387.470 2981.020 2387.790 2981.080 ;
        RECT 2388.390 2981.020 2388.710 2981.080 ;
        RECT 2387.470 2980.880 2388.710 2981.020 ;
        RECT 2387.470 2980.820 2387.790 2980.880 ;
        RECT 2388.390 2980.820 2388.710 2980.880 ;
        RECT 2387.485 2946.340 2387.775 2946.385 ;
        RECT 2387.930 2946.340 2388.250 2946.400 ;
        RECT 2387.485 2946.200 2388.250 2946.340 ;
        RECT 2387.485 2946.155 2387.775 2946.200 ;
        RECT 2387.930 2946.140 2388.250 2946.200 ;
        RECT 2387.470 2898.400 2387.790 2898.460 ;
        RECT 2387.275 2898.260 2387.790 2898.400 ;
        RECT 2387.470 2898.200 2387.790 2898.260 ;
        RECT 2387.930 2849.440 2388.250 2849.500 ;
        RECT 2387.735 2849.300 2388.250 2849.440 ;
        RECT 2387.930 2849.240 2388.250 2849.300 ;
        RECT 2387.945 2815.440 2388.235 2815.485 ;
        RECT 2388.850 2815.440 2389.170 2815.500 ;
        RECT 2387.945 2815.300 2389.170 2815.440 ;
        RECT 2387.945 2815.255 2388.235 2815.300 ;
        RECT 2388.850 2815.240 2389.170 2815.300 ;
        RECT 2387.930 2753.220 2388.250 2753.280 ;
        RECT 2389.310 2753.220 2389.630 2753.280 ;
        RECT 2387.930 2753.080 2389.630 2753.220 ;
        RECT 2387.930 2753.020 2388.250 2753.080 ;
        RECT 2389.310 2753.020 2389.630 2753.080 ;
        RECT 2389.310 2719.220 2389.630 2719.280 ;
        RECT 2388.940 2719.080 2389.630 2719.220 ;
        RECT 2388.940 2718.600 2389.080 2719.080 ;
        RECT 2389.310 2719.020 2389.630 2719.080 ;
        RECT 2388.850 2718.340 2389.170 2718.600 ;
        RECT 2387.930 2656.660 2388.250 2656.720 ;
        RECT 2389.310 2656.660 2389.630 2656.720 ;
        RECT 2387.930 2656.520 2389.630 2656.660 ;
        RECT 2387.930 2656.460 2388.250 2656.520 ;
        RECT 2389.310 2656.460 2389.630 2656.520 ;
        RECT 2388.390 2608.380 2388.710 2608.440 ;
        RECT 2389.310 2608.380 2389.630 2608.440 ;
        RECT 2388.390 2608.240 2389.630 2608.380 ;
        RECT 2388.390 2608.180 2388.710 2608.240 ;
        RECT 2389.310 2608.180 2389.630 2608.240 ;
        RECT 1986.350 2578.460 1986.670 2578.520 ;
        RECT 2388.390 2578.460 2388.710 2578.520 ;
        RECT 1986.350 2578.320 2388.710 2578.460 ;
        RECT 1986.350 2578.260 1986.670 2578.320 ;
        RECT 2388.390 2578.260 2388.710 2578.320 ;
      LAYER via ;
        RECT 2387.500 3463.960 2387.760 3464.220 ;
        RECT 2393.020 3463.960 2393.280 3464.220 ;
        RECT 2387.500 3367.400 2387.760 3367.660 ;
        RECT 2388.420 3367.400 2388.680 3367.660 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 2387.500 3077.380 2387.760 3077.640 ;
        RECT 2388.420 3077.380 2388.680 3077.640 ;
        RECT 2387.500 2980.820 2387.760 2981.080 ;
        RECT 2388.420 2980.820 2388.680 2981.080 ;
        RECT 2387.960 2946.140 2388.220 2946.400 ;
        RECT 2387.500 2898.200 2387.760 2898.460 ;
        RECT 2387.960 2849.240 2388.220 2849.500 ;
        RECT 2388.880 2815.240 2389.140 2815.500 ;
        RECT 2387.960 2753.020 2388.220 2753.280 ;
        RECT 2389.340 2753.020 2389.600 2753.280 ;
        RECT 2389.340 2719.020 2389.600 2719.280 ;
        RECT 2388.880 2718.340 2389.140 2718.600 ;
        RECT 2387.960 2656.460 2388.220 2656.720 ;
        RECT 2389.340 2656.460 2389.600 2656.720 ;
        RECT 2388.420 2608.180 2388.680 2608.440 ;
        RECT 2389.340 2608.180 2389.600 2608.440 ;
        RECT 1986.380 2578.260 1986.640 2578.520 ;
        RECT 2388.420 2578.260 2388.680 2578.520 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3464.250 2393.220 3517.230 ;
        RECT 2387.500 3463.930 2387.760 3464.250 ;
        RECT 2393.020 3463.930 2393.280 3464.250 ;
        RECT 2387.560 3415.370 2387.700 3463.930 ;
        RECT 2387.560 3415.230 2388.620 3415.370 ;
        RECT 2388.480 3367.690 2388.620 3415.230 ;
        RECT 2387.500 3367.370 2387.760 3367.690 ;
        RECT 2388.420 3367.370 2388.680 3367.690 ;
        RECT 2387.560 3318.810 2387.700 3367.370 ;
        RECT 2387.560 3318.670 2388.620 3318.810 ;
        RECT 2388.480 3270.790 2388.620 3318.670 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3077.670 2388.620 3125.550 ;
        RECT 2387.500 3077.350 2387.760 3077.670 ;
        RECT 2388.420 3077.350 2388.680 3077.670 ;
        RECT 2387.560 3029.130 2387.700 3077.350 ;
        RECT 2387.560 3028.990 2388.620 3029.130 ;
        RECT 2388.480 2981.110 2388.620 3028.990 ;
        RECT 2387.500 2980.850 2387.760 2981.110 ;
        RECT 2387.500 2980.790 2388.160 2980.850 ;
        RECT 2388.420 2980.790 2388.680 2981.110 ;
        RECT 2387.560 2980.710 2388.160 2980.790 ;
        RECT 2388.020 2980.170 2388.160 2980.710 ;
        RECT 2388.020 2980.030 2388.620 2980.170 ;
        RECT 2388.480 2959.770 2388.620 2980.030 ;
        RECT 2388.020 2959.630 2388.620 2959.770 ;
        RECT 2388.020 2946.430 2388.160 2959.630 ;
        RECT 2387.960 2946.110 2388.220 2946.430 ;
        RECT 2387.500 2898.170 2387.760 2898.490 ;
        RECT 2387.560 2863.210 2387.700 2898.170 ;
        RECT 2387.560 2863.070 2388.160 2863.210 ;
        RECT 2388.020 2849.530 2388.160 2863.070 ;
        RECT 2387.960 2849.210 2388.220 2849.530 ;
        RECT 2388.880 2815.210 2389.140 2815.530 ;
        RECT 2388.940 2801.445 2389.080 2815.210 ;
        RECT 2387.950 2801.075 2388.230 2801.445 ;
        RECT 2388.870 2801.075 2389.150 2801.445 ;
        RECT 2388.020 2753.310 2388.160 2801.075 ;
        RECT 2387.960 2752.990 2388.220 2753.310 ;
        RECT 2389.340 2752.990 2389.600 2753.310 ;
        RECT 2389.400 2719.310 2389.540 2752.990 ;
        RECT 2389.340 2718.990 2389.600 2719.310 ;
        RECT 2388.880 2718.310 2389.140 2718.630 ;
        RECT 2388.940 2704.885 2389.080 2718.310 ;
        RECT 2387.950 2704.515 2388.230 2704.885 ;
        RECT 2388.870 2704.515 2389.150 2704.885 ;
        RECT 2388.020 2656.750 2388.160 2704.515 ;
        RECT 2387.960 2656.430 2388.220 2656.750 ;
        RECT 2389.340 2656.430 2389.600 2656.750 ;
        RECT 2389.400 2608.470 2389.540 2656.430 ;
        RECT 2388.420 2608.150 2388.680 2608.470 ;
        RECT 2389.340 2608.150 2389.600 2608.470 ;
        RECT 2388.480 2578.550 2388.620 2608.150 ;
        RECT 1986.380 2578.230 1986.640 2578.550 ;
        RECT 2388.420 2578.230 2388.680 2578.550 ;
        RECT 1986.440 2562.185 1986.580 2578.230 ;
        RECT 1986.270 2561.900 1986.580 2562.185 ;
        RECT 1986.270 2558.185 1986.550 2561.900 ;
      LAYER via2 ;
        RECT 2387.950 2801.120 2388.230 2801.400 ;
        RECT 2388.870 2801.120 2389.150 2801.400 ;
        RECT 2387.950 2704.560 2388.230 2704.840 ;
        RECT 2388.870 2704.560 2389.150 2704.840 ;
      LAYER met3 ;
        RECT 2387.925 2801.410 2388.255 2801.425 ;
        RECT 2388.845 2801.410 2389.175 2801.425 ;
        RECT 2387.925 2801.110 2389.175 2801.410 ;
        RECT 2387.925 2801.095 2388.255 2801.110 ;
        RECT 2388.845 2801.095 2389.175 2801.110 ;
        RECT 2387.925 2704.850 2388.255 2704.865 ;
        RECT 2388.845 2704.850 2389.175 2704.865 ;
        RECT 2387.925 2704.550 2389.175 2704.850 ;
        RECT 2387.925 2704.535 2388.255 2704.550 ;
        RECT 2388.845 2704.535 2389.175 2704.550 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2063.245 3416.065 2063.415 3463.835 ;
        RECT 2065.085 3332.765 2065.255 3415.555 ;
        RECT 2064.165 3008.405 2064.335 3042.915 ;
        RECT 2065.085 2946.525 2065.255 2994.635 ;
        RECT 2063.705 2753.065 2063.875 2801.175 ;
      LAYER mcon ;
        RECT 2063.245 3463.665 2063.415 3463.835 ;
        RECT 2065.085 3415.385 2065.255 3415.555 ;
        RECT 2064.165 3042.745 2064.335 3042.915 ;
        RECT 2065.085 2994.465 2065.255 2994.635 ;
        RECT 2063.705 2801.005 2063.875 2801.175 ;
      LAYER met1 ;
        RECT 2065.010 3491.360 2065.330 3491.420 ;
        RECT 2068.690 3491.360 2069.010 3491.420 ;
        RECT 2065.010 3491.220 2069.010 3491.360 ;
        RECT 2065.010 3491.160 2065.330 3491.220 ;
        RECT 2068.690 3491.160 2069.010 3491.220 ;
        RECT 2064.090 3470.620 2064.410 3470.680 ;
        RECT 2065.010 3470.620 2065.330 3470.680 ;
        RECT 2064.090 3470.480 2065.330 3470.620 ;
        RECT 2064.090 3470.420 2064.410 3470.480 ;
        RECT 2065.010 3470.420 2065.330 3470.480 ;
        RECT 2063.185 3463.820 2063.475 3463.865 ;
        RECT 2064.090 3463.820 2064.410 3463.880 ;
        RECT 2063.185 3463.680 2064.410 3463.820 ;
        RECT 2063.185 3463.635 2063.475 3463.680 ;
        RECT 2064.090 3463.620 2064.410 3463.680 ;
        RECT 2063.170 3416.220 2063.490 3416.280 ;
        RECT 2063.170 3416.080 2063.685 3416.220 ;
        RECT 2063.170 3416.020 2063.490 3416.080 ;
        RECT 2063.170 3415.540 2063.490 3415.600 ;
        RECT 2065.025 3415.540 2065.315 3415.585 ;
        RECT 2063.170 3415.400 2065.315 3415.540 ;
        RECT 2063.170 3415.340 2063.490 3415.400 ;
        RECT 2065.025 3415.355 2065.315 3415.400 ;
        RECT 2065.025 3332.920 2065.315 3332.965 ;
        RECT 2065.470 3332.920 2065.790 3332.980 ;
        RECT 2065.025 3332.780 2065.790 3332.920 ;
        RECT 2065.025 3332.735 2065.315 3332.780 ;
        RECT 2065.470 3332.720 2065.790 3332.780 ;
        RECT 2064.090 3236.360 2064.410 3236.420 ;
        RECT 2064.550 3236.360 2064.870 3236.420 ;
        RECT 2064.090 3236.220 2064.870 3236.360 ;
        RECT 2064.090 3236.160 2064.410 3236.220 ;
        RECT 2064.550 3236.160 2064.870 3236.220 ;
        RECT 2064.090 3202.020 2064.410 3202.080 ;
        RECT 2064.550 3202.020 2064.870 3202.080 ;
        RECT 2064.090 3201.880 2064.870 3202.020 ;
        RECT 2064.090 3201.820 2064.410 3201.880 ;
        RECT 2064.550 3201.820 2064.870 3201.880 ;
        RECT 2063.630 3153.400 2063.950 3153.460 ;
        RECT 2064.550 3153.400 2064.870 3153.460 ;
        RECT 2063.630 3153.260 2064.870 3153.400 ;
        RECT 2063.630 3153.200 2063.950 3153.260 ;
        RECT 2064.550 3153.200 2064.870 3153.260 ;
        RECT 2063.630 3056.840 2063.950 3056.900 ;
        RECT 2064.550 3056.840 2064.870 3056.900 ;
        RECT 2063.630 3056.700 2064.870 3056.840 ;
        RECT 2063.630 3056.640 2063.950 3056.700 ;
        RECT 2064.550 3056.640 2064.870 3056.700 ;
        RECT 2064.090 3042.900 2064.410 3042.960 ;
        RECT 2063.895 3042.760 2064.410 3042.900 ;
        RECT 2064.090 3042.700 2064.410 3042.760 ;
        RECT 2064.105 3008.560 2064.395 3008.605 ;
        RECT 2065.010 3008.560 2065.330 3008.620 ;
        RECT 2064.105 3008.420 2065.330 3008.560 ;
        RECT 2064.105 3008.375 2064.395 3008.420 ;
        RECT 2065.010 3008.360 2065.330 3008.420 ;
        RECT 2065.010 2994.620 2065.330 2994.680 ;
        RECT 2064.815 2994.480 2065.330 2994.620 ;
        RECT 2065.010 2994.420 2065.330 2994.480 ;
        RECT 2065.025 2946.680 2065.315 2946.725 ;
        RECT 2065.470 2946.680 2065.790 2946.740 ;
        RECT 2065.025 2946.540 2065.790 2946.680 ;
        RECT 2065.025 2946.495 2065.315 2946.540 ;
        RECT 2065.470 2946.480 2065.790 2946.540 ;
        RECT 2065.470 2912.340 2065.790 2912.400 ;
        RECT 2065.100 2912.200 2065.790 2912.340 ;
        RECT 2065.100 2911.720 2065.240 2912.200 ;
        RECT 2065.470 2912.140 2065.790 2912.200 ;
        RECT 2065.010 2911.460 2065.330 2911.720 ;
        RECT 2063.630 2815.580 2063.950 2815.840 ;
        RECT 2063.720 2815.160 2063.860 2815.580 ;
        RECT 2063.630 2814.900 2063.950 2815.160 ;
        RECT 2063.630 2801.160 2063.950 2801.220 ;
        RECT 2063.435 2801.020 2063.950 2801.160 ;
        RECT 2063.630 2800.960 2063.950 2801.020 ;
        RECT 2063.645 2753.220 2063.935 2753.265 ;
        RECT 2064.550 2753.220 2064.870 2753.280 ;
        RECT 2063.645 2753.080 2064.870 2753.220 ;
        RECT 2063.645 2753.035 2063.935 2753.080 ;
        RECT 2064.550 2753.020 2064.870 2753.080 ;
        RECT 2063.630 2718.200 2063.950 2718.260 ;
        RECT 2064.550 2718.200 2064.870 2718.260 ;
        RECT 2063.630 2718.060 2064.870 2718.200 ;
        RECT 2063.630 2718.000 2063.950 2718.060 ;
        RECT 2064.550 2718.000 2064.870 2718.060 ;
        RECT 1809.250 2577.440 1809.570 2577.500 ;
        RECT 2064.550 2577.440 2064.870 2577.500 ;
        RECT 1809.250 2577.300 2064.870 2577.440 ;
        RECT 1809.250 2577.240 1809.570 2577.300 ;
        RECT 2064.550 2577.240 2064.870 2577.300 ;
      LAYER via ;
        RECT 2065.040 3491.160 2065.300 3491.420 ;
        RECT 2068.720 3491.160 2068.980 3491.420 ;
        RECT 2064.120 3470.420 2064.380 3470.680 ;
        RECT 2065.040 3470.420 2065.300 3470.680 ;
        RECT 2064.120 3463.620 2064.380 3463.880 ;
        RECT 2063.200 3416.020 2063.460 3416.280 ;
        RECT 2063.200 3415.340 2063.460 3415.600 ;
        RECT 2065.500 3332.720 2065.760 3332.980 ;
        RECT 2064.120 3236.160 2064.380 3236.420 ;
        RECT 2064.580 3236.160 2064.840 3236.420 ;
        RECT 2064.120 3201.820 2064.380 3202.080 ;
        RECT 2064.580 3201.820 2064.840 3202.080 ;
        RECT 2063.660 3153.200 2063.920 3153.460 ;
        RECT 2064.580 3153.200 2064.840 3153.460 ;
        RECT 2063.660 3056.640 2063.920 3056.900 ;
        RECT 2064.580 3056.640 2064.840 3056.900 ;
        RECT 2064.120 3042.700 2064.380 3042.960 ;
        RECT 2065.040 3008.360 2065.300 3008.620 ;
        RECT 2065.040 2994.420 2065.300 2994.680 ;
        RECT 2065.500 2946.480 2065.760 2946.740 ;
        RECT 2065.500 2912.140 2065.760 2912.400 ;
        RECT 2065.040 2911.460 2065.300 2911.720 ;
        RECT 2063.660 2815.580 2063.920 2815.840 ;
        RECT 2063.660 2814.900 2063.920 2815.160 ;
        RECT 2063.660 2800.960 2063.920 2801.220 ;
        RECT 2064.580 2753.020 2064.840 2753.280 ;
        RECT 2063.660 2718.000 2063.920 2718.260 ;
        RECT 2064.580 2718.000 2064.840 2718.260 ;
        RECT 1809.280 2577.240 1809.540 2577.500 ;
        RECT 2064.580 2577.240 2064.840 2577.500 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2068.320 3517.230 2068.920 3517.370 ;
        RECT 2068.780 3491.450 2068.920 3517.230 ;
        RECT 2065.040 3491.130 2065.300 3491.450 ;
        RECT 2068.720 3491.130 2068.980 3491.450 ;
        RECT 2065.100 3470.710 2065.240 3491.130 ;
        RECT 2064.120 3470.390 2064.380 3470.710 ;
        RECT 2065.040 3470.390 2065.300 3470.710 ;
        RECT 2064.180 3463.910 2064.320 3470.390 ;
        RECT 2064.120 3463.590 2064.380 3463.910 ;
        RECT 2063.200 3415.990 2063.460 3416.310 ;
        RECT 2063.260 3415.630 2063.400 3415.990 ;
        RECT 2063.200 3415.310 2063.460 3415.630 ;
        RECT 2065.500 3332.690 2065.760 3333.010 ;
        RECT 2065.560 3298.410 2065.700 3332.690 ;
        RECT 2064.640 3298.270 2065.700 3298.410 ;
        RECT 2064.640 3236.450 2064.780 3298.270 ;
        RECT 2064.120 3236.130 2064.380 3236.450 ;
        RECT 2064.580 3236.130 2064.840 3236.450 ;
        RECT 2064.180 3202.110 2064.320 3236.130 ;
        RECT 2064.120 3201.790 2064.380 3202.110 ;
        RECT 2064.580 3201.790 2064.840 3202.110 ;
        RECT 2064.640 3153.490 2064.780 3201.790 ;
        RECT 2063.660 3153.170 2063.920 3153.490 ;
        RECT 2064.580 3153.170 2064.840 3153.490 ;
        RECT 2063.720 3152.890 2063.860 3153.170 ;
        RECT 2063.720 3152.750 2064.320 3152.890 ;
        RECT 2064.180 3105.290 2064.320 3152.750 ;
        RECT 2064.180 3105.150 2064.780 3105.290 ;
        RECT 2064.640 3056.930 2064.780 3105.150 ;
        RECT 2063.660 3056.610 2063.920 3056.930 ;
        RECT 2064.580 3056.610 2064.840 3056.930 ;
        RECT 2063.720 3056.330 2063.860 3056.610 ;
        RECT 2063.720 3056.190 2064.320 3056.330 ;
        RECT 2064.180 3042.990 2064.320 3056.190 ;
        RECT 2064.120 3042.670 2064.380 3042.990 ;
        RECT 2065.040 3008.330 2065.300 3008.650 ;
        RECT 2065.100 2994.710 2065.240 3008.330 ;
        RECT 2065.040 2994.390 2065.300 2994.710 ;
        RECT 2065.500 2946.450 2065.760 2946.770 ;
        RECT 2065.560 2912.430 2065.700 2946.450 ;
        RECT 2065.500 2912.110 2065.760 2912.430 ;
        RECT 2065.040 2911.430 2065.300 2911.750 ;
        RECT 2065.100 2863.210 2065.240 2911.430 ;
        RECT 2064.180 2863.070 2065.240 2863.210 ;
        RECT 2064.180 2849.610 2064.320 2863.070 ;
        RECT 2063.720 2849.470 2064.320 2849.610 ;
        RECT 2063.720 2815.870 2063.860 2849.470 ;
        RECT 2063.660 2815.550 2063.920 2815.870 ;
        RECT 2063.660 2814.870 2063.920 2815.190 ;
        RECT 2063.720 2801.250 2063.860 2814.870 ;
        RECT 2063.660 2800.930 2063.920 2801.250 ;
        RECT 2064.580 2752.990 2064.840 2753.310 ;
        RECT 2064.640 2718.290 2064.780 2752.990 ;
        RECT 2063.660 2717.970 2063.920 2718.290 ;
        RECT 2064.580 2717.970 2064.840 2718.290 ;
        RECT 2063.720 2670.090 2063.860 2717.970 ;
        RECT 2063.720 2669.950 2064.320 2670.090 ;
        RECT 2064.180 2622.490 2064.320 2669.950 ;
        RECT 2064.180 2622.350 2064.780 2622.490 ;
        RECT 2064.640 2577.530 2064.780 2622.350 ;
        RECT 1809.280 2577.210 1809.540 2577.530 ;
        RECT 2064.580 2577.210 2064.840 2577.530 ;
        RECT 1809.340 2562.185 1809.480 2577.210 ;
        RECT 1809.170 2561.900 1809.480 2562.185 ;
        RECT 1809.170 2558.185 1809.450 2561.900 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1738.945 2898.245 1739.115 2946.355 ;
        RECT 1739.405 2815.285 1739.575 2849.455 ;
      LAYER mcon ;
        RECT 1738.945 2946.185 1739.115 2946.355 ;
        RECT 1739.405 2849.285 1739.575 2849.455 ;
      LAYER met1 ;
        RECT 1738.870 3464.160 1739.190 3464.220 ;
        RECT 1744.390 3464.160 1744.710 3464.220 ;
        RECT 1738.870 3464.020 1744.710 3464.160 ;
        RECT 1738.870 3463.960 1739.190 3464.020 ;
        RECT 1744.390 3463.960 1744.710 3464.020 ;
        RECT 1738.870 3367.600 1739.190 3367.660 ;
        RECT 1739.790 3367.600 1740.110 3367.660 ;
        RECT 1738.870 3367.460 1740.110 3367.600 ;
        RECT 1738.870 3367.400 1739.190 3367.460 ;
        RECT 1739.790 3367.400 1740.110 3367.460 ;
        RECT 1738.870 3270.700 1739.190 3270.760 ;
        RECT 1739.790 3270.700 1740.110 3270.760 ;
        RECT 1738.870 3270.560 1740.110 3270.700 ;
        RECT 1738.870 3270.500 1739.190 3270.560 ;
        RECT 1739.790 3270.500 1740.110 3270.560 ;
        RECT 1738.870 3174.140 1739.190 3174.200 ;
        RECT 1739.790 3174.140 1740.110 3174.200 ;
        RECT 1738.870 3174.000 1740.110 3174.140 ;
        RECT 1738.870 3173.940 1739.190 3174.000 ;
        RECT 1739.790 3173.940 1740.110 3174.000 ;
        RECT 1738.870 3077.580 1739.190 3077.640 ;
        RECT 1739.790 3077.580 1740.110 3077.640 ;
        RECT 1738.870 3077.440 1740.110 3077.580 ;
        RECT 1738.870 3077.380 1739.190 3077.440 ;
        RECT 1739.790 3077.380 1740.110 3077.440 ;
        RECT 1738.870 2981.020 1739.190 2981.080 ;
        RECT 1739.790 2981.020 1740.110 2981.080 ;
        RECT 1738.870 2980.880 1740.110 2981.020 ;
        RECT 1738.870 2980.820 1739.190 2980.880 ;
        RECT 1739.790 2980.820 1740.110 2980.880 ;
        RECT 1738.885 2946.340 1739.175 2946.385 ;
        RECT 1739.330 2946.340 1739.650 2946.400 ;
        RECT 1738.885 2946.200 1739.650 2946.340 ;
        RECT 1738.885 2946.155 1739.175 2946.200 ;
        RECT 1739.330 2946.140 1739.650 2946.200 ;
        RECT 1738.870 2898.400 1739.190 2898.460 ;
        RECT 1738.870 2898.260 1739.385 2898.400 ;
        RECT 1738.870 2898.200 1739.190 2898.260 ;
        RECT 1739.330 2849.440 1739.650 2849.500 ;
        RECT 1739.135 2849.300 1739.650 2849.440 ;
        RECT 1739.330 2849.240 1739.650 2849.300 ;
        RECT 1739.345 2815.440 1739.635 2815.485 ;
        RECT 1740.250 2815.440 1740.570 2815.500 ;
        RECT 1739.345 2815.300 1740.570 2815.440 ;
        RECT 1739.345 2815.255 1739.635 2815.300 ;
        RECT 1740.250 2815.240 1740.570 2815.300 ;
        RECT 1739.330 2753.220 1739.650 2753.280 ;
        RECT 1740.710 2753.220 1741.030 2753.280 ;
        RECT 1739.330 2753.080 1741.030 2753.220 ;
        RECT 1739.330 2753.020 1739.650 2753.080 ;
        RECT 1740.710 2753.020 1741.030 2753.080 ;
        RECT 1740.710 2719.220 1741.030 2719.280 ;
        RECT 1740.340 2719.080 1741.030 2719.220 ;
        RECT 1740.340 2718.600 1740.480 2719.080 ;
        RECT 1740.710 2719.020 1741.030 2719.080 ;
        RECT 1740.250 2718.340 1740.570 2718.600 ;
        RECT 1739.330 2656.660 1739.650 2656.720 ;
        RECT 1740.710 2656.660 1741.030 2656.720 ;
        RECT 1739.330 2656.520 1741.030 2656.660 ;
        RECT 1739.330 2656.460 1739.650 2656.520 ;
        RECT 1740.710 2656.460 1741.030 2656.520 ;
        RECT 1739.790 2608.380 1740.110 2608.440 ;
        RECT 1740.710 2608.380 1741.030 2608.440 ;
        RECT 1739.790 2608.240 1741.030 2608.380 ;
        RECT 1739.790 2608.180 1740.110 2608.240 ;
        RECT 1740.710 2608.180 1741.030 2608.240 ;
        RECT 1632.610 2577.440 1632.930 2577.500 ;
        RECT 1739.790 2577.440 1740.110 2577.500 ;
        RECT 1632.610 2577.300 1740.110 2577.440 ;
        RECT 1632.610 2577.240 1632.930 2577.300 ;
        RECT 1739.790 2577.240 1740.110 2577.300 ;
      LAYER via ;
        RECT 1738.900 3463.960 1739.160 3464.220 ;
        RECT 1744.420 3463.960 1744.680 3464.220 ;
        RECT 1738.900 3367.400 1739.160 3367.660 ;
        RECT 1739.820 3367.400 1740.080 3367.660 ;
        RECT 1738.900 3270.500 1739.160 3270.760 ;
        RECT 1739.820 3270.500 1740.080 3270.760 ;
        RECT 1738.900 3173.940 1739.160 3174.200 ;
        RECT 1739.820 3173.940 1740.080 3174.200 ;
        RECT 1738.900 3077.380 1739.160 3077.640 ;
        RECT 1739.820 3077.380 1740.080 3077.640 ;
        RECT 1738.900 2980.820 1739.160 2981.080 ;
        RECT 1739.820 2980.820 1740.080 2981.080 ;
        RECT 1739.360 2946.140 1739.620 2946.400 ;
        RECT 1738.900 2898.200 1739.160 2898.460 ;
        RECT 1739.360 2849.240 1739.620 2849.500 ;
        RECT 1740.280 2815.240 1740.540 2815.500 ;
        RECT 1739.360 2753.020 1739.620 2753.280 ;
        RECT 1740.740 2753.020 1741.000 2753.280 ;
        RECT 1740.740 2719.020 1741.000 2719.280 ;
        RECT 1740.280 2718.340 1740.540 2718.600 ;
        RECT 1739.360 2656.460 1739.620 2656.720 ;
        RECT 1740.740 2656.460 1741.000 2656.720 ;
        RECT 1739.820 2608.180 1740.080 2608.440 ;
        RECT 1740.740 2608.180 1741.000 2608.440 ;
        RECT 1632.640 2577.240 1632.900 2577.500 ;
        RECT 1739.820 2577.240 1740.080 2577.500 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3517.370 1744.160 3517.600 ;
        RECT 1744.020 3517.230 1744.620 3517.370 ;
        RECT 1744.480 3464.250 1744.620 3517.230 ;
        RECT 1738.900 3463.930 1739.160 3464.250 ;
        RECT 1744.420 3463.930 1744.680 3464.250 ;
        RECT 1738.960 3415.370 1739.100 3463.930 ;
        RECT 1738.960 3415.230 1740.020 3415.370 ;
        RECT 1739.880 3367.690 1740.020 3415.230 ;
        RECT 1738.900 3367.370 1739.160 3367.690 ;
        RECT 1739.820 3367.370 1740.080 3367.690 ;
        RECT 1738.960 3318.810 1739.100 3367.370 ;
        RECT 1738.960 3318.670 1740.020 3318.810 ;
        RECT 1739.880 3270.790 1740.020 3318.670 ;
        RECT 1738.900 3270.470 1739.160 3270.790 ;
        RECT 1739.820 3270.470 1740.080 3270.790 ;
        RECT 1738.960 3222.250 1739.100 3270.470 ;
        RECT 1738.960 3222.110 1740.020 3222.250 ;
        RECT 1739.880 3174.230 1740.020 3222.110 ;
        RECT 1738.900 3173.910 1739.160 3174.230 ;
        RECT 1739.820 3173.910 1740.080 3174.230 ;
        RECT 1738.960 3125.690 1739.100 3173.910 ;
        RECT 1738.960 3125.550 1740.020 3125.690 ;
        RECT 1739.880 3077.670 1740.020 3125.550 ;
        RECT 1738.900 3077.350 1739.160 3077.670 ;
        RECT 1739.820 3077.350 1740.080 3077.670 ;
        RECT 1738.960 3029.130 1739.100 3077.350 ;
        RECT 1738.960 3028.990 1740.020 3029.130 ;
        RECT 1739.880 2981.110 1740.020 3028.990 ;
        RECT 1738.900 2980.850 1739.160 2981.110 ;
        RECT 1738.900 2980.790 1739.560 2980.850 ;
        RECT 1739.820 2980.790 1740.080 2981.110 ;
        RECT 1738.960 2980.710 1739.560 2980.790 ;
        RECT 1739.420 2980.170 1739.560 2980.710 ;
        RECT 1739.420 2980.030 1740.020 2980.170 ;
        RECT 1739.880 2959.770 1740.020 2980.030 ;
        RECT 1739.420 2959.630 1740.020 2959.770 ;
        RECT 1739.420 2946.430 1739.560 2959.630 ;
        RECT 1739.360 2946.110 1739.620 2946.430 ;
        RECT 1738.900 2898.170 1739.160 2898.490 ;
        RECT 1738.960 2863.210 1739.100 2898.170 ;
        RECT 1738.960 2863.070 1739.560 2863.210 ;
        RECT 1739.420 2849.530 1739.560 2863.070 ;
        RECT 1739.360 2849.210 1739.620 2849.530 ;
        RECT 1740.280 2815.210 1740.540 2815.530 ;
        RECT 1740.340 2801.445 1740.480 2815.210 ;
        RECT 1739.350 2801.075 1739.630 2801.445 ;
        RECT 1740.270 2801.075 1740.550 2801.445 ;
        RECT 1739.420 2753.310 1739.560 2801.075 ;
        RECT 1739.360 2752.990 1739.620 2753.310 ;
        RECT 1740.740 2752.990 1741.000 2753.310 ;
        RECT 1740.800 2719.310 1740.940 2752.990 ;
        RECT 1740.740 2718.990 1741.000 2719.310 ;
        RECT 1740.280 2718.310 1740.540 2718.630 ;
        RECT 1740.340 2704.885 1740.480 2718.310 ;
        RECT 1739.350 2704.515 1739.630 2704.885 ;
        RECT 1740.270 2704.515 1740.550 2704.885 ;
        RECT 1739.420 2656.750 1739.560 2704.515 ;
        RECT 1739.360 2656.430 1739.620 2656.750 ;
        RECT 1740.740 2656.430 1741.000 2656.750 ;
        RECT 1740.800 2608.470 1740.940 2656.430 ;
        RECT 1739.820 2608.150 1740.080 2608.470 ;
        RECT 1740.740 2608.150 1741.000 2608.470 ;
        RECT 1739.880 2577.530 1740.020 2608.150 ;
        RECT 1632.640 2577.210 1632.900 2577.530 ;
        RECT 1739.820 2577.210 1740.080 2577.530 ;
        RECT 1632.700 2562.185 1632.840 2577.210 ;
        RECT 1632.530 2561.900 1632.840 2562.185 ;
        RECT 1632.530 2558.185 1632.810 2561.900 ;
      LAYER via2 ;
        RECT 1739.350 2801.120 1739.630 2801.400 ;
        RECT 1740.270 2801.120 1740.550 2801.400 ;
        RECT 1739.350 2704.560 1739.630 2704.840 ;
        RECT 1740.270 2704.560 1740.550 2704.840 ;
      LAYER met3 ;
        RECT 1739.325 2801.410 1739.655 2801.425 ;
        RECT 1740.245 2801.410 1740.575 2801.425 ;
        RECT 1739.325 2801.110 1740.575 2801.410 ;
        RECT 1739.325 2801.095 1739.655 2801.110 ;
        RECT 1740.245 2801.095 1740.575 2801.110 ;
        RECT 1739.325 2704.850 1739.655 2704.865 ;
        RECT 1740.245 2704.850 1740.575 2704.865 ;
        RECT 1739.325 2704.550 1740.575 2704.850 ;
        RECT 1739.325 2704.535 1739.655 2704.550 ;
        RECT 1740.245 2704.535 1740.575 2704.550 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1420.165 3381.045 1420.335 3429.155 ;
        RECT 1420.165 2898.585 1420.335 2946.355 ;
        RECT 1420.165 2718.725 1420.335 2752.895 ;
      LAYER mcon ;
        RECT 1420.165 3428.985 1420.335 3429.155 ;
        RECT 1420.165 2946.185 1420.335 2946.355 ;
        RECT 1420.165 2752.725 1420.335 2752.895 ;
      LAYER met1 ;
        RECT 1419.170 3477.760 1419.490 3477.820 ;
        RECT 1419.630 3477.760 1419.950 3477.820 ;
        RECT 1419.170 3477.620 1419.950 3477.760 ;
        RECT 1419.170 3477.560 1419.490 3477.620 ;
        RECT 1419.630 3477.560 1419.950 3477.620 ;
        RECT 1419.630 3443.080 1419.950 3443.140 ;
        RECT 1420.550 3443.080 1420.870 3443.140 ;
        RECT 1419.630 3442.940 1420.870 3443.080 ;
        RECT 1419.630 3442.880 1419.950 3442.940 ;
        RECT 1420.550 3442.880 1420.870 3442.940 ;
        RECT 1420.105 3429.140 1420.395 3429.185 ;
        RECT 1420.550 3429.140 1420.870 3429.200 ;
        RECT 1420.105 3429.000 1420.870 3429.140 ;
        RECT 1420.105 3428.955 1420.395 3429.000 ;
        RECT 1420.550 3428.940 1420.870 3429.000 ;
        RECT 1420.090 3381.200 1420.410 3381.260 ;
        RECT 1419.895 3381.060 1420.410 3381.200 ;
        RECT 1420.090 3381.000 1420.410 3381.060 ;
        RECT 1420.090 3367.600 1420.410 3367.660 ;
        RECT 1421.010 3367.600 1421.330 3367.660 ;
        RECT 1420.090 3367.460 1421.330 3367.600 ;
        RECT 1420.090 3367.400 1420.410 3367.460 ;
        RECT 1421.010 3367.400 1421.330 3367.460 ;
        RECT 1420.090 3270.700 1420.410 3270.760 ;
        RECT 1421.010 3270.700 1421.330 3270.760 ;
        RECT 1420.090 3270.560 1421.330 3270.700 ;
        RECT 1420.090 3270.500 1420.410 3270.560 ;
        RECT 1421.010 3270.500 1421.330 3270.560 ;
        RECT 1420.090 3174.140 1420.410 3174.200 ;
        RECT 1421.010 3174.140 1421.330 3174.200 ;
        RECT 1420.090 3174.000 1421.330 3174.140 ;
        RECT 1420.090 3173.940 1420.410 3174.000 ;
        RECT 1421.010 3173.940 1421.330 3174.000 ;
        RECT 1420.090 3077.580 1420.410 3077.640 ;
        RECT 1421.010 3077.580 1421.330 3077.640 ;
        RECT 1420.090 3077.440 1421.330 3077.580 ;
        RECT 1420.090 3077.380 1420.410 3077.440 ;
        RECT 1421.010 3077.380 1421.330 3077.440 ;
        RECT 1420.090 2981.020 1420.410 2981.080 ;
        RECT 1421.010 2981.020 1421.330 2981.080 ;
        RECT 1420.090 2980.880 1421.330 2981.020 ;
        RECT 1420.090 2980.820 1420.410 2980.880 ;
        RECT 1421.010 2980.820 1421.330 2980.880 ;
        RECT 1420.090 2946.340 1420.410 2946.400 ;
        RECT 1419.895 2946.200 1420.410 2946.340 ;
        RECT 1420.090 2946.140 1420.410 2946.200 ;
        RECT 1420.090 2898.740 1420.410 2898.800 ;
        RECT 1419.895 2898.600 1420.410 2898.740 ;
        RECT 1420.090 2898.540 1420.410 2898.600 ;
        RECT 1419.630 2898.060 1419.950 2898.120 ;
        RECT 1420.550 2898.060 1420.870 2898.120 ;
        RECT 1419.630 2897.920 1420.870 2898.060 ;
        RECT 1419.630 2897.860 1419.950 2897.920 ;
        RECT 1420.550 2897.860 1420.870 2897.920 ;
        RECT 1419.630 2814.760 1419.950 2814.820 ;
        RECT 1420.550 2814.760 1420.870 2814.820 ;
        RECT 1419.630 2814.620 1420.870 2814.760 ;
        RECT 1419.630 2814.560 1419.950 2814.620 ;
        RECT 1420.550 2814.560 1420.870 2814.620 ;
        RECT 1420.090 2752.880 1420.410 2752.940 ;
        RECT 1419.895 2752.740 1420.410 2752.880 ;
        RECT 1420.090 2752.680 1420.410 2752.740 ;
        RECT 1420.105 2718.880 1420.395 2718.925 ;
        RECT 1421.010 2718.880 1421.330 2718.940 ;
        RECT 1420.105 2718.740 1421.330 2718.880 ;
        RECT 1420.105 2718.695 1420.395 2718.740 ;
        RECT 1421.010 2718.680 1421.330 2718.740 ;
        RECT 1420.550 2621.640 1420.870 2621.700 ;
        RECT 1421.470 2621.640 1421.790 2621.700 ;
        RECT 1420.550 2621.500 1421.790 2621.640 ;
        RECT 1420.550 2621.440 1420.870 2621.500 ;
        RECT 1421.470 2621.440 1421.790 2621.500 ;
        RECT 1420.550 2580.500 1420.870 2580.560 ;
        RECT 1455.510 2580.500 1455.830 2580.560 ;
        RECT 1420.550 2580.360 1455.830 2580.500 ;
        RECT 1420.550 2580.300 1420.870 2580.360 ;
        RECT 1455.510 2580.300 1455.830 2580.360 ;
      LAYER via ;
        RECT 1419.200 3477.560 1419.460 3477.820 ;
        RECT 1419.660 3477.560 1419.920 3477.820 ;
        RECT 1419.660 3442.880 1419.920 3443.140 ;
        RECT 1420.580 3442.880 1420.840 3443.140 ;
        RECT 1420.580 3428.940 1420.840 3429.200 ;
        RECT 1420.120 3381.000 1420.380 3381.260 ;
        RECT 1420.120 3367.400 1420.380 3367.660 ;
        RECT 1421.040 3367.400 1421.300 3367.660 ;
        RECT 1420.120 3270.500 1420.380 3270.760 ;
        RECT 1421.040 3270.500 1421.300 3270.760 ;
        RECT 1420.120 3173.940 1420.380 3174.200 ;
        RECT 1421.040 3173.940 1421.300 3174.200 ;
        RECT 1420.120 3077.380 1420.380 3077.640 ;
        RECT 1421.040 3077.380 1421.300 3077.640 ;
        RECT 1420.120 2980.820 1420.380 2981.080 ;
        RECT 1421.040 2980.820 1421.300 2981.080 ;
        RECT 1420.120 2946.140 1420.380 2946.400 ;
        RECT 1420.120 2898.540 1420.380 2898.800 ;
        RECT 1419.660 2897.860 1419.920 2898.120 ;
        RECT 1420.580 2897.860 1420.840 2898.120 ;
        RECT 1419.660 2814.560 1419.920 2814.820 ;
        RECT 1420.580 2814.560 1420.840 2814.820 ;
        RECT 1420.120 2752.680 1420.380 2752.940 ;
        RECT 1421.040 2718.680 1421.300 2718.940 ;
        RECT 1420.580 2621.440 1420.840 2621.700 ;
        RECT 1421.500 2621.440 1421.760 2621.700 ;
        RECT 1420.580 2580.300 1420.840 2580.560 ;
        RECT 1455.540 2580.300 1455.800 2580.560 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3477.850 1419.400 3517.600 ;
        RECT 1419.200 3477.530 1419.460 3477.850 ;
        RECT 1419.660 3477.530 1419.920 3477.850 ;
        RECT 1419.720 3443.170 1419.860 3477.530 ;
        RECT 1419.660 3442.850 1419.920 3443.170 ;
        RECT 1420.580 3442.850 1420.840 3443.170 ;
        RECT 1420.640 3429.230 1420.780 3442.850 ;
        RECT 1420.580 3428.910 1420.840 3429.230 ;
        RECT 1420.120 3380.970 1420.380 3381.290 ;
        RECT 1420.180 3367.690 1420.320 3380.970 ;
        RECT 1420.120 3367.370 1420.380 3367.690 ;
        RECT 1421.040 3367.370 1421.300 3367.690 ;
        RECT 1421.100 3318.810 1421.240 3367.370 ;
        RECT 1420.180 3318.670 1421.240 3318.810 ;
        RECT 1420.180 3270.790 1420.320 3318.670 ;
        RECT 1420.120 3270.470 1420.380 3270.790 ;
        RECT 1421.040 3270.470 1421.300 3270.790 ;
        RECT 1421.100 3222.250 1421.240 3270.470 ;
        RECT 1420.180 3222.110 1421.240 3222.250 ;
        RECT 1420.180 3174.230 1420.320 3222.110 ;
        RECT 1420.120 3173.910 1420.380 3174.230 ;
        RECT 1421.040 3173.910 1421.300 3174.230 ;
        RECT 1421.100 3125.690 1421.240 3173.910 ;
        RECT 1420.180 3125.550 1421.240 3125.690 ;
        RECT 1420.180 3077.670 1420.320 3125.550 ;
        RECT 1420.120 3077.350 1420.380 3077.670 ;
        RECT 1421.040 3077.350 1421.300 3077.670 ;
        RECT 1421.100 3029.130 1421.240 3077.350 ;
        RECT 1420.180 3028.990 1421.240 3029.130 ;
        RECT 1420.180 2981.110 1420.320 3028.990 ;
        RECT 1420.120 2980.790 1420.380 2981.110 ;
        RECT 1421.040 2980.850 1421.300 2981.110 ;
        RECT 1420.640 2980.790 1421.300 2980.850 ;
        RECT 1420.640 2980.710 1421.240 2980.790 ;
        RECT 1420.640 2959.770 1420.780 2980.710 ;
        RECT 1420.180 2959.630 1420.780 2959.770 ;
        RECT 1420.180 2946.430 1420.320 2959.630 ;
        RECT 1420.120 2946.110 1420.380 2946.430 ;
        RECT 1420.120 2898.570 1420.380 2898.830 ;
        RECT 1419.720 2898.510 1420.380 2898.570 ;
        RECT 1419.720 2898.430 1420.320 2898.510 ;
        RECT 1419.720 2898.150 1419.860 2898.430 ;
        RECT 1419.660 2897.830 1419.920 2898.150 ;
        RECT 1420.580 2897.830 1420.840 2898.150 ;
        RECT 1420.640 2814.850 1420.780 2897.830 ;
        RECT 1419.660 2814.530 1419.920 2814.850 ;
        RECT 1420.580 2814.530 1420.840 2814.850 ;
        RECT 1419.720 2766.650 1419.860 2814.530 ;
        RECT 1419.720 2766.510 1420.320 2766.650 ;
        RECT 1420.180 2752.970 1420.320 2766.510 ;
        RECT 1420.120 2752.650 1420.380 2752.970 ;
        RECT 1421.040 2718.650 1421.300 2718.970 ;
        RECT 1421.100 2704.885 1421.240 2718.650 ;
        RECT 1421.030 2704.515 1421.310 2704.885 ;
        RECT 1421.950 2704.515 1422.230 2704.885 ;
        RECT 1422.020 2669.410 1422.160 2704.515 ;
        RECT 1420.640 2669.270 1422.160 2669.410 ;
        RECT 1420.640 2656.605 1420.780 2669.270 ;
        RECT 1420.570 2656.235 1420.850 2656.605 ;
        RECT 1421.490 2656.235 1421.770 2656.605 ;
        RECT 1421.560 2621.730 1421.700 2656.235 ;
        RECT 1420.580 2621.410 1420.840 2621.730 ;
        RECT 1421.500 2621.410 1421.760 2621.730 ;
        RECT 1420.640 2580.590 1420.780 2621.410 ;
        RECT 1420.580 2580.270 1420.840 2580.590 ;
        RECT 1455.540 2580.270 1455.800 2580.590 ;
        RECT 1455.600 2562.185 1455.740 2580.270 ;
        RECT 1455.430 2561.900 1455.740 2562.185 ;
        RECT 1455.430 2558.185 1455.710 2561.900 ;
      LAYER via2 ;
        RECT 1421.030 2704.560 1421.310 2704.840 ;
        RECT 1421.950 2704.560 1422.230 2704.840 ;
        RECT 1420.570 2656.280 1420.850 2656.560 ;
        RECT 1421.490 2656.280 1421.770 2656.560 ;
      LAYER met3 ;
        RECT 1421.005 2704.850 1421.335 2704.865 ;
        RECT 1421.925 2704.850 1422.255 2704.865 ;
        RECT 1421.005 2704.550 1422.255 2704.850 ;
        RECT 1421.005 2704.535 1421.335 2704.550 ;
        RECT 1421.925 2704.535 1422.255 2704.550 ;
        RECT 1420.545 2656.570 1420.875 2656.585 ;
        RECT 1421.465 2656.570 1421.795 2656.585 ;
        RECT 1420.545 2656.270 1421.795 2656.570 ;
        RECT 1420.545 2656.255 1420.875 2656.270 ;
        RECT 1421.465 2656.255 1421.795 2656.270 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 386.140 2267.270 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2266.950 386.000 2901.150 386.140 ;
        RECT 2266.950 385.940 2267.270 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2266.980 385.940 2267.240 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2266.970 1120.115 2267.250 1120.485 ;
        RECT 2267.040 386.230 2267.180 1120.115 ;
        RECT 2266.980 385.910 2267.240 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2266.970 1120.160 2267.250 1120.440 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2266.945 1120.450 2267.275 1120.465 ;
        RECT 2250.780 1120.440 2267.275 1120.450 ;
        RECT 2247.465 1120.150 2267.275 1120.440 ;
        RECT 2247.465 1119.840 2251.465 1120.150 ;
        RECT 2266.945 1120.135 2267.275 1120.150 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1096.785 3084.225 1096.955 3132.675 ;
        RECT 1095.405 3043.425 1095.575 3057.195 ;
        RECT 1096.325 3007.725 1096.495 3042.915 ;
        RECT 1095.865 2946.525 1096.035 2994.635 ;
        RECT 1094.485 2849.625 1094.655 2898.075 ;
        RECT 1094.945 2753.065 1095.115 2801.175 ;
        RECT 1095.405 2608.225 1095.575 2622.335 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1096.785 3132.505 1096.955 3132.675 ;
        RECT 1095.405 3057.025 1095.575 3057.195 ;
        RECT 1096.325 3042.745 1096.495 3042.915 ;
        RECT 1095.865 2994.465 1096.035 2994.635 ;
        RECT 1094.485 2897.905 1094.655 2898.075 ;
        RECT 1094.945 2801.005 1095.115 2801.175 ;
        RECT 1095.405 2622.165 1095.575 2622.335 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.790 3187.740 1096.110 3187.800 ;
        RECT 1095.330 3187.600 1096.110 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.790 3187.540 1096.110 3187.600 ;
        RECT 1096.710 3132.660 1097.030 3132.720 ;
        RECT 1096.515 3132.520 1097.030 3132.660 ;
        RECT 1096.710 3132.460 1097.030 3132.520 ;
        RECT 1096.710 3084.380 1097.030 3084.440 ;
        RECT 1096.515 3084.240 1097.030 3084.380 ;
        RECT 1096.710 3084.180 1097.030 3084.240 ;
        RECT 1095.345 3057.180 1095.635 3057.225 ;
        RECT 1096.710 3057.180 1097.030 3057.240 ;
        RECT 1095.345 3057.040 1097.030 3057.180 ;
        RECT 1095.345 3056.995 1095.635 3057.040 ;
        RECT 1096.710 3056.980 1097.030 3057.040 ;
        RECT 1095.330 3043.580 1095.650 3043.640 ;
        RECT 1095.135 3043.440 1095.650 3043.580 ;
        RECT 1095.330 3043.380 1095.650 3043.440 ;
        RECT 1095.330 3042.900 1095.650 3042.960 ;
        RECT 1096.265 3042.900 1096.555 3042.945 ;
        RECT 1095.330 3042.760 1096.555 3042.900 ;
        RECT 1095.330 3042.700 1095.650 3042.760 ;
        RECT 1096.265 3042.715 1096.555 3042.760 ;
        RECT 1096.250 3007.880 1096.570 3007.940 ;
        RECT 1096.055 3007.740 1096.570 3007.880 ;
        RECT 1096.250 3007.680 1096.570 3007.740 ;
        RECT 1095.805 2994.620 1096.095 2994.665 ;
        RECT 1096.250 2994.620 1096.570 2994.680 ;
        RECT 1095.805 2994.480 1096.570 2994.620 ;
        RECT 1095.805 2994.435 1096.095 2994.480 ;
        RECT 1096.250 2994.420 1096.570 2994.480 ;
        RECT 1095.790 2946.680 1096.110 2946.740 ;
        RECT 1095.595 2946.540 1096.110 2946.680 ;
        RECT 1095.790 2946.480 1096.110 2946.540 ;
        RECT 1094.870 2912.000 1095.190 2912.060 ;
        RECT 1095.790 2912.000 1096.110 2912.060 ;
        RECT 1094.870 2911.860 1096.110 2912.000 ;
        RECT 1094.870 2911.800 1095.190 2911.860 ;
        RECT 1095.790 2911.800 1096.110 2911.860 ;
        RECT 1094.425 2898.060 1094.715 2898.105 ;
        RECT 1094.870 2898.060 1095.190 2898.120 ;
        RECT 1094.425 2897.920 1095.190 2898.060 ;
        RECT 1094.425 2897.875 1094.715 2897.920 ;
        RECT 1094.870 2897.860 1095.190 2897.920 ;
        RECT 1094.410 2849.780 1094.730 2849.840 ;
        RECT 1094.215 2849.640 1094.730 2849.780 ;
        RECT 1094.410 2849.580 1094.730 2849.640 ;
        RECT 1094.410 2815.240 1094.730 2815.500 ;
        RECT 1094.500 2814.760 1094.640 2815.240 ;
        RECT 1094.870 2814.760 1095.190 2814.820 ;
        RECT 1094.500 2814.620 1095.190 2814.760 ;
        RECT 1094.870 2814.560 1095.190 2814.620 ;
        RECT 1094.870 2801.160 1095.190 2801.220 ;
        RECT 1094.675 2801.020 1095.190 2801.160 ;
        RECT 1094.870 2800.960 1095.190 2801.020 ;
        RECT 1094.885 2753.220 1095.175 2753.265 ;
        RECT 1095.790 2753.220 1096.110 2753.280 ;
        RECT 1094.885 2753.080 1096.110 2753.220 ;
        RECT 1094.885 2753.035 1095.175 2753.080 ;
        RECT 1095.790 2753.020 1096.110 2753.080 ;
        RECT 1094.870 2718.200 1095.190 2718.260 ;
        RECT 1095.790 2718.200 1096.110 2718.260 ;
        RECT 1094.870 2718.060 1096.110 2718.200 ;
        RECT 1094.870 2718.000 1095.190 2718.060 ;
        RECT 1095.790 2718.000 1096.110 2718.060 ;
        RECT 1094.870 2670.260 1095.190 2670.320 ;
        RECT 1095.790 2670.260 1096.110 2670.320 ;
        RECT 1094.870 2670.120 1096.110 2670.260 ;
        RECT 1094.870 2670.060 1095.190 2670.120 ;
        RECT 1095.790 2670.060 1096.110 2670.120 ;
        RECT 1095.330 2622.320 1095.650 2622.380 ;
        RECT 1095.135 2622.180 1095.650 2622.320 ;
        RECT 1095.330 2622.120 1095.650 2622.180 ;
        RECT 1095.330 2608.380 1095.650 2608.440 ;
        RECT 1095.135 2608.240 1095.650 2608.380 ;
        RECT 1095.330 2608.180 1095.650 2608.240 ;
        RECT 1095.330 2577.100 1095.650 2577.160 ;
        RECT 1278.870 2577.100 1279.190 2577.160 ;
        RECT 1095.330 2576.960 1279.190 2577.100 ;
        RECT 1095.330 2576.900 1095.650 2576.960 ;
        RECT 1278.870 2576.900 1279.190 2576.960 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1095.820 3187.540 1096.080 3187.800 ;
        RECT 1096.740 3132.460 1097.000 3132.720 ;
        RECT 1096.740 3084.180 1097.000 3084.440 ;
        RECT 1096.740 3056.980 1097.000 3057.240 ;
        RECT 1095.360 3043.380 1095.620 3043.640 ;
        RECT 1095.360 3042.700 1095.620 3042.960 ;
        RECT 1096.280 3007.680 1096.540 3007.940 ;
        RECT 1096.280 2994.420 1096.540 2994.680 ;
        RECT 1095.820 2946.480 1096.080 2946.740 ;
        RECT 1094.900 2911.800 1095.160 2912.060 ;
        RECT 1095.820 2911.800 1096.080 2912.060 ;
        RECT 1094.900 2897.860 1095.160 2898.120 ;
        RECT 1094.440 2849.580 1094.700 2849.840 ;
        RECT 1094.440 2815.240 1094.700 2815.500 ;
        RECT 1094.900 2814.560 1095.160 2814.820 ;
        RECT 1094.900 2800.960 1095.160 2801.220 ;
        RECT 1095.820 2753.020 1096.080 2753.280 ;
        RECT 1094.900 2718.000 1095.160 2718.260 ;
        RECT 1095.820 2718.000 1096.080 2718.260 ;
        RECT 1094.900 2670.060 1095.160 2670.320 ;
        RECT 1095.820 2670.060 1096.080 2670.320 ;
        RECT 1095.360 2622.120 1095.620 2622.380 ;
        RECT 1095.360 2608.180 1095.620 2608.440 ;
        RECT 1095.360 2576.900 1095.620 2577.160 ;
        RECT 1278.900 2576.900 1279.160 2577.160 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1095.820 3187.510 1096.080 3187.830 ;
        RECT 1095.880 3152.890 1096.020 3187.510 ;
        RECT 1095.880 3152.750 1096.940 3152.890 ;
        RECT 1096.800 3132.750 1096.940 3152.750 ;
        RECT 1096.740 3132.430 1097.000 3132.750 ;
        RECT 1096.740 3084.150 1097.000 3084.470 ;
        RECT 1096.800 3057.270 1096.940 3084.150 ;
        RECT 1096.740 3056.950 1097.000 3057.270 ;
        RECT 1095.360 3043.350 1095.620 3043.670 ;
        RECT 1095.420 3042.990 1095.560 3043.350 ;
        RECT 1095.360 3042.670 1095.620 3042.990 ;
        RECT 1096.280 3007.650 1096.540 3007.970 ;
        RECT 1096.340 2994.710 1096.480 3007.650 ;
        RECT 1096.280 2994.390 1096.540 2994.710 ;
        RECT 1095.820 2946.450 1096.080 2946.770 ;
        RECT 1095.880 2912.090 1096.020 2946.450 ;
        RECT 1094.900 2911.770 1095.160 2912.090 ;
        RECT 1095.820 2911.770 1096.080 2912.090 ;
        RECT 1094.960 2898.150 1095.100 2911.770 ;
        RECT 1094.900 2897.830 1095.160 2898.150 ;
        RECT 1094.440 2849.550 1094.700 2849.870 ;
        RECT 1094.500 2815.530 1094.640 2849.550 ;
        RECT 1094.440 2815.210 1094.700 2815.530 ;
        RECT 1094.900 2814.530 1095.160 2814.850 ;
        RECT 1094.960 2801.250 1095.100 2814.530 ;
        RECT 1094.900 2800.930 1095.160 2801.250 ;
        RECT 1095.820 2752.990 1096.080 2753.310 ;
        RECT 1095.880 2718.290 1096.020 2752.990 ;
        RECT 1094.900 2717.970 1095.160 2718.290 ;
        RECT 1095.820 2717.970 1096.080 2718.290 ;
        RECT 1094.960 2670.350 1095.100 2717.970 ;
        RECT 1094.900 2670.030 1095.160 2670.350 ;
        RECT 1095.820 2670.030 1096.080 2670.350 ;
        RECT 1095.880 2656.490 1096.020 2670.030 ;
        RECT 1095.420 2656.350 1096.020 2656.490 ;
        RECT 1095.420 2622.410 1095.560 2656.350 ;
        RECT 1095.360 2622.090 1095.620 2622.410 ;
        RECT 1095.360 2608.150 1095.620 2608.470 ;
        RECT 1095.420 2577.190 1095.560 2608.150 ;
        RECT 1095.360 2576.870 1095.620 2577.190 ;
        RECT 1278.900 2576.870 1279.160 2577.190 ;
        RECT 1278.960 2562.185 1279.100 2576.870 ;
        RECT 1278.790 2561.900 1279.100 2562.185 ;
        RECT 1278.790 2558.185 1279.070 2561.900 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
        RECT 771.565 2898.585 771.735 2946.355 ;
        RECT 771.565 2718.725 771.735 2752.895 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
        RECT 771.565 2946.185 771.735 2946.355 ;
        RECT 771.565 2752.725 771.735 2752.895 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 2981.020 771.810 2981.080 ;
        RECT 772.410 2981.020 772.730 2981.080 ;
        RECT 771.490 2980.880 772.730 2981.020 ;
        RECT 771.490 2980.820 771.810 2980.880 ;
        RECT 772.410 2980.820 772.730 2980.880 ;
        RECT 771.490 2946.340 771.810 2946.400 ;
        RECT 771.295 2946.200 771.810 2946.340 ;
        RECT 771.490 2946.140 771.810 2946.200 ;
        RECT 771.490 2898.740 771.810 2898.800 ;
        RECT 771.295 2898.600 771.810 2898.740 ;
        RECT 771.490 2898.540 771.810 2898.600 ;
        RECT 771.030 2898.060 771.350 2898.120 ;
        RECT 771.950 2898.060 772.270 2898.120 ;
        RECT 771.030 2897.920 772.270 2898.060 ;
        RECT 771.030 2897.860 771.350 2897.920 ;
        RECT 771.950 2897.860 772.270 2897.920 ;
        RECT 771.030 2814.760 771.350 2814.820 ;
        RECT 771.950 2814.760 772.270 2814.820 ;
        RECT 771.030 2814.620 772.270 2814.760 ;
        RECT 771.030 2814.560 771.350 2814.620 ;
        RECT 771.950 2814.560 772.270 2814.620 ;
        RECT 771.490 2752.880 771.810 2752.940 ;
        RECT 771.295 2752.740 771.810 2752.880 ;
        RECT 771.490 2752.680 771.810 2752.740 ;
        RECT 771.505 2718.880 771.795 2718.925 ;
        RECT 772.410 2718.880 772.730 2718.940 ;
        RECT 771.505 2718.740 772.730 2718.880 ;
        RECT 771.505 2718.695 771.795 2718.740 ;
        RECT 772.410 2718.680 772.730 2718.740 ;
        RECT 771.030 2656.660 771.350 2656.720 ;
        RECT 771.490 2656.660 771.810 2656.720 ;
        RECT 771.030 2656.520 771.810 2656.660 ;
        RECT 771.030 2656.460 771.350 2656.520 ;
        RECT 771.490 2656.460 771.810 2656.520 ;
        RECT 771.490 2622.120 771.810 2622.380 ;
        RECT 771.580 2621.640 771.720 2622.120 ;
        RECT 771.950 2621.640 772.270 2621.700 ;
        RECT 771.580 2621.500 772.270 2621.640 ;
        RECT 771.950 2621.440 772.270 2621.500 ;
        RECT 771.950 2577.440 772.270 2577.500 ;
        RECT 1102.230 2577.440 1102.550 2577.500 ;
        RECT 771.950 2577.300 1102.550 2577.440 ;
        RECT 771.950 2577.240 772.270 2577.300 ;
        RECT 1102.230 2577.240 1102.550 2577.300 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 2980.820 771.780 2981.080 ;
        RECT 772.440 2980.820 772.700 2981.080 ;
        RECT 771.520 2946.140 771.780 2946.400 ;
        RECT 771.520 2898.540 771.780 2898.800 ;
        RECT 771.060 2897.860 771.320 2898.120 ;
        RECT 771.980 2897.860 772.240 2898.120 ;
        RECT 771.060 2814.560 771.320 2814.820 ;
        RECT 771.980 2814.560 772.240 2814.820 ;
        RECT 771.520 2752.680 771.780 2752.940 ;
        RECT 772.440 2718.680 772.700 2718.940 ;
        RECT 771.060 2656.460 771.320 2656.720 ;
        RECT 771.520 2656.460 771.780 2656.720 ;
        RECT 771.520 2622.120 771.780 2622.380 ;
        RECT 771.980 2621.440 772.240 2621.700 ;
        RECT 771.980 2577.240 772.240 2577.500 ;
        RECT 1102.260 2577.240 1102.520 2577.500 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 2981.110 771.720 3028.990 ;
        RECT 771.520 2980.790 771.780 2981.110 ;
        RECT 772.440 2980.850 772.700 2981.110 ;
        RECT 772.040 2980.790 772.700 2980.850 ;
        RECT 772.040 2980.710 772.640 2980.790 ;
        RECT 772.040 2959.770 772.180 2980.710 ;
        RECT 771.580 2959.630 772.180 2959.770 ;
        RECT 771.580 2946.430 771.720 2959.630 ;
        RECT 771.520 2946.110 771.780 2946.430 ;
        RECT 771.520 2898.570 771.780 2898.830 ;
        RECT 771.120 2898.510 771.780 2898.570 ;
        RECT 771.120 2898.430 771.720 2898.510 ;
        RECT 771.120 2898.150 771.260 2898.430 ;
        RECT 771.060 2897.830 771.320 2898.150 ;
        RECT 771.980 2897.830 772.240 2898.150 ;
        RECT 772.040 2814.850 772.180 2897.830 ;
        RECT 771.060 2814.530 771.320 2814.850 ;
        RECT 771.980 2814.530 772.240 2814.850 ;
        RECT 771.120 2766.650 771.260 2814.530 ;
        RECT 771.120 2766.510 771.720 2766.650 ;
        RECT 771.580 2752.970 771.720 2766.510 ;
        RECT 771.520 2752.650 771.780 2752.970 ;
        RECT 772.440 2718.650 772.700 2718.970 ;
        RECT 772.500 2704.885 772.640 2718.650 ;
        RECT 771.050 2704.515 771.330 2704.885 ;
        RECT 772.430 2704.515 772.710 2704.885 ;
        RECT 771.120 2656.750 771.260 2704.515 ;
        RECT 771.060 2656.430 771.320 2656.750 ;
        RECT 771.520 2656.430 771.780 2656.750 ;
        RECT 771.580 2622.410 771.720 2656.430 ;
        RECT 771.520 2622.090 771.780 2622.410 ;
        RECT 771.980 2621.410 772.240 2621.730 ;
        RECT 772.040 2577.530 772.180 2621.410 ;
        RECT 771.980 2577.210 772.240 2577.530 ;
        RECT 1102.260 2577.210 1102.520 2577.530 ;
        RECT 1102.320 2562.185 1102.460 2577.210 ;
        RECT 1102.150 2561.900 1102.460 2562.185 ;
        RECT 1102.150 2558.185 1102.430 2561.900 ;
      LAYER via2 ;
        RECT 771.050 2704.560 771.330 2704.840 ;
        RECT 772.430 2704.560 772.710 2704.840 ;
      LAYER met3 ;
        RECT 771.025 2704.850 771.355 2704.865 ;
        RECT 772.405 2704.850 772.735 2704.865 ;
        RECT 771.025 2704.550 772.735 2704.850 ;
        RECT 771.025 2704.535 771.355 2704.550 ;
        RECT 772.405 2704.535 772.735 2704.550 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2578.460 448.430 2578.520 ;
        RECT 925.130 2578.460 925.450 2578.520 ;
        RECT 448.110 2578.320 925.450 2578.460 ;
        RECT 448.110 2578.260 448.430 2578.320 ;
        RECT 925.130 2578.260 925.450 2578.320 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2578.260 448.400 2578.520 ;
        RECT 925.160 2578.260 925.420 2578.520 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2578.550 448.340 3498.270 ;
        RECT 448.140 2578.230 448.400 2578.550 ;
        RECT 925.160 2578.230 925.420 2578.550 ;
        RECT 925.220 2562.185 925.360 2578.230 ;
        RECT 925.050 2561.900 925.360 2562.185 ;
        RECT 925.050 2558.185 925.330 2561.900 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2577.440 124.130 2577.500 ;
        RECT 748.490 2577.440 748.810 2577.500 ;
        RECT 123.810 2577.300 748.810 2577.440 ;
        RECT 123.810 2577.240 124.130 2577.300 ;
        RECT 748.490 2577.240 748.810 2577.300 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2577.240 124.100 2577.500 ;
        RECT 748.520 2577.240 748.780 2577.500 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2577.530 124.040 3498.270 ;
        RECT 123.840 2577.210 124.100 2577.530 ;
        RECT 748.520 2577.210 748.780 2577.530 ;
        RECT 748.580 2562.185 748.720 2577.210 ;
        RECT 748.410 2561.900 748.720 2562.185 ;
        RECT 748.410 2558.185 748.690 2561.900 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2511.480 17.410 2511.540 ;
        RECT 641.770 2511.480 642.090 2511.540 ;
        RECT 17.090 2511.340 642.090 2511.480 ;
        RECT 17.090 2511.280 17.410 2511.340 ;
        RECT 641.770 2511.280 642.090 2511.340 ;
      LAYER via ;
        RECT 17.120 2511.280 17.380 2511.540 ;
        RECT 641.800 2511.280 642.060 2511.540 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 2511.570 17.320 3339.635 ;
        RECT 17.120 2511.250 17.380 2511.570 ;
        RECT 641.800 2511.250 642.060 2511.570 ;
        RECT 641.860 2504.965 642.000 2511.250 ;
        RECT 641.790 2504.595 642.070 2504.965 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 641.790 2504.640 642.070 2504.920 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 641.765 2504.930 642.095 2504.945 ;
        RECT 641.765 2504.920 660.100 2504.930 ;
        RECT 641.765 2504.630 664.000 2504.920 ;
        RECT 641.765 2504.615 642.095 2504.630 ;
        RECT 660.000 2504.320 664.000 2504.630 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2394.180 17.870 2394.240 ;
        RECT 641.770 2394.180 642.090 2394.240 ;
        RECT 17.550 2394.040 642.090 2394.180 ;
        RECT 17.550 2393.980 17.870 2394.040 ;
        RECT 641.770 2393.980 642.090 2394.040 ;
      LAYER via ;
        RECT 17.580 2393.980 17.840 2394.240 ;
        RECT 641.800 2393.980 642.060 2394.240 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 2394.270 17.780 3051.995 ;
        RECT 17.580 2393.950 17.840 2394.270 ;
        RECT 641.800 2393.950 642.060 2394.270 ;
        RECT 641.860 2390.725 642.000 2393.950 ;
        RECT 641.790 2390.355 642.070 2390.725 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 641.790 2390.400 642.070 2390.680 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 641.765 2390.690 642.095 2390.705 ;
        RECT 641.765 2390.680 660.100 2390.690 ;
        RECT 641.765 2390.390 664.000 2390.680 ;
        RECT 641.765 2390.375 642.095 2390.390 ;
        RECT 660.000 2390.080 664.000 2390.390 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 2276.880 18.330 2276.940 ;
        RECT 641.770 2276.880 642.090 2276.940 ;
        RECT 18.010 2276.740 642.090 2276.880 ;
        RECT 18.010 2276.680 18.330 2276.740 ;
        RECT 641.770 2276.680 642.090 2276.740 ;
      LAYER via ;
        RECT 18.040 2276.680 18.300 2276.940 ;
        RECT 641.800 2276.680 642.060 2276.940 ;
      LAYER met2 ;
        RECT 18.030 2765.035 18.310 2765.405 ;
        RECT 18.100 2276.970 18.240 2765.035 ;
        RECT 18.040 2276.650 18.300 2276.970 ;
        RECT 641.800 2276.650 642.060 2276.970 ;
        RECT 641.860 2276.485 642.000 2276.650 ;
        RECT 641.790 2276.115 642.070 2276.485 ;
      LAYER via2 ;
        RECT 18.030 2765.080 18.310 2765.360 ;
        RECT 641.790 2276.160 642.070 2276.440 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.005 2765.370 18.335 2765.385 ;
        RECT -4.800 2765.070 18.335 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.005 2765.055 18.335 2765.070 ;
        RECT 641.765 2276.450 642.095 2276.465 ;
        RECT 641.765 2276.440 660.100 2276.450 ;
        RECT 641.765 2276.150 664.000 2276.440 ;
        RECT 641.765 2276.135 642.095 2276.150 ;
        RECT 660.000 2275.840 664.000 2276.150 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2166.380 17.410 2166.440 ;
        RECT 641.770 2166.380 642.090 2166.440 ;
        RECT 17.090 2166.240 642.090 2166.380 ;
        RECT 17.090 2166.180 17.410 2166.240 ;
        RECT 641.770 2166.180 642.090 2166.240 ;
      LAYER via ;
        RECT 17.120 2166.180 17.380 2166.440 ;
        RECT 641.800 2166.180 642.060 2166.440 ;
      LAYER met2 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
        RECT 17.180 2166.470 17.320 2477.395 ;
        RECT 17.120 2166.150 17.380 2166.470 ;
        RECT 641.800 2166.150 642.060 2166.470 ;
        RECT 641.860 2161.565 642.000 2166.150 ;
        RECT 641.790 2161.195 642.070 2161.565 ;
      LAYER via2 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
        RECT 641.790 2161.240 642.070 2161.520 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
        RECT 641.765 2161.530 642.095 2161.545 ;
        RECT 641.765 2161.520 660.100 2161.530 ;
        RECT 641.765 2161.230 664.000 2161.520 ;
        RECT 641.765 2161.215 642.095 2161.230 ;
        RECT 660.000 2160.920 664.000 2161.230 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 2049.080 18.330 2049.140 ;
        RECT 641.770 2049.080 642.090 2049.140 ;
        RECT 18.010 2048.940 642.090 2049.080 ;
        RECT 18.010 2048.880 18.330 2048.940 ;
        RECT 641.770 2048.880 642.090 2048.940 ;
      LAYER via ;
        RECT 18.040 2048.880 18.300 2049.140 ;
        RECT 641.800 2048.880 642.060 2049.140 ;
      LAYER met2 ;
        RECT 18.030 2189.755 18.310 2190.125 ;
        RECT 18.100 2049.170 18.240 2189.755 ;
        RECT 18.040 2048.850 18.300 2049.170 ;
        RECT 641.800 2048.850 642.060 2049.170 ;
        RECT 641.860 2047.325 642.000 2048.850 ;
        RECT 641.790 2046.955 642.070 2047.325 ;
      LAYER via2 ;
        RECT 18.030 2189.800 18.310 2190.080 ;
        RECT 641.790 2047.000 642.070 2047.280 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.005 2190.090 18.335 2190.105 ;
        RECT -4.800 2189.790 18.335 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.005 2189.775 18.335 2189.790 ;
        RECT 641.765 2047.290 642.095 2047.305 ;
        RECT 641.765 2047.280 660.100 2047.290 ;
        RECT 641.765 2046.990 664.000 2047.280 ;
        RECT 641.765 2046.975 642.095 2046.990 ;
        RECT 660.000 2046.680 664.000 2046.990 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 644.990 1904.240 645.310 1904.300 ;
        RECT 16.170 1904.100 645.310 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 644.990 1904.040 645.310 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 645.020 1904.040 645.280 1904.300 ;
      LAYER met2 ;
        RECT 645.010 1932.715 645.290 1933.085 ;
        RECT 645.080 1904.330 645.220 1932.715 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 645.020 1904.010 645.280 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 645.010 1932.760 645.290 1933.040 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 644.985 1933.050 645.315 1933.065 ;
        RECT 644.985 1933.040 660.100 1933.050 ;
        RECT 644.985 1932.750 664.000 1933.040 ;
        RECT 644.985 1932.735 645.315 1932.750 ;
        RECT 660.000 1932.440 664.000 1932.750 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.410 620.740 2267.730 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2267.410 620.600 2901.150 620.740 ;
        RECT 2267.410 620.540 2267.730 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2267.440 620.540 2267.700 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2267.430 1226.875 2267.710 1227.245 ;
        RECT 2267.500 620.830 2267.640 1226.875 ;
        RECT 2267.440 620.510 2267.700 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2267.430 1226.920 2267.710 1227.200 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2267.405 1227.210 2267.735 1227.225 ;
        RECT 2250.780 1227.200 2267.735 1227.210 ;
        RECT 2247.465 1226.910 2267.735 1227.200 ;
        RECT 2247.465 1226.600 2251.465 1226.910 ;
        RECT 2267.405 1226.895 2267.735 1226.910 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1621.360 17.870 1621.420 ;
        RECT 644.990 1621.360 645.310 1621.420 ;
        RECT 17.550 1621.220 645.310 1621.360 ;
        RECT 17.550 1621.160 17.870 1621.220 ;
        RECT 644.990 1621.160 645.310 1621.220 ;
      LAYER via ;
        RECT 17.580 1621.160 17.840 1621.420 ;
        RECT 645.020 1621.160 645.280 1621.420 ;
      LAYER met2 ;
        RECT 645.010 1818.475 645.290 1818.845 ;
        RECT 645.080 1621.450 645.220 1818.475 ;
        RECT 17.580 1621.130 17.840 1621.450 ;
        RECT 645.020 1621.130 645.280 1621.450 ;
        RECT 17.640 1615.525 17.780 1621.130 ;
        RECT 17.570 1615.155 17.850 1615.525 ;
      LAYER via2 ;
        RECT 645.010 1818.520 645.290 1818.800 ;
        RECT 17.570 1615.200 17.850 1615.480 ;
      LAYER met3 ;
        RECT 644.985 1818.810 645.315 1818.825 ;
        RECT 644.985 1818.800 660.100 1818.810 ;
        RECT 644.985 1818.510 664.000 1818.800 ;
        RECT 644.985 1818.495 645.315 1818.510 ;
        RECT 660.000 1818.200 664.000 1818.510 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 17.545 1615.490 17.875 1615.505 ;
        RECT -4.800 1615.190 17.875 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 17.545 1615.175 17.875 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 645.450 1400.700 645.770 1400.760 ;
        RECT 17.090 1400.560 645.770 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 645.450 1400.500 645.770 1400.560 ;
      LAYER via ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 645.480 1400.500 645.740 1400.760 ;
      LAYER met2 ;
        RECT 645.470 1703.555 645.750 1703.925 ;
        RECT 645.540 1400.790 645.680 1703.555 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 645.480 1400.470 645.740 1400.790 ;
      LAYER via2 ;
        RECT 645.470 1703.600 645.750 1703.880 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 645.445 1703.890 645.775 1703.905 ;
        RECT 645.445 1703.880 660.100 1703.890 ;
        RECT 645.445 1703.590 664.000 1703.880 ;
        RECT 645.445 1703.575 645.775 1703.590 ;
        RECT 660.000 1703.280 664.000 1703.590 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1186.840 17.870 1186.900 ;
        RECT 644.990 1186.840 645.310 1186.900 ;
        RECT 17.550 1186.700 645.310 1186.840 ;
        RECT 17.550 1186.640 17.870 1186.700 ;
        RECT 644.990 1186.640 645.310 1186.700 ;
      LAYER via ;
        RECT 17.580 1186.640 17.840 1186.900 ;
        RECT 645.020 1186.640 645.280 1186.900 ;
      LAYER met2 ;
        RECT 645.010 1589.315 645.290 1589.685 ;
        RECT 645.080 1186.930 645.220 1589.315 ;
        RECT 17.580 1186.610 17.840 1186.930 ;
        RECT 645.020 1186.610 645.280 1186.930 ;
        RECT 17.640 1185.085 17.780 1186.610 ;
        RECT 17.570 1184.715 17.850 1185.085 ;
      LAYER via2 ;
        RECT 645.010 1589.360 645.290 1589.640 ;
        RECT 17.570 1184.760 17.850 1185.040 ;
      LAYER met3 ;
        RECT 644.985 1589.650 645.315 1589.665 ;
        RECT 644.985 1589.640 660.100 1589.650 ;
        RECT 644.985 1589.350 664.000 1589.640 ;
        RECT 644.985 1589.335 645.315 1589.350 ;
        RECT 660.000 1589.040 664.000 1589.350 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.545 1185.050 17.875 1185.065 ;
        RECT -4.800 1184.750 17.875 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.545 1184.735 17.875 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 972.640 14.650 972.700 ;
        RECT 646.830 972.640 647.150 972.700 ;
        RECT 14.330 972.500 647.150 972.640 ;
        RECT 14.330 972.440 14.650 972.500 ;
        RECT 646.830 972.440 647.150 972.500 ;
      LAYER via ;
        RECT 14.360 972.440 14.620 972.700 ;
        RECT 646.860 972.440 647.120 972.700 ;
      LAYER met2 ;
        RECT 646.850 1475.075 647.130 1475.445 ;
        RECT 646.920 972.730 647.060 1475.075 ;
        RECT 14.360 972.410 14.620 972.730 ;
        RECT 646.860 972.410 647.120 972.730 ;
        RECT 14.420 969.525 14.560 972.410 ;
        RECT 14.350 969.155 14.630 969.525 ;
      LAYER via2 ;
        RECT 646.850 1475.120 647.130 1475.400 ;
        RECT 14.350 969.200 14.630 969.480 ;
      LAYER met3 ;
        RECT 646.825 1475.410 647.155 1475.425 ;
        RECT 646.825 1475.400 660.100 1475.410 ;
        RECT 646.825 1475.110 664.000 1475.400 ;
        RECT 646.825 1475.095 647.155 1475.110 ;
        RECT 660.000 1474.800 664.000 1475.110 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 14.325 969.490 14.655 969.505 ;
        RECT -4.800 969.190 14.655 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 14.325 969.175 14.655 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 646.370 758.780 646.690 758.840 ;
        RECT 15.710 758.640 646.690 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 646.370 758.580 646.690 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 646.400 758.580 646.660 758.840 ;
      LAYER met2 ;
        RECT 646.390 1360.155 646.670 1360.525 ;
        RECT 646.460 758.870 646.600 1360.155 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 646.400 758.550 646.660 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 646.390 1360.200 646.670 1360.480 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 646.365 1360.490 646.695 1360.505 ;
        RECT 646.365 1360.480 660.100 1360.490 ;
        RECT 646.365 1360.190 664.000 1360.480 ;
        RECT 646.365 1360.175 646.695 1360.190 ;
        RECT 660.000 1359.880 664.000 1360.190 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 645.910 544.920 646.230 544.980 ;
        RECT 16.170 544.780 646.230 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 645.910 544.720 646.230 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 645.940 544.720 646.200 544.980 ;
      LAYER met2 ;
        RECT 645.930 1245.915 646.210 1246.285 ;
        RECT 646.000 545.010 646.140 1245.915 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 645.940 544.690 646.200 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 645.930 1245.960 646.210 1246.240 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 645.905 1246.250 646.235 1246.265 ;
        RECT 645.905 1246.240 660.100 1246.250 ;
        RECT 645.905 1245.950 664.000 1246.240 ;
        RECT 645.905 1245.935 646.235 1245.950 ;
        RECT 660.000 1245.640 664.000 1245.950 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 645.450 324.260 645.770 324.320 ;
        RECT 16.630 324.120 645.770 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 645.450 324.060 645.770 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 645.480 324.060 645.740 324.320 ;
      LAYER met2 ;
        RECT 645.470 1131.675 645.750 1132.045 ;
        RECT 645.540 324.350 645.680 1131.675 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 645.480 324.030 645.740 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 645.470 1131.720 645.750 1132.000 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 645.445 1132.010 645.775 1132.025 ;
        RECT 645.445 1132.000 660.100 1132.010 ;
        RECT 645.445 1131.710 664.000 1132.000 ;
        RECT 645.445 1131.695 645.775 1131.710 ;
        RECT 660.000 1131.400 664.000 1131.710 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 644.990 110.400 645.310 110.460 ;
        RECT 15.710 110.260 645.310 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 644.990 110.200 645.310 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 645.020 110.200 645.280 110.460 ;
      LAYER met2 ;
        RECT 645.010 1017.435 645.290 1017.805 ;
        RECT 645.080 110.490 645.220 1017.435 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 645.020 110.170 645.280 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 645.010 1017.480 645.290 1017.760 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 644.985 1017.770 645.315 1017.785 ;
        RECT 644.985 1017.760 660.100 1017.770 ;
        RECT 644.985 1017.470 664.000 1017.760 ;
        RECT 644.985 1017.455 645.315 1017.470 ;
        RECT 660.000 1017.160 664.000 1017.470 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.870 855.340 2268.190 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2267.870 855.200 2901.150 855.340 ;
        RECT 2267.870 855.140 2268.190 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2267.900 855.140 2268.160 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2267.890 1333.635 2268.170 1334.005 ;
        RECT 2267.960 855.430 2268.100 1333.635 ;
        RECT 2267.900 855.110 2268.160 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2267.890 1333.680 2268.170 1333.960 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2267.865 1333.970 2268.195 1333.985 ;
        RECT 2250.780 1333.960 2268.195 1333.970 ;
        RECT 2247.465 1333.670 2268.195 1333.960 ;
        RECT 2247.465 1333.360 2251.465 1333.670 ;
        RECT 2267.865 1333.655 2268.195 1333.670 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.490 1089.940 2266.810 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2266.490 1089.800 2901.150 1089.940 ;
        RECT 2266.490 1089.740 2266.810 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2266.520 1089.740 2266.780 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2266.510 1440.395 2266.790 1440.765 ;
        RECT 2266.580 1090.030 2266.720 1440.395 ;
        RECT 2266.520 1089.710 2266.780 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2266.510 1440.440 2266.790 1440.720 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2266.485 1440.730 2266.815 1440.745 ;
        RECT 2250.780 1440.720 2266.815 1440.730 ;
        RECT 2247.465 1440.430 2266.815 1440.720 ;
        RECT 2247.465 1440.120 2251.465 1440.430 ;
        RECT 2266.485 1440.415 2266.815 1440.430 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.410 1324.540 2267.730 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2267.410 1324.400 2901.150 1324.540 ;
        RECT 2267.410 1324.340 2267.730 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2267.440 1324.340 2267.700 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2267.430 1547.155 2267.710 1547.525 ;
        RECT 2267.500 1324.630 2267.640 1547.155 ;
        RECT 2267.440 1324.310 2267.700 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2267.430 1547.200 2267.710 1547.480 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2267.405 1547.490 2267.735 1547.505 ;
        RECT 2250.780 1547.480 2267.735 1547.490 ;
        RECT 2247.465 1547.190 2267.735 1547.480 ;
        RECT 2247.465 1546.880 2251.465 1547.190 ;
        RECT 2267.405 1547.175 2267.735 1547.190 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 1559.140 2267.270 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2266.950 1559.000 2901.150 1559.140 ;
        RECT 2266.950 1558.940 2267.270 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2266.980 1558.940 2267.240 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2266.970 1653.915 2267.250 1654.285 ;
        RECT 2267.040 1559.230 2267.180 1653.915 ;
        RECT 2266.980 1558.910 2267.240 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2266.970 1653.960 2267.250 1654.240 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2266.945 1654.250 2267.275 1654.265 ;
        RECT 2250.780 1654.240 2267.275 1654.250 ;
        RECT 2247.465 1653.950 2267.275 1654.240 ;
        RECT 2247.465 1653.640 2251.465 1653.950 ;
        RECT 2266.945 1653.935 2267.275 1653.950 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2268.790 1766.200 2269.110 1766.260 ;
        RECT 2901.290 1766.200 2901.610 1766.260 ;
        RECT 2268.790 1766.060 2901.610 1766.200 ;
        RECT 2268.790 1766.000 2269.110 1766.060 ;
        RECT 2901.290 1766.000 2901.610 1766.060 ;
      LAYER via ;
        RECT 2268.820 1766.000 2269.080 1766.260 ;
        RECT 2901.320 1766.000 2901.580 1766.260 ;
      LAYER met2 ;
        RECT 2901.310 1789.235 2901.590 1789.605 ;
        RECT 2901.380 1766.290 2901.520 1789.235 ;
        RECT 2268.820 1765.970 2269.080 1766.290 ;
        RECT 2901.320 1765.970 2901.580 1766.290 ;
        RECT 2268.880 1761.045 2269.020 1765.970 ;
        RECT 2268.810 1760.675 2269.090 1761.045 ;
      LAYER via2 ;
        RECT 2901.310 1789.280 2901.590 1789.560 ;
        RECT 2268.810 1760.720 2269.090 1761.000 ;
      LAYER met3 ;
        RECT 2901.285 1789.570 2901.615 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.285 1789.270 2924.800 1789.570 ;
        RECT 2901.285 1789.255 2901.615 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2268.785 1761.010 2269.115 1761.025 ;
        RECT 2250.780 1761.000 2269.115 1761.010 ;
        RECT 2247.465 1760.710 2269.115 1761.000 ;
        RECT 2247.465 1760.400 2251.465 1760.710 ;
        RECT 2268.785 1760.695 2269.115 1760.710 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 1869.900 2267.270 1869.960 ;
        RECT 2901.750 1869.900 2902.070 1869.960 ;
        RECT 2266.950 1869.760 2902.070 1869.900 ;
        RECT 2266.950 1869.700 2267.270 1869.760 ;
        RECT 2901.750 1869.700 2902.070 1869.760 ;
      LAYER via ;
        RECT 2266.980 1869.700 2267.240 1869.960 ;
        RECT 2901.780 1869.700 2902.040 1869.960 ;
      LAYER met2 ;
        RECT 2901.770 2023.835 2902.050 2024.205 ;
        RECT 2901.840 1869.990 2901.980 2023.835 ;
        RECT 2266.980 1869.670 2267.240 1869.990 ;
        RECT 2901.780 1869.670 2902.040 1869.990 ;
        RECT 2267.040 1867.805 2267.180 1869.670 ;
        RECT 2266.970 1867.435 2267.250 1867.805 ;
      LAYER via2 ;
        RECT 2901.770 2023.880 2902.050 2024.160 ;
        RECT 2266.970 1867.480 2267.250 1867.760 ;
      LAYER met3 ;
        RECT 2901.745 2024.170 2902.075 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.745 2023.870 2924.800 2024.170 ;
        RECT 2901.745 2023.855 2902.075 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2266.945 1867.770 2267.275 1867.785 ;
        RECT 2250.780 1867.760 2267.275 1867.770 ;
        RECT 2247.465 1867.470 2267.275 1867.760 ;
        RECT 2247.465 1867.160 2251.465 1867.470 ;
        RECT 2266.945 1867.455 2267.275 1867.470 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2268.790 1980.060 2269.110 1980.120 ;
        RECT 2901.290 1980.060 2901.610 1980.120 ;
        RECT 2268.790 1979.920 2901.610 1980.060 ;
        RECT 2268.790 1979.860 2269.110 1979.920 ;
        RECT 2901.290 1979.860 2901.610 1979.920 ;
      LAYER via ;
        RECT 2268.820 1979.860 2269.080 1980.120 ;
        RECT 2901.320 1979.860 2901.580 1980.120 ;
      LAYER met2 ;
        RECT 2901.310 2258.435 2901.590 2258.805 ;
        RECT 2901.380 1980.150 2901.520 2258.435 ;
        RECT 2268.820 1979.830 2269.080 1980.150 ;
        RECT 2901.320 1979.830 2901.580 1980.150 ;
        RECT 2268.880 1974.565 2269.020 1979.830 ;
        RECT 2268.810 1974.195 2269.090 1974.565 ;
      LAYER via2 ;
        RECT 2901.310 2258.480 2901.590 2258.760 ;
        RECT 2268.810 1974.240 2269.090 1974.520 ;
      LAYER met3 ;
        RECT 2901.285 2258.770 2901.615 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2901.285 2258.470 2924.800 2258.770 ;
        RECT 2901.285 2258.455 2901.615 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2268.785 1974.530 2269.115 1974.545 ;
        RECT 2250.780 1974.520 2269.115 1974.530 ;
        RECT 2247.465 1974.230 2269.115 1974.520 ;
        RECT 2247.465 1973.920 2251.465 1974.230 ;
        RECT 2268.785 1974.215 2269.115 1974.230 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 15.540 633.350 15.600 ;
        RECT 669.370 15.540 669.690 15.600 ;
        RECT 633.030 15.400 669.690 15.540 ;
        RECT 633.030 15.340 633.350 15.400 ;
        RECT 669.370 15.340 669.690 15.400 ;
      LAYER via ;
        RECT 633.060 15.340 633.320 15.600 ;
        RECT 669.400 15.340 669.660 15.600 ;
      LAYER met2 ;
        RECT 669.750 960.570 670.030 964.000 ;
        RECT 669.460 960.430 670.030 960.570 ;
        RECT 669.460 15.630 669.600 960.430 ;
        RECT 669.750 960.000 670.030 960.430 ;
        RECT 633.060 15.310 633.320 15.630 ;
        RECT 669.400 15.310 669.660 15.630 ;
        RECT 633.120 2.400 633.260 15.310 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1907.230 945.440 1907.550 945.500 ;
        RECT 1910.910 945.440 1911.230 945.500 ;
        RECT 1907.230 945.300 1911.230 945.440 ;
        RECT 1907.230 945.240 1907.550 945.300 ;
        RECT 1910.910 945.240 1911.230 945.300 ;
        RECT 1910.910 24.040 1911.230 24.100 ;
        RECT 2417.370 24.040 2417.690 24.100 ;
        RECT 1910.910 23.900 2417.690 24.040 ;
        RECT 1910.910 23.840 1911.230 23.900 ;
        RECT 2417.370 23.840 2417.690 23.900 ;
      LAYER via ;
        RECT 1907.260 945.240 1907.520 945.500 ;
        RECT 1910.940 945.240 1911.200 945.500 ;
        RECT 1910.940 23.840 1911.200 24.100 ;
        RECT 2417.400 23.840 2417.660 24.100 ;
      LAYER met2 ;
        RECT 1907.150 960.500 1907.430 964.000 ;
        RECT 1907.150 960.000 1907.460 960.500 ;
        RECT 1907.320 945.530 1907.460 960.000 ;
        RECT 1907.260 945.210 1907.520 945.530 ;
        RECT 1910.940 945.210 1911.200 945.530 ;
        RECT 1911.000 24.130 1911.140 945.210 ;
        RECT 1910.940 23.810 1911.200 24.130 ;
        RECT 2417.400 23.810 2417.660 24.130 ;
        RECT 2417.460 2.400 2417.600 23.810 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1919.190 948.840 1919.510 948.900 ;
        RECT 2428.870 948.840 2429.190 948.900 ;
        RECT 1919.190 948.700 2429.190 948.840 ;
        RECT 1919.190 948.640 1919.510 948.700 ;
        RECT 2428.870 948.640 2429.190 948.700 ;
        RECT 2428.870 17.920 2429.190 17.980 ;
        RECT 2434.850 17.920 2435.170 17.980 ;
        RECT 2428.870 17.780 2435.170 17.920 ;
        RECT 2428.870 17.720 2429.190 17.780 ;
        RECT 2434.850 17.720 2435.170 17.780 ;
      LAYER via ;
        RECT 1919.220 948.640 1919.480 948.900 ;
        RECT 2428.900 948.640 2429.160 948.900 ;
        RECT 2428.900 17.720 2429.160 17.980 ;
        RECT 2434.880 17.720 2435.140 17.980 ;
      LAYER met2 ;
        RECT 1919.110 960.500 1919.390 964.000 ;
        RECT 1919.110 960.000 1919.420 960.500 ;
        RECT 1919.280 948.930 1919.420 960.000 ;
        RECT 1919.220 948.610 1919.480 948.930 ;
        RECT 2428.900 948.610 2429.160 948.930 ;
        RECT 2428.960 18.010 2429.100 948.610 ;
        RECT 2428.900 17.690 2429.160 18.010 ;
        RECT 2434.880 17.690 2435.140 18.010 ;
        RECT 2434.940 2.400 2435.080 17.690 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.610 30.840 1931.930 30.900 ;
        RECT 2452.790 30.840 2453.110 30.900 ;
        RECT 1931.610 30.700 2453.110 30.840 ;
        RECT 1931.610 30.640 1931.930 30.700 ;
        RECT 2452.790 30.640 2453.110 30.700 ;
      LAYER via ;
        RECT 1931.640 30.640 1931.900 30.900 ;
        RECT 2452.820 30.640 2453.080 30.900 ;
      LAYER met2 ;
        RECT 1931.530 960.500 1931.810 964.000 ;
        RECT 1931.530 960.000 1931.840 960.500 ;
        RECT 1931.700 30.930 1931.840 960.000 ;
        RECT 1931.640 30.610 1931.900 30.930 ;
        RECT 2452.820 30.610 2453.080 30.930 ;
        RECT 2452.880 2.400 2453.020 30.610 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.030 941.700 1944.350 941.760 ;
        RECT 2470.270 941.700 2470.590 941.760 ;
        RECT 1944.030 941.560 2470.590 941.700 ;
        RECT 1944.030 941.500 1944.350 941.560 ;
        RECT 2470.270 941.500 2470.590 941.560 ;
      LAYER via ;
        RECT 1944.060 941.500 1944.320 941.760 ;
        RECT 2470.300 941.500 2470.560 941.760 ;
      LAYER met2 ;
        RECT 1943.950 960.500 1944.230 964.000 ;
        RECT 1943.950 960.000 1944.260 960.500 ;
        RECT 1944.120 941.790 1944.260 960.000 ;
        RECT 1944.060 941.470 1944.320 941.790 ;
        RECT 2470.300 941.470 2470.560 941.790 ;
        RECT 2470.360 17.410 2470.500 941.470 ;
        RECT 2470.360 17.270 2470.960 17.410 ;
        RECT 2470.820 2.400 2470.960 17.270 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1959.210 58.720 1959.530 58.780 ;
        RECT 2484.070 58.720 2484.390 58.780 ;
        RECT 1959.210 58.580 2484.390 58.720 ;
        RECT 1959.210 58.520 1959.530 58.580 ;
        RECT 2484.070 58.520 2484.390 58.580 ;
      LAYER via ;
        RECT 1959.240 58.520 1959.500 58.780 ;
        RECT 2484.100 58.520 2484.360 58.780 ;
      LAYER met2 ;
        RECT 1956.370 960.570 1956.650 964.000 ;
        RECT 1956.370 960.430 1959.440 960.570 ;
        RECT 1956.370 960.000 1956.650 960.430 ;
        RECT 1959.300 58.810 1959.440 960.430 ;
        RECT 1959.240 58.490 1959.500 58.810 ;
        RECT 2484.100 58.490 2484.360 58.810 ;
        RECT 2484.160 17.410 2484.300 58.490 ;
        RECT 2484.160 17.270 2488.900 17.410 ;
        RECT 2488.760 2.400 2488.900 17.270 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1968.870 934.900 1969.190 934.960 ;
        RECT 2504.770 934.900 2505.090 934.960 ;
        RECT 1968.870 934.760 2505.090 934.900 ;
        RECT 1968.870 934.700 1969.190 934.760 ;
        RECT 2504.770 934.700 2505.090 934.760 ;
        RECT 2504.770 2.960 2505.090 3.020 ;
        RECT 2506.150 2.960 2506.470 3.020 ;
        RECT 2504.770 2.820 2506.470 2.960 ;
        RECT 2504.770 2.760 2505.090 2.820 ;
        RECT 2506.150 2.760 2506.470 2.820 ;
      LAYER via ;
        RECT 1968.900 934.700 1969.160 934.960 ;
        RECT 2504.800 934.700 2505.060 934.960 ;
        RECT 2504.800 2.760 2505.060 3.020 ;
        RECT 2506.180 2.760 2506.440 3.020 ;
      LAYER met2 ;
        RECT 1968.790 960.500 1969.070 964.000 ;
        RECT 1968.790 960.000 1969.100 960.500 ;
        RECT 1968.960 934.990 1969.100 960.000 ;
        RECT 1968.900 934.670 1969.160 934.990 ;
        RECT 2504.800 934.670 2505.060 934.990 ;
        RECT 2504.860 3.050 2505.000 934.670 ;
        RECT 2504.800 2.730 2505.060 3.050 ;
        RECT 2506.180 2.730 2506.440 3.050 ;
        RECT 2506.240 2.400 2506.380 2.730 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1981.290 928.100 1981.610 928.160 ;
        RECT 2518.570 928.100 2518.890 928.160 ;
        RECT 1981.290 927.960 2518.890 928.100 ;
        RECT 1981.290 927.900 1981.610 927.960 ;
        RECT 2518.570 927.900 2518.890 927.960 ;
        RECT 2518.570 2.960 2518.890 3.020 ;
        RECT 2524.090 2.960 2524.410 3.020 ;
        RECT 2518.570 2.820 2524.410 2.960 ;
        RECT 2518.570 2.760 2518.890 2.820 ;
        RECT 2524.090 2.760 2524.410 2.820 ;
      LAYER via ;
        RECT 1981.320 927.900 1981.580 928.160 ;
        RECT 2518.600 927.900 2518.860 928.160 ;
        RECT 2518.600 2.760 2518.860 3.020 ;
        RECT 2524.120 2.760 2524.380 3.020 ;
      LAYER met2 ;
        RECT 1981.210 960.500 1981.490 964.000 ;
        RECT 1981.210 960.000 1981.520 960.500 ;
        RECT 1981.380 928.190 1981.520 960.000 ;
        RECT 1981.320 927.870 1981.580 928.190 ;
        RECT 2518.600 927.870 2518.860 928.190 ;
        RECT 2518.660 3.050 2518.800 927.870 ;
        RECT 2518.600 2.730 2518.860 3.050 ;
        RECT 2524.120 2.730 2524.380 3.050 ;
        RECT 2524.180 2.400 2524.320 2.730 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 37.980 1994.030 38.040 ;
        RECT 2542.030 37.980 2542.350 38.040 ;
        RECT 1993.710 37.840 2542.350 37.980 ;
        RECT 1993.710 37.780 1994.030 37.840 ;
        RECT 2542.030 37.780 2542.350 37.840 ;
      LAYER via ;
        RECT 1993.740 37.780 1994.000 38.040 ;
        RECT 2542.060 37.780 2542.320 38.040 ;
      LAYER met2 ;
        RECT 1993.630 960.500 1993.910 964.000 ;
        RECT 1993.630 960.000 1993.940 960.500 ;
        RECT 1993.800 38.070 1993.940 960.000 ;
        RECT 1993.740 37.750 1994.000 38.070 ;
        RECT 2542.060 37.750 2542.320 38.070 ;
        RECT 2542.120 2.400 2542.260 37.750 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.130 920.960 2006.450 921.020 ;
        RECT 2559.970 920.960 2560.290 921.020 ;
        RECT 2006.130 920.820 2560.290 920.960 ;
        RECT 2006.130 920.760 2006.450 920.820 ;
        RECT 2559.970 920.760 2560.290 920.820 ;
      LAYER via ;
        RECT 2006.160 920.760 2006.420 921.020 ;
        RECT 2560.000 920.760 2560.260 921.020 ;
      LAYER met2 ;
        RECT 2006.050 960.500 2006.330 964.000 ;
        RECT 2006.050 960.000 2006.360 960.500 ;
        RECT 2006.220 921.050 2006.360 960.000 ;
        RECT 2006.160 920.730 2006.420 921.050 ;
        RECT 2560.000 920.730 2560.260 921.050 ;
        RECT 2560.060 2.400 2560.200 920.730 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 65.520 2021.630 65.580 ;
        RECT 2573.770 65.520 2574.090 65.580 ;
        RECT 2021.310 65.380 2574.090 65.520 ;
        RECT 2021.310 65.320 2021.630 65.380 ;
        RECT 2573.770 65.320 2574.090 65.380 ;
      LAYER via ;
        RECT 2021.340 65.320 2021.600 65.580 ;
        RECT 2573.800 65.320 2574.060 65.580 ;
      LAYER met2 ;
        RECT 2018.470 960.570 2018.750 964.000 ;
        RECT 2018.470 960.430 2021.540 960.570 ;
        RECT 2018.470 960.000 2018.750 960.430 ;
        RECT 2021.400 65.610 2021.540 960.430 ;
        RECT 2021.340 65.290 2021.600 65.610 ;
        RECT 2573.800 65.290 2574.060 65.610 ;
        RECT 2573.860 17.410 2574.000 65.290 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 949.180 793.890 949.240 ;
        RECT 799.550 949.180 799.870 949.240 ;
        RECT 793.570 949.040 799.870 949.180 ;
        RECT 793.570 948.980 793.890 949.040 ;
        RECT 799.550 948.980 799.870 949.040 ;
        RECT 799.550 20.300 799.870 20.360 ;
        RECT 811.510 20.300 811.830 20.360 ;
        RECT 799.550 20.160 811.830 20.300 ;
        RECT 799.550 20.100 799.870 20.160 ;
        RECT 811.510 20.100 811.830 20.160 ;
      LAYER via ;
        RECT 793.600 948.980 793.860 949.240 ;
        RECT 799.580 948.980 799.840 949.240 ;
        RECT 799.580 20.100 799.840 20.360 ;
        RECT 811.540 20.100 811.800 20.360 ;
      LAYER met2 ;
        RECT 793.490 960.500 793.770 964.000 ;
        RECT 793.490 960.000 793.800 960.500 ;
        RECT 793.660 949.270 793.800 960.000 ;
        RECT 793.600 948.950 793.860 949.270 ;
        RECT 799.580 948.950 799.840 949.270 ;
        RECT 799.640 20.390 799.780 948.950 ;
        RECT 799.580 20.070 799.840 20.390 ;
        RECT 811.540 20.070 811.800 20.390 ;
        RECT 811.600 2.400 811.740 20.070 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2030.510 914.160 2030.830 914.220 ;
        RECT 2594.470 914.160 2594.790 914.220 ;
        RECT 2030.510 914.020 2594.790 914.160 ;
        RECT 2030.510 913.960 2030.830 914.020 ;
        RECT 2594.470 913.960 2594.790 914.020 ;
      LAYER via ;
        RECT 2030.540 913.960 2030.800 914.220 ;
        RECT 2594.500 913.960 2594.760 914.220 ;
      LAYER met2 ;
        RECT 2030.430 960.500 2030.710 964.000 ;
        RECT 2030.430 960.000 2030.740 960.500 ;
        RECT 2030.600 914.250 2030.740 960.000 ;
        RECT 2030.540 913.930 2030.800 914.250 ;
        RECT 2594.500 913.930 2594.760 914.250 ;
        RECT 2594.560 17.410 2594.700 913.930 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.930 950.880 2043.250 950.940 ;
        RECT 2048.450 950.880 2048.770 950.940 ;
        RECT 2042.930 950.740 2048.770 950.880 ;
        RECT 2042.930 950.680 2043.250 950.740 ;
        RECT 2048.450 950.680 2048.770 950.740 ;
        RECT 2048.450 900.560 2048.770 900.620 ;
        RECT 2608.270 900.560 2608.590 900.620 ;
        RECT 2048.450 900.420 2608.590 900.560 ;
        RECT 2048.450 900.360 2048.770 900.420 ;
        RECT 2608.270 900.360 2608.590 900.420 ;
      LAYER via ;
        RECT 2042.960 950.680 2043.220 950.940 ;
        RECT 2048.480 950.680 2048.740 950.940 ;
        RECT 2048.480 900.360 2048.740 900.620 ;
        RECT 2608.300 900.360 2608.560 900.620 ;
      LAYER met2 ;
        RECT 2042.850 960.500 2043.130 964.000 ;
        RECT 2042.850 960.000 2043.160 960.500 ;
        RECT 2043.020 950.970 2043.160 960.000 ;
        RECT 2042.960 950.650 2043.220 950.970 ;
        RECT 2048.480 950.650 2048.740 950.970 ;
        RECT 2048.540 900.650 2048.680 950.650 ;
        RECT 2048.480 900.330 2048.740 900.650 ;
        RECT 2608.300 900.330 2608.560 900.650 ;
        RECT 2608.360 17.410 2608.500 900.330 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.350 949.180 2055.670 949.240 ;
        RECT 2259.590 949.180 2259.910 949.240 ;
        RECT 2055.350 949.040 2259.910 949.180 ;
        RECT 2055.350 948.980 2055.670 949.040 ;
        RECT 2259.590 948.980 2259.910 949.040 ;
        RECT 2259.590 44.780 2259.910 44.840 ;
        RECT 2631.270 44.780 2631.590 44.840 ;
        RECT 2259.590 44.640 2631.590 44.780 ;
        RECT 2259.590 44.580 2259.910 44.640 ;
        RECT 2631.270 44.580 2631.590 44.640 ;
      LAYER via ;
        RECT 2055.380 948.980 2055.640 949.240 ;
        RECT 2259.620 948.980 2259.880 949.240 ;
        RECT 2259.620 44.580 2259.880 44.840 ;
        RECT 2631.300 44.580 2631.560 44.840 ;
      LAYER met2 ;
        RECT 2055.270 960.500 2055.550 964.000 ;
        RECT 2055.270 960.000 2055.580 960.500 ;
        RECT 2055.440 949.270 2055.580 960.000 ;
        RECT 2055.380 948.950 2055.640 949.270 ;
        RECT 2259.620 948.950 2259.880 949.270 ;
        RECT 2259.680 44.870 2259.820 948.950 ;
        RECT 2259.620 44.550 2259.880 44.870 ;
        RECT 2631.300 44.550 2631.560 44.870 ;
        RECT 2631.360 2.400 2631.500 44.550 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.150 893.420 2069.470 893.480 ;
        RECT 2642.770 893.420 2643.090 893.480 ;
        RECT 2069.150 893.280 2643.090 893.420 ;
        RECT 2069.150 893.220 2069.470 893.280 ;
        RECT 2642.770 893.220 2643.090 893.280 ;
        RECT 2642.770 17.920 2643.090 17.980 ;
        RECT 2649.210 17.920 2649.530 17.980 ;
        RECT 2642.770 17.780 2649.530 17.920 ;
        RECT 2642.770 17.720 2643.090 17.780 ;
        RECT 2649.210 17.720 2649.530 17.780 ;
      LAYER via ;
        RECT 2069.180 893.220 2069.440 893.480 ;
        RECT 2642.800 893.220 2643.060 893.480 ;
        RECT 2642.800 17.720 2643.060 17.980 ;
        RECT 2649.240 17.720 2649.500 17.980 ;
      LAYER met2 ;
        RECT 2067.690 960.570 2067.970 964.000 ;
        RECT 2067.690 960.430 2069.380 960.570 ;
        RECT 2067.690 960.000 2067.970 960.430 ;
        RECT 2069.240 893.510 2069.380 960.430 ;
        RECT 2069.180 893.190 2069.440 893.510 ;
        RECT 2642.800 893.190 2643.060 893.510 ;
        RECT 2642.860 18.010 2643.000 893.190 ;
        RECT 2642.800 17.690 2643.060 18.010 ;
        RECT 2649.240 17.690 2649.500 18.010 ;
        RECT 2649.300 2.400 2649.440 17.690 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 99.860 2083.730 99.920 ;
        RECT 2663.470 99.860 2663.790 99.920 ;
        RECT 2083.410 99.720 2663.790 99.860 ;
        RECT 2083.410 99.660 2083.730 99.720 ;
        RECT 2663.470 99.660 2663.790 99.720 ;
      LAYER via ;
        RECT 2083.440 99.660 2083.700 99.920 ;
        RECT 2663.500 99.660 2663.760 99.920 ;
      LAYER met2 ;
        RECT 2080.110 960.570 2080.390 964.000 ;
        RECT 2080.110 960.430 2083.640 960.570 ;
        RECT 2080.110 960.000 2080.390 960.430 ;
        RECT 2083.500 99.950 2083.640 960.430 ;
        RECT 2083.440 99.630 2083.700 99.950 ;
        RECT 2663.500 99.630 2663.760 99.950 ;
        RECT 2663.560 17.410 2663.700 99.630 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2092.610 945.440 2092.930 945.500 ;
        RECT 2100.890 945.440 2101.210 945.500 ;
        RECT 2092.610 945.300 2101.210 945.440 ;
        RECT 2092.610 945.240 2092.930 945.300 ;
        RECT 2100.890 945.240 2101.210 945.300 ;
        RECT 2100.890 886.620 2101.210 886.680 ;
        RECT 2684.170 886.620 2684.490 886.680 ;
        RECT 2100.890 886.480 2684.490 886.620 ;
        RECT 2100.890 886.420 2101.210 886.480 ;
        RECT 2684.170 886.420 2684.490 886.480 ;
      LAYER via ;
        RECT 2092.640 945.240 2092.900 945.500 ;
        RECT 2100.920 945.240 2101.180 945.500 ;
        RECT 2100.920 886.420 2101.180 886.680 ;
        RECT 2684.200 886.420 2684.460 886.680 ;
      LAYER met2 ;
        RECT 2092.530 960.500 2092.810 964.000 ;
        RECT 2092.530 960.000 2092.840 960.500 ;
        RECT 2092.700 945.530 2092.840 960.000 ;
        RECT 2092.640 945.210 2092.900 945.530 ;
        RECT 2100.920 945.210 2101.180 945.530 ;
        RECT 2100.980 886.710 2101.120 945.210 ;
        RECT 2100.920 886.390 2101.180 886.710 ;
        RECT 2684.200 886.390 2684.460 886.710 ;
        RECT 2684.260 17.410 2684.400 886.390 ;
        RECT 2684.260 17.270 2684.860 17.410 ;
        RECT 2684.720 2.400 2684.860 17.270 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.030 945.440 2105.350 945.500 ;
        RECT 2110.550 945.440 2110.870 945.500 ;
        RECT 2105.030 945.300 2110.870 945.440 ;
        RECT 2105.030 945.240 2105.350 945.300 ;
        RECT 2110.550 945.240 2110.870 945.300 ;
        RECT 2110.550 879.820 2110.870 879.880 ;
        RECT 2697.970 879.820 2698.290 879.880 ;
        RECT 2110.550 879.680 2698.290 879.820 ;
        RECT 2110.550 879.620 2110.870 879.680 ;
        RECT 2697.970 879.620 2698.290 879.680 ;
      LAYER via ;
        RECT 2105.060 945.240 2105.320 945.500 ;
        RECT 2110.580 945.240 2110.840 945.500 ;
        RECT 2110.580 879.620 2110.840 879.880 ;
        RECT 2698.000 879.620 2698.260 879.880 ;
      LAYER met2 ;
        RECT 2104.950 960.500 2105.230 964.000 ;
        RECT 2104.950 960.000 2105.260 960.500 ;
        RECT 2105.120 945.530 2105.260 960.000 ;
        RECT 2105.060 945.210 2105.320 945.530 ;
        RECT 2110.580 945.210 2110.840 945.530 ;
        RECT 2110.640 879.910 2110.780 945.210 ;
        RECT 2110.580 879.590 2110.840 879.910 ;
        RECT 2698.000 879.590 2698.260 879.910 ;
        RECT 2698.060 17.410 2698.200 879.590 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 51.580 2118.230 51.640 ;
        RECT 2718.670 51.580 2718.990 51.640 ;
        RECT 2117.910 51.440 2718.990 51.580 ;
        RECT 2117.910 51.380 2118.230 51.440 ;
        RECT 2718.670 51.380 2718.990 51.440 ;
      LAYER via ;
        RECT 2117.940 51.380 2118.200 51.640 ;
        RECT 2718.700 51.380 2718.960 51.640 ;
      LAYER met2 ;
        RECT 2117.370 960.570 2117.650 964.000 ;
        RECT 2117.370 960.430 2118.140 960.570 ;
        RECT 2117.370 960.000 2117.650 960.430 ;
        RECT 2118.000 51.670 2118.140 960.430 ;
        RECT 2117.940 51.350 2118.200 51.670 ;
        RECT 2718.700 51.350 2718.960 51.670 ;
        RECT 2718.760 17.410 2718.900 51.350 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.250 872.680 2131.570 872.740 ;
        RECT 2732.470 872.680 2732.790 872.740 ;
        RECT 2131.250 872.540 2732.790 872.680 ;
        RECT 2131.250 872.480 2131.570 872.540 ;
        RECT 2732.470 872.480 2732.790 872.540 ;
        RECT 2732.470 17.920 2732.790 17.980 ;
        RECT 2738.450 17.920 2738.770 17.980 ;
        RECT 2732.470 17.780 2738.770 17.920 ;
        RECT 2732.470 17.720 2732.790 17.780 ;
        RECT 2738.450 17.720 2738.770 17.780 ;
      LAYER via ;
        RECT 2131.280 872.480 2131.540 872.740 ;
        RECT 2732.500 872.480 2732.760 872.740 ;
        RECT 2732.500 17.720 2732.760 17.980 ;
        RECT 2738.480 17.720 2738.740 17.980 ;
      LAYER met2 ;
        RECT 2129.790 960.570 2130.070 964.000 ;
        RECT 2129.790 960.430 2131.480 960.570 ;
        RECT 2129.790 960.000 2130.070 960.430 ;
        RECT 2131.340 872.770 2131.480 960.430 ;
        RECT 2131.280 872.450 2131.540 872.770 ;
        RECT 2732.500 872.450 2732.760 872.770 ;
        RECT 2732.560 18.010 2732.700 872.450 ;
        RECT 2732.500 17.690 2732.760 18.010 ;
        RECT 2738.480 17.690 2738.740 18.010 ;
        RECT 2738.540 2.400 2738.680 17.690 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.830 945.440 2142.150 945.500 ;
        RECT 2145.510 945.440 2145.830 945.500 ;
        RECT 2141.830 945.300 2145.830 945.440 ;
        RECT 2141.830 945.240 2142.150 945.300 ;
        RECT 2145.510 945.240 2145.830 945.300 ;
        RECT 2145.510 127.740 2145.830 127.800 ;
        RECT 2753.170 127.740 2753.490 127.800 ;
        RECT 2145.510 127.600 2753.490 127.740 ;
        RECT 2145.510 127.540 2145.830 127.600 ;
        RECT 2753.170 127.540 2753.490 127.600 ;
      LAYER via ;
        RECT 2141.860 945.240 2142.120 945.500 ;
        RECT 2145.540 945.240 2145.800 945.500 ;
        RECT 2145.540 127.540 2145.800 127.800 ;
        RECT 2753.200 127.540 2753.460 127.800 ;
      LAYER met2 ;
        RECT 2141.750 960.500 2142.030 964.000 ;
        RECT 2141.750 960.000 2142.060 960.500 ;
        RECT 2141.920 945.530 2142.060 960.000 ;
        RECT 2141.860 945.210 2142.120 945.530 ;
        RECT 2145.540 945.210 2145.800 945.530 ;
        RECT 2145.600 127.830 2145.740 945.210 ;
        RECT 2145.540 127.510 2145.800 127.830 ;
        RECT 2753.200 127.510 2753.460 127.830 ;
        RECT 2753.260 17.410 2753.400 127.510 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.450 17.240 806.770 17.300 ;
        RECT 829.450 17.240 829.770 17.300 ;
        RECT 806.450 17.100 829.770 17.240 ;
        RECT 806.450 17.040 806.770 17.100 ;
        RECT 829.450 17.040 829.770 17.100 ;
      LAYER via ;
        RECT 806.480 17.040 806.740 17.300 ;
        RECT 829.480 17.040 829.740 17.300 ;
      LAYER met2 ;
        RECT 805.910 960.570 806.190 964.000 ;
        RECT 805.910 960.430 806.680 960.570 ;
        RECT 805.910 960.000 806.190 960.430 ;
        RECT 806.540 17.330 806.680 960.430 ;
        RECT 806.480 17.010 806.740 17.330 ;
        RECT 829.480 17.010 829.740 17.330 ;
        RECT 829.540 2.400 829.680 17.010 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2154.250 945.440 2154.570 945.500 ;
        RECT 2158.850 945.440 2159.170 945.500 ;
        RECT 2154.250 945.300 2159.170 945.440 ;
        RECT 2154.250 945.240 2154.570 945.300 ;
        RECT 2158.850 945.240 2159.170 945.300 ;
        RECT 2158.850 865.880 2159.170 865.940 ;
        RECT 2773.870 865.880 2774.190 865.940 ;
        RECT 2158.850 865.740 2774.190 865.880 ;
        RECT 2158.850 865.680 2159.170 865.740 ;
        RECT 2773.870 865.680 2774.190 865.740 ;
      LAYER via ;
        RECT 2154.280 945.240 2154.540 945.500 ;
        RECT 2158.880 945.240 2159.140 945.500 ;
        RECT 2158.880 865.680 2159.140 865.940 ;
        RECT 2773.900 865.680 2774.160 865.940 ;
      LAYER met2 ;
        RECT 2154.170 960.500 2154.450 964.000 ;
        RECT 2154.170 960.000 2154.480 960.500 ;
        RECT 2154.340 945.530 2154.480 960.000 ;
        RECT 2154.280 945.210 2154.540 945.530 ;
        RECT 2158.880 945.210 2159.140 945.530 ;
        RECT 2158.940 865.970 2159.080 945.210 ;
        RECT 2158.880 865.650 2159.140 865.970 ;
        RECT 2773.900 865.650 2774.160 865.970 ;
        RECT 2773.960 2.400 2774.100 865.650 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.670 950.540 2166.990 950.600 ;
        RECT 2172.650 950.540 2172.970 950.600 ;
        RECT 2166.670 950.400 2172.970 950.540 ;
        RECT 2166.670 950.340 2166.990 950.400 ;
        RECT 2172.650 950.340 2172.970 950.400 ;
        RECT 2172.650 859.080 2172.970 859.140 ;
        RECT 2787.670 859.080 2787.990 859.140 ;
        RECT 2172.650 858.940 2787.990 859.080 ;
        RECT 2172.650 858.880 2172.970 858.940 ;
        RECT 2787.670 858.880 2787.990 858.940 ;
      LAYER via ;
        RECT 2166.700 950.340 2166.960 950.600 ;
        RECT 2172.680 950.340 2172.940 950.600 ;
        RECT 2172.680 858.880 2172.940 859.140 ;
        RECT 2787.700 858.880 2787.960 859.140 ;
      LAYER met2 ;
        RECT 2166.590 960.500 2166.870 964.000 ;
        RECT 2166.590 960.000 2166.900 960.500 ;
        RECT 2166.760 950.630 2166.900 960.000 ;
        RECT 2166.700 950.310 2166.960 950.630 ;
        RECT 2172.680 950.310 2172.940 950.630 ;
        RECT 2172.740 859.170 2172.880 950.310 ;
        RECT 2172.680 858.850 2172.940 859.170 ;
        RECT 2787.700 858.850 2787.960 859.170 ;
        RECT 2787.760 17.410 2787.900 858.850 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 72.320 2180.330 72.380 ;
        RECT 2808.370 72.320 2808.690 72.380 ;
        RECT 2180.010 72.180 2808.690 72.320 ;
        RECT 2180.010 72.120 2180.330 72.180 ;
        RECT 2808.370 72.120 2808.690 72.180 ;
      LAYER via ;
        RECT 2180.040 72.120 2180.300 72.380 ;
        RECT 2808.400 72.120 2808.660 72.380 ;
      LAYER met2 ;
        RECT 2179.010 960.570 2179.290 964.000 ;
        RECT 2179.010 960.430 2180.240 960.570 ;
        RECT 2179.010 960.000 2179.290 960.430 ;
        RECT 2180.100 72.410 2180.240 960.430 ;
        RECT 2180.040 72.090 2180.300 72.410 ;
        RECT 2808.400 72.090 2808.660 72.410 ;
        RECT 2808.460 17.410 2808.600 72.090 ;
        RECT 2808.460 17.270 2809.980 17.410 ;
        RECT 2809.840 2.400 2809.980 17.270 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2193.350 845.140 2193.670 845.200 ;
        RECT 2822.170 845.140 2822.490 845.200 ;
        RECT 2193.350 845.000 2822.490 845.140 ;
        RECT 2193.350 844.940 2193.670 845.000 ;
        RECT 2822.170 844.940 2822.490 845.000 ;
      LAYER via ;
        RECT 2193.380 844.940 2193.640 845.200 ;
        RECT 2822.200 844.940 2822.460 845.200 ;
      LAYER met2 ;
        RECT 2191.430 960.570 2191.710 964.000 ;
        RECT 2191.430 960.430 2193.580 960.570 ;
        RECT 2191.430 960.000 2191.710 960.430 ;
        RECT 2193.440 845.230 2193.580 960.430 ;
        RECT 2193.380 844.910 2193.640 845.230 ;
        RECT 2822.200 844.910 2822.460 845.230 ;
        RECT 2822.260 17.410 2822.400 844.910 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2207.610 155.280 2207.930 155.340 ;
        RECT 2842.870 155.280 2843.190 155.340 ;
        RECT 2207.610 155.140 2843.190 155.280 ;
        RECT 2207.610 155.080 2207.930 155.140 ;
        RECT 2842.870 155.080 2843.190 155.140 ;
      LAYER via ;
        RECT 2207.640 155.080 2207.900 155.340 ;
        RECT 2842.900 155.080 2843.160 155.340 ;
      LAYER met2 ;
        RECT 2203.850 960.570 2204.130 964.000 ;
        RECT 2203.850 960.430 2207.840 960.570 ;
        RECT 2203.850 960.000 2204.130 960.430 ;
        RECT 2207.700 155.370 2207.840 960.430 ;
        RECT 2207.640 155.050 2207.900 155.370 ;
        RECT 2842.900 155.050 2843.160 155.370 ;
        RECT 2842.960 6.530 2843.100 155.050 ;
        RECT 2842.960 6.390 2845.400 6.530 ;
        RECT 2845.260 2.400 2845.400 6.390 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2216.350 945.440 2216.670 945.500 ;
        RECT 2220.950 945.440 2221.270 945.500 ;
        RECT 2216.350 945.300 2221.270 945.440 ;
        RECT 2216.350 945.240 2216.670 945.300 ;
        RECT 2220.950 945.240 2221.270 945.300 ;
        RECT 2220.950 838.340 2221.270 838.400 ;
        RECT 2856.670 838.340 2856.990 838.400 ;
        RECT 2220.950 838.200 2856.990 838.340 ;
        RECT 2220.950 838.140 2221.270 838.200 ;
        RECT 2856.670 838.140 2856.990 838.200 ;
        RECT 2856.670 16.560 2856.990 16.620 ;
        RECT 2863.110 16.560 2863.430 16.620 ;
        RECT 2856.670 16.420 2863.430 16.560 ;
        RECT 2856.670 16.360 2856.990 16.420 ;
        RECT 2863.110 16.360 2863.430 16.420 ;
      LAYER via ;
        RECT 2216.380 945.240 2216.640 945.500 ;
        RECT 2220.980 945.240 2221.240 945.500 ;
        RECT 2220.980 838.140 2221.240 838.400 ;
        RECT 2856.700 838.140 2856.960 838.400 ;
        RECT 2856.700 16.360 2856.960 16.620 ;
        RECT 2863.140 16.360 2863.400 16.620 ;
      LAYER met2 ;
        RECT 2216.270 960.500 2216.550 964.000 ;
        RECT 2216.270 960.000 2216.580 960.500 ;
        RECT 2216.440 945.530 2216.580 960.000 ;
        RECT 2216.380 945.210 2216.640 945.530 ;
        RECT 2220.980 945.210 2221.240 945.530 ;
        RECT 2221.040 838.430 2221.180 945.210 ;
        RECT 2220.980 838.110 2221.240 838.430 ;
        RECT 2856.700 838.110 2856.960 838.430 ;
        RECT 2856.760 16.650 2856.900 838.110 ;
        RECT 2856.700 16.330 2856.960 16.650 ;
        RECT 2863.140 16.330 2863.400 16.650 ;
        RECT 2863.200 2.400 2863.340 16.330 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2228.770 949.860 2229.090 949.920 ;
        RECT 2234.750 949.860 2235.070 949.920 ;
        RECT 2228.770 949.720 2235.070 949.860 ;
        RECT 2228.770 949.660 2229.090 949.720 ;
        RECT 2234.750 949.660 2235.070 949.720 ;
        RECT 2234.750 831.540 2235.070 831.600 ;
        RECT 2877.370 831.540 2877.690 831.600 ;
        RECT 2234.750 831.400 2877.690 831.540 ;
        RECT 2234.750 831.340 2235.070 831.400 ;
        RECT 2877.370 831.340 2877.690 831.400 ;
      LAYER via ;
        RECT 2228.800 949.660 2229.060 949.920 ;
        RECT 2234.780 949.660 2235.040 949.920 ;
        RECT 2234.780 831.340 2235.040 831.600 ;
        RECT 2877.400 831.340 2877.660 831.600 ;
      LAYER met2 ;
        RECT 2228.690 960.500 2228.970 964.000 ;
        RECT 2228.690 960.000 2229.000 960.500 ;
        RECT 2228.860 949.950 2229.000 960.000 ;
        RECT 2228.800 949.630 2229.060 949.950 ;
        RECT 2234.780 949.630 2235.040 949.950 ;
        RECT 2234.840 831.630 2234.980 949.630 ;
        RECT 2234.780 831.310 2235.040 831.630 ;
        RECT 2877.400 831.310 2877.660 831.630 ;
        RECT 2877.460 17.410 2877.600 831.310 ;
        RECT 2877.460 17.270 2881.280 17.410 ;
        RECT 2881.140 2.400 2881.280 17.270 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2241.650 824.400 2241.970 824.460 ;
        RECT 2894.390 824.400 2894.710 824.460 ;
        RECT 2241.650 824.260 2894.710 824.400 ;
        RECT 2241.650 824.200 2241.970 824.260 ;
        RECT 2894.390 824.200 2894.710 824.260 ;
        RECT 2894.390 16.560 2894.710 16.620 ;
        RECT 2898.990 16.560 2899.310 16.620 ;
        RECT 2894.390 16.420 2899.310 16.560 ;
        RECT 2894.390 16.360 2894.710 16.420 ;
        RECT 2898.990 16.360 2899.310 16.420 ;
      LAYER via ;
        RECT 2241.680 824.200 2241.940 824.460 ;
        RECT 2894.420 824.200 2894.680 824.460 ;
        RECT 2894.420 16.360 2894.680 16.620 ;
        RECT 2899.020 16.360 2899.280 16.620 ;
      LAYER met2 ;
        RECT 2241.110 960.570 2241.390 964.000 ;
        RECT 2241.110 960.430 2241.880 960.570 ;
        RECT 2241.110 960.000 2241.390 960.430 ;
        RECT 2241.740 824.490 2241.880 960.430 ;
        RECT 2241.680 824.170 2241.940 824.490 ;
        RECT 2894.420 824.170 2894.680 824.490 ;
        RECT 2894.480 16.650 2894.620 824.170 ;
        RECT 2894.420 16.330 2894.680 16.650 ;
        RECT 2899.020 16.330 2899.280 16.650 ;
        RECT 2899.080 2.400 2899.220 16.330 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 820.710 15.880 821.030 15.940 ;
        RECT 846.930 15.880 847.250 15.940 ;
        RECT 820.710 15.740 847.250 15.880 ;
        RECT 820.710 15.680 821.030 15.740 ;
        RECT 846.930 15.680 847.250 15.740 ;
      LAYER via ;
        RECT 820.740 15.680 821.000 15.940 ;
        RECT 846.960 15.680 847.220 15.940 ;
      LAYER met2 ;
        RECT 818.330 960.570 818.610 964.000 ;
        RECT 818.330 960.430 820.940 960.570 ;
        RECT 818.330 960.000 818.610 960.430 ;
        RECT 820.800 15.970 820.940 960.430 ;
        RECT 820.740 15.650 821.000 15.970 ;
        RECT 846.960 15.650 847.220 15.970 ;
        RECT 847.020 2.400 847.160 15.650 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 830.830 945.440 831.150 945.500 ;
        RECT 834.510 945.440 834.830 945.500 ;
        RECT 830.830 945.300 834.830 945.440 ;
        RECT 830.830 945.240 831.150 945.300 ;
        RECT 834.510 945.240 834.830 945.300 ;
        RECT 834.510 20.640 834.830 20.700 ;
        RECT 864.870 20.640 865.190 20.700 ;
        RECT 834.510 20.500 865.190 20.640 ;
        RECT 834.510 20.440 834.830 20.500 ;
        RECT 864.870 20.440 865.190 20.500 ;
      LAYER via ;
        RECT 830.860 945.240 831.120 945.500 ;
        RECT 834.540 945.240 834.800 945.500 ;
        RECT 834.540 20.440 834.800 20.700 ;
        RECT 864.900 20.440 865.160 20.700 ;
      LAYER met2 ;
        RECT 830.750 960.500 831.030 964.000 ;
        RECT 830.750 960.000 831.060 960.500 ;
        RECT 830.920 945.530 831.060 960.000 ;
        RECT 830.860 945.210 831.120 945.530 ;
        RECT 834.540 945.210 834.800 945.530 ;
        RECT 834.600 20.730 834.740 945.210 ;
        RECT 834.540 20.410 834.800 20.730 ;
        RECT 864.900 20.410 865.160 20.730 ;
        RECT 864.960 2.400 865.100 20.410 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 843.250 951.560 843.570 951.620 ;
        RECT 847.850 951.560 848.170 951.620 ;
        RECT 843.250 951.420 848.170 951.560 ;
        RECT 843.250 951.360 843.570 951.420 ;
        RECT 847.850 951.360 848.170 951.420 ;
        RECT 847.850 19.620 848.170 19.680 ;
        RECT 882.350 19.620 882.670 19.680 ;
        RECT 847.850 19.480 882.670 19.620 ;
        RECT 847.850 19.420 848.170 19.480 ;
        RECT 882.350 19.420 882.670 19.480 ;
      LAYER via ;
        RECT 843.280 951.360 843.540 951.620 ;
        RECT 847.880 951.360 848.140 951.620 ;
        RECT 847.880 19.420 848.140 19.680 ;
        RECT 882.380 19.420 882.640 19.680 ;
      LAYER met2 ;
        RECT 843.170 960.500 843.450 964.000 ;
        RECT 843.170 960.000 843.480 960.500 ;
        RECT 843.340 951.650 843.480 960.000 ;
        RECT 843.280 951.330 843.540 951.650 ;
        RECT 847.880 951.330 848.140 951.650 ;
        RECT 847.940 19.710 848.080 951.330 ;
        RECT 847.880 19.390 848.140 19.710 ;
        RECT 882.380 19.450 882.640 19.710 ;
        RECT 882.380 19.390 883.040 19.450 ;
        RECT 882.440 19.310 883.040 19.390 ;
        RECT 882.900 2.400 883.040 19.310 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.670 945.440 855.990 945.500 ;
        RECT 862.110 945.440 862.430 945.500 ;
        RECT 855.670 945.300 862.430 945.440 ;
        RECT 855.670 945.240 855.990 945.300 ;
        RECT 862.110 945.240 862.430 945.300 ;
        RECT 862.110 14.860 862.430 14.920 ;
        RECT 900.750 14.860 901.070 14.920 ;
        RECT 862.110 14.720 901.070 14.860 ;
        RECT 862.110 14.660 862.430 14.720 ;
        RECT 900.750 14.660 901.070 14.720 ;
      LAYER via ;
        RECT 855.700 945.240 855.960 945.500 ;
        RECT 862.140 945.240 862.400 945.500 ;
        RECT 862.140 14.660 862.400 14.920 ;
        RECT 900.780 14.660 901.040 14.920 ;
      LAYER met2 ;
        RECT 855.590 960.500 855.870 964.000 ;
        RECT 855.590 960.000 855.900 960.500 ;
        RECT 855.760 945.530 855.900 960.000 ;
        RECT 855.700 945.210 855.960 945.530 ;
        RECT 862.140 945.210 862.400 945.530 ;
        RECT 862.200 14.950 862.340 945.210 ;
        RECT 862.140 14.630 862.400 14.950 ;
        RECT 900.780 14.630 901.040 14.950 ;
        RECT 900.840 2.400 900.980 14.630 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 868.550 24.040 868.870 24.100 ;
        RECT 918.690 24.040 919.010 24.100 ;
        RECT 868.550 23.900 919.010 24.040 ;
        RECT 868.550 23.840 868.870 23.900 ;
        RECT 918.690 23.840 919.010 23.900 ;
      LAYER via ;
        RECT 868.580 23.840 868.840 24.100 ;
        RECT 918.720 23.840 918.980 24.100 ;
      LAYER met2 ;
        RECT 868.010 960.570 868.290 964.000 ;
        RECT 868.010 960.430 868.780 960.570 ;
        RECT 868.010 960.000 868.290 960.430 ;
        RECT 868.640 24.130 868.780 960.430 ;
        RECT 868.580 23.810 868.840 24.130 ;
        RECT 918.720 23.810 918.980 24.130 ;
        RECT 918.780 2.400 918.920 23.810 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 30.840 882.670 30.900 ;
        RECT 936.170 30.840 936.490 30.900 ;
        RECT 882.350 30.700 936.490 30.840 ;
        RECT 882.350 30.640 882.670 30.700 ;
        RECT 936.170 30.640 936.490 30.700 ;
      LAYER via ;
        RECT 882.380 30.640 882.640 30.900 ;
        RECT 936.200 30.640 936.460 30.900 ;
      LAYER met2 ;
        RECT 880.430 960.570 880.710 964.000 ;
        RECT 880.430 960.430 882.580 960.570 ;
        RECT 880.430 960.000 880.710 960.430 ;
        RECT 882.440 30.930 882.580 960.430 ;
        RECT 882.380 30.610 882.640 30.930 ;
        RECT 936.200 30.610 936.460 30.930 ;
        RECT 936.260 2.400 936.400 30.610 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 892.470 949.180 892.790 949.240 ;
        RECT 941.690 949.180 942.010 949.240 ;
        RECT 892.470 949.040 942.010 949.180 ;
        RECT 892.470 948.980 892.790 949.040 ;
        RECT 941.690 948.980 942.010 949.040 ;
        RECT 941.690 24.380 942.010 24.440 ;
        RECT 954.110 24.380 954.430 24.440 ;
        RECT 941.690 24.240 954.430 24.380 ;
        RECT 941.690 24.180 942.010 24.240 ;
        RECT 954.110 24.180 954.430 24.240 ;
      LAYER via ;
        RECT 892.500 948.980 892.760 949.240 ;
        RECT 941.720 948.980 941.980 949.240 ;
        RECT 941.720 24.180 941.980 24.440 ;
        RECT 954.140 24.180 954.400 24.440 ;
      LAYER met2 ;
        RECT 892.390 960.500 892.670 964.000 ;
        RECT 892.390 960.000 892.700 960.500 ;
        RECT 892.560 949.270 892.700 960.000 ;
        RECT 892.500 948.950 892.760 949.270 ;
        RECT 941.720 948.950 941.980 949.270 ;
        RECT 941.780 24.470 941.920 948.950 ;
        RECT 941.720 24.150 941.980 24.470 ;
        RECT 954.140 24.150 954.400 24.470 ;
        RECT 954.200 2.400 954.340 24.150 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 904.890 948.840 905.210 948.900 ;
        RECT 962.390 948.840 962.710 948.900 ;
        RECT 904.890 948.700 962.710 948.840 ;
        RECT 904.890 948.640 905.210 948.700 ;
        RECT 962.390 948.640 962.710 948.700 ;
        RECT 962.390 20.980 962.710 21.040 ;
        RECT 972.050 20.980 972.370 21.040 ;
        RECT 962.390 20.840 972.370 20.980 ;
        RECT 962.390 20.780 962.710 20.840 ;
        RECT 972.050 20.780 972.370 20.840 ;
      LAYER via ;
        RECT 904.920 948.640 905.180 948.900 ;
        RECT 962.420 948.640 962.680 948.900 ;
        RECT 962.420 20.780 962.680 21.040 ;
        RECT 972.080 20.780 972.340 21.040 ;
      LAYER met2 ;
        RECT 904.810 960.500 905.090 964.000 ;
        RECT 904.810 960.000 905.120 960.500 ;
        RECT 904.980 948.930 905.120 960.000 ;
        RECT 904.920 948.610 905.180 948.930 ;
        RECT 962.420 948.610 962.680 948.930 ;
        RECT 962.480 21.070 962.620 948.610 ;
        RECT 962.420 20.750 962.680 21.070 ;
        RECT 972.080 20.750 972.340 21.070 ;
        RECT 972.140 2.400 972.280 20.750 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 676.805 737.885 676.975 772.735 ;
        RECT 677.725 657.305 677.895 717.655 ;
        RECT 678.185 530.825 678.355 613.955 ;
        RECT 678.185 448.205 678.355 524.195 ;
        RECT 678.645 386.325 678.815 427.635 ;
        RECT 677.265 289.425 677.435 304.215 ;
        RECT 677.725 58.565 677.895 137.955 ;
      LAYER mcon ;
        RECT 676.805 772.565 676.975 772.735 ;
        RECT 677.725 717.485 677.895 717.655 ;
        RECT 678.185 613.785 678.355 613.955 ;
        RECT 678.185 524.025 678.355 524.195 ;
        RECT 678.645 427.465 678.815 427.635 ;
        RECT 677.265 304.045 677.435 304.215 ;
        RECT 677.725 137.785 677.895 137.955 ;
      LAYER met1 ;
        RECT 677.650 917.560 677.970 917.620 ;
        RECT 678.110 917.560 678.430 917.620 ;
        RECT 677.650 917.420 678.430 917.560 ;
        RECT 677.650 917.360 677.970 917.420 ;
        RECT 678.110 917.360 678.430 917.420 ;
        RECT 676.730 772.720 677.050 772.780 ;
        RECT 676.535 772.580 677.050 772.720 ;
        RECT 676.730 772.520 677.050 772.580 ;
        RECT 676.745 738.040 677.035 738.085 ;
        RECT 677.190 738.040 677.510 738.100 ;
        RECT 676.745 737.900 677.510 738.040 ;
        RECT 676.745 737.855 677.035 737.900 ;
        RECT 677.190 737.840 677.510 737.900 ;
        RECT 677.190 717.640 677.510 717.700 ;
        RECT 677.665 717.640 677.955 717.685 ;
        RECT 677.190 717.500 677.955 717.640 ;
        RECT 677.190 717.440 677.510 717.500 ;
        RECT 677.665 717.455 677.955 717.500 ;
        RECT 677.665 657.460 677.955 657.505 ;
        RECT 678.110 657.460 678.430 657.520 ;
        RECT 677.665 657.320 678.430 657.460 ;
        RECT 677.665 657.275 677.955 657.320 ;
        RECT 678.110 657.260 678.430 657.320 ;
        RECT 678.110 620.740 678.430 620.800 ;
        RECT 679.030 620.740 679.350 620.800 ;
        RECT 678.110 620.600 679.350 620.740 ;
        RECT 678.110 620.540 678.430 620.600 ;
        RECT 679.030 620.540 679.350 620.600 ;
        RECT 678.125 613.940 678.415 613.985 ;
        RECT 679.030 613.940 679.350 614.000 ;
        RECT 678.125 613.800 679.350 613.940 ;
        RECT 678.125 613.755 678.415 613.800 ;
        RECT 679.030 613.740 679.350 613.800 ;
        RECT 678.110 530.980 678.430 531.040 ;
        RECT 677.915 530.840 678.430 530.980 ;
        RECT 678.110 530.780 678.430 530.840 ;
        RECT 678.110 524.180 678.430 524.240 ;
        RECT 677.915 524.040 678.430 524.180 ;
        RECT 678.110 523.980 678.430 524.040 ;
        RECT 677.650 448.360 677.970 448.420 ;
        RECT 678.125 448.360 678.415 448.405 ;
        RECT 677.650 448.220 678.415 448.360 ;
        RECT 677.650 448.160 677.970 448.220 ;
        RECT 678.125 448.175 678.415 448.220 ;
        RECT 677.190 434.760 677.510 434.820 ;
        RECT 678.570 434.760 678.890 434.820 ;
        RECT 677.190 434.620 678.890 434.760 ;
        RECT 677.190 434.560 677.510 434.620 ;
        RECT 678.570 434.560 678.890 434.620 ;
        RECT 678.570 427.620 678.890 427.680 ;
        RECT 678.375 427.480 678.890 427.620 ;
        RECT 678.570 427.420 678.890 427.480 ;
        RECT 678.570 386.480 678.890 386.540 ;
        RECT 678.375 386.340 678.890 386.480 ;
        RECT 678.570 386.280 678.890 386.340 ;
        RECT 677.190 331.400 677.510 331.460 ;
        RECT 678.570 331.400 678.890 331.460 ;
        RECT 677.190 331.260 678.890 331.400 ;
        RECT 677.190 331.200 677.510 331.260 ;
        RECT 678.570 331.200 678.890 331.260 ;
        RECT 677.190 304.200 677.510 304.260 ;
        RECT 676.995 304.060 677.510 304.200 ;
        RECT 677.190 304.000 677.510 304.060 ;
        RECT 677.190 289.580 677.510 289.640 ;
        RECT 676.995 289.440 677.510 289.580 ;
        RECT 677.190 289.380 677.510 289.440 ;
        RECT 677.190 137.940 677.510 138.000 ;
        RECT 677.665 137.940 677.955 137.985 ;
        RECT 677.190 137.800 677.955 137.940 ;
        RECT 677.190 137.740 677.510 137.800 ;
        RECT 677.665 137.755 677.955 137.800 ;
        RECT 677.650 58.720 677.970 58.780 ;
        RECT 677.455 58.580 677.970 58.720 ;
        RECT 677.650 58.520 677.970 58.580 ;
        RECT 650.970 20.300 651.290 20.360 ;
        RECT 677.650 20.300 677.970 20.360 ;
        RECT 650.970 20.160 677.970 20.300 ;
        RECT 650.970 20.100 651.290 20.160 ;
        RECT 677.650 20.100 677.970 20.160 ;
      LAYER via ;
        RECT 677.680 917.360 677.940 917.620 ;
        RECT 678.140 917.360 678.400 917.620 ;
        RECT 676.760 772.520 677.020 772.780 ;
        RECT 677.220 737.840 677.480 738.100 ;
        RECT 677.220 717.440 677.480 717.700 ;
        RECT 678.140 657.260 678.400 657.520 ;
        RECT 678.140 620.540 678.400 620.800 ;
        RECT 679.060 620.540 679.320 620.800 ;
        RECT 679.060 613.740 679.320 614.000 ;
        RECT 678.140 530.780 678.400 531.040 ;
        RECT 678.140 523.980 678.400 524.240 ;
        RECT 677.680 448.160 677.940 448.420 ;
        RECT 677.220 434.560 677.480 434.820 ;
        RECT 678.600 434.560 678.860 434.820 ;
        RECT 678.600 427.420 678.860 427.680 ;
        RECT 678.600 386.280 678.860 386.540 ;
        RECT 677.220 331.200 677.480 331.460 ;
        RECT 678.600 331.200 678.860 331.460 ;
        RECT 677.220 304.000 677.480 304.260 ;
        RECT 677.220 289.380 677.480 289.640 ;
        RECT 677.220 137.740 677.480 138.000 ;
        RECT 677.680 58.520 677.940 58.780 ;
        RECT 651.000 20.100 651.260 20.360 ;
        RECT 677.680 20.100 677.940 20.360 ;
      LAYER met2 ;
        RECT 682.170 961.250 682.450 964.000 ;
        RECT 678.660 961.110 682.450 961.250 ;
        RECT 678.660 946.290 678.800 961.110 ;
        RECT 682.170 960.000 682.450 961.110 ;
        RECT 678.200 946.150 678.800 946.290 ;
        RECT 678.200 931.330 678.340 946.150 ;
        RECT 677.740 931.190 678.340 931.330 ;
        RECT 677.740 917.650 677.880 931.190 ;
        RECT 677.680 917.330 677.940 917.650 ;
        RECT 678.140 917.330 678.400 917.650 ;
        RECT 678.200 834.770 678.340 917.330 ;
        RECT 677.280 834.630 678.340 834.770 ;
        RECT 677.280 796.690 677.420 834.630 ;
        RECT 676.820 796.550 677.420 796.690 ;
        RECT 676.820 772.810 676.960 796.550 ;
        RECT 676.760 772.490 677.020 772.810 ;
        RECT 677.220 737.810 677.480 738.130 ;
        RECT 677.280 717.730 677.420 737.810 ;
        RECT 677.220 717.410 677.480 717.730 ;
        RECT 678.140 657.230 678.400 657.550 ;
        RECT 678.200 620.830 678.340 657.230 ;
        RECT 678.140 620.510 678.400 620.830 ;
        RECT 679.060 620.510 679.320 620.830 ;
        RECT 679.120 614.030 679.260 620.510 ;
        RECT 679.060 613.710 679.320 614.030 ;
        RECT 678.140 530.750 678.400 531.070 ;
        RECT 678.200 524.270 678.340 530.750 ;
        RECT 678.140 523.950 678.400 524.270 ;
        RECT 677.680 448.130 677.940 448.450 ;
        RECT 677.740 434.930 677.880 448.130 ;
        RECT 677.280 434.850 677.880 434.930 ;
        RECT 677.220 434.790 677.880 434.850 ;
        RECT 677.220 434.530 677.480 434.790 ;
        RECT 678.600 434.530 678.860 434.850 ;
        RECT 678.660 427.710 678.800 434.530 ;
        RECT 678.600 427.390 678.860 427.710 ;
        RECT 678.600 386.250 678.860 386.570 ;
        RECT 678.660 331.490 678.800 386.250 ;
        RECT 677.220 331.170 677.480 331.490 ;
        RECT 678.600 331.170 678.860 331.490 ;
        RECT 677.280 304.290 677.420 331.170 ;
        RECT 677.220 303.970 677.480 304.290 ;
        RECT 677.220 289.350 677.480 289.670 ;
        RECT 677.280 217.330 677.420 289.350 ;
        RECT 677.280 217.190 677.880 217.330 ;
        RECT 677.740 158.170 677.880 217.190 ;
        RECT 677.280 158.030 677.880 158.170 ;
        RECT 677.280 138.030 677.420 158.030 ;
        RECT 677.220 137.710 677.480 138.030 ;
        RECT 677.680 58.490 677.940 58.810 ;
        RECT 677.740 20.390 677.880 58.490 ;
        RECT 651.000 20.070 651.260 20.390 ;
        RECT 677.680 20.070 677.940 20.390 ;
        RECT 651.060 2.400 651.200 20.070 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 916.850 37.980 917.170 38.040 ;
        RECT 989.990 37.980 990.310 38.040 ;
        RECT 916.850 37.840 990.310 37.980 ;
        RECT 916.850 37.780 917.170 37.840 ;
        RECT 989.990 37.780 990.310 37.840 ;
      LAYER via ;
        RECT 916.880 37.780 917.140 38.040 ;
        RECT 990.020 37.780 990.280 38.040 ;
      LAYER met2 ;
        RECT 917.230 960.570 917.510 964.000 ;
        RECT 916.940 960.430 917.510 960.570 ;
        RECT 916.940 38.070 917.080 960.430 ;
        RECT 917.230 960.000 917.510 960.430 ;
        RECT 916.880 37.750 917.140 38.070 ;
        RECT 990.020 37.750 990.280 38.070 ;
        RECT 990.080 2.400 990.220 37.750 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 930.650 31.180 930.970 31.240 ;
        RECT 1007.930 31.180 1008.250 31.240 ;
        RECT 930.650 31.040 1008.250 31.180 ;
        RECT 930.650 30.980 930.970 31.040 ;
        RECT 1007.930 30.980 1008.250 31.040 ;
      LAYER via ;
        RECT 930.680 30.980 930.940 31.240 ;
        RECT 1007.960 30.980 1008.220 31.240 ;
      LAYER met2 ;
        RECT 929.650 960.570 929.930 964.000 ;
        RECT 929.650 960.430 930.880 960.570 ;
        RECT 929.650 960.000 929.930 960.430 ;
        RECT 930.740 31.270 930.880 960.430 ;
        RECT 930.680 30.950 930.940 31.270 ;
        RECT 1007.960 30.950 1008.220 31.270 ;
        RECT 1008.020 16.730 1008.160 30.950 ;
        RECT 1007.560 16.590 1008.160 16.730 ;
        RECT 1007.560 2.400 1007.700 16.590 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 944.910 51.580 945.230 51.640 ;
        RECT 1021.270 51.580 1021.590 51.640 ;
        RECT 944.910 51.440 1021.590 51.580 ;
        RECT 944.910 51.380 945.230 51.440 ;
        RECT 1021.270 51.380 1021.590 51.440 ;
      LAYER via ;
        RECT 944.940 51.380 945.200 51.640 ;
        RECT 1021.300 51.380 1021.560 51.640 ;
      LAYER met2 ;
        RECT 942.070 960.570 942.350 964.000 ;
        RECT 942.070 960.430 945.140 960.570 ;
        RECT 942.070 960.000 942.350 960.430 ;
        RECT 945.000 51.670 945.140 960.430 ;
        RECT 944.940 51.350 945.200 51.670 ;
        RECT 1021.300 51.350 1021.560 51.670 ;
        RECT 1021.360 16.730 1021.500 51.350 ;
        RECT 1021.360 16.590 1025.640 16.730 ;
        RECT 1025.500 2.400 1025.640 16.590 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.570 945.440 954.890 945.500 ;
        RECT 958.710 945.440 959.030 945.500 ;
        RECT 954.570 945.300 959.030 945.440 ;
        RECT 954.570 945.240 954.890 945.300 ;
        RECT 958.710 945.240 959.030 945.300 ;
        RECT 958.710 44.780 959.030 44.840 ;
        RECT 1043.350 44.780 1043.670 44.840 ;
        RECT 958.710 44.640 1043.670 44.780 ;
        RECT 958.710 44.580 959.030 44.640 ;
        RECT 1043.350 44.580 1043.670 44.640 ;
      LAYER via ;
        RECT 954.600 945.240 954.860 945.500 ;
        RECT 958.740 945.240 959.000 945.500 ;
        RECT 958.740 44.580 959.000 44.840 ;
        RECT 1043.380 44.580 1043.640 44.840 ;
      LAYER met2 ;
        RECT 954.490 960.500 954.770 964.000 ;
        RECT 954.490 960.000 954.800 960.500 ;
        RECT 954.660 945.530 954.800 960.000 ;
        RECT 954.600 945.210 954.860 945.530 ;
        RECT 958.740 945.210 959.000 945.530 ;
        RECT 958.800 44.870 958.940 945.210 ;
        RECT 958.740 44.550 959.000 44.870 ;
        RECT 1043.380 44.550 1043.640 44.870 ;
        RECT 1043.440 2.400 1043.580 44.550 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.990 946.460 967.310 946.520 ;
        RECT 972.510 946.460 972.830 946.520 ;
        RECT 966.990 946.320 972.830 946.460 ;
        RECT 966.990 946.260 967.310 946.320 ;
        RECT 972.510 946.260 972.830 946.320 ;
        RECT 972.510 24.040 972.830 24.100 ;
        RECT 1061.290 24.040 1061.610 24.100 ;
        RECT 972.510 23.900 1061.610 24.040 ;
        RECT 972.510 23.840 972.830 23.900 ;
        RECT 1061.290 23.840 1061.610 23.900 ;
      LAYER via ;
        RECT 967.020 946.260 967.280 946.520 ;
        RECT 972.540 946.260 972.800 946.520 ;
        RECT 972.540 23.840 972.800 24.100 ;
        RECT 1061.320 23.840 1061.580 24.100 ;
      LAYER met2 ;
        RECT 966.910 960.500 967.190 964.000 ;
        RECT 966.910 960.000 967.220 960.500 ;
        RECT 967.080 946.550 967.220 960.000 ;
        RECT 967.020 946.230 967.280 946.550 ;
        RECT 972.540 946.230 972.800 946.550 ;
        RECT 972.600 24.130 972.740 946.230 ;
        RECT 972.540 23.810 972.800 24.130 ;
        RECT 1061.320 23.810 1061.580 24.130 ;
        RECT 1061.380 2.400 1061.520 23.810 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.410 948.840 979.730 948.900 ;
        RECT 1065.890 948.840 1066.210 948.900 ;
        RECT 979.410 948.700 1066.210 948.840 ;
        RECT 979.410 948.640 979.730 948.700 ;
        RECT 1065.890 948.640 1066.210 948.700 ;
        RECT 1065.890 20.980 1066.210 21.040 ;
        RECT 1079.230 20.980 1079.550 21.040 ;
        RECT 1065.890 20.840 1079.550 20.980 ;
        RECT 1065.890 20.780 1066.210 20.840 ;
        RECT 1079.230 20.780 1079.550 20.840 ;
      LAYER via ;
        RECT 979.440 948.640 979.700 948.900 ;
        RECT 1065.920 948.640 1066.180 948.900 ;
        RECT 1065.920 20.780 1066.180 21.040 ;
        RECT 1079.260 20.780 1079.520 21.040 ;
      LAYER met2 ;
        RECT 979.330 960.500 979.610 964.000 ;
        RECT 979.330 960.000 979.640 960.500 ;
        RECT 979.500 948.930 979.640 960.000 ;
        RECT 979.440 948.610 979.700 948.930 ;
        RECT 1065.920 948.610 1066.180 948.930 ;
        RECT 1065.980 21.070 1066.120 948.610 ;
        RECT 1065.920 20.750 1066.180 21.070 ;
        RECT 1079.260 20.750 1079.520 21.070 ;
        RECT 1079.320 2.400 1079.460 20.750 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 992.750 37.980 993.070 38.040 ;
        RECT 992.750 37.840 1049.100 37.980 ;
        RECT 992.750 37.780 993.070 37.840 ;
        RECT 1048.960 37.640 1049.100 37.840 ;
        RECT 1048.960 37.500 1097.400 37.640 ;
        RECT 1096.710 36.960 1097.030 37.020 ;
        RECT 1097.260 36.960 1097.400 37.500 ;
        RECT 1096.710 36.820 1097.400 36.960 ;
        RECT 1096.710 36.760 1097.030 36.820 ;
      LAYER via ;
        RECT 992.780 37.780 993.040 38.040 ;
        RECT 1096.740 36.760 1097.000 37.020 ;
      LAYER met2 ;
        RECT 991.750 960.570 992.030 964.000 ;
        RECT 991.750 960.430 992.980 960.570 ;
        RECT 991.750 960.000 992.030 960.430 ;
        RECT 992.840 38.070 992.980 960.430 ;
        RECT 992.780 37.750 993.040 38.070 ;
        RECT 1096.740 36.730 1097.000 37.050 ;
        RECT 1096.800 2.400 1096.940 36.730 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 30.840 1007.330 30.900 ;
        RECT 1114.650 30.840 1114.970 30.900 ;
        RECT 1007.010 30.700 1114.970 30.840 ;
        RECT 1007.010 30.640 1007.330 30.700 ;
        RECT 1114.650 30.640 1114.970 30.700 ;
      LAYER via ;
        RECT 1007.040 30.640 1007.300 30.900 ;
        RECT 1114.680 30.640 1114.940 30.900 ;
      LAYER met2 ;
        RECT 1003.710 960.570 1003.990 964.000 ;
        RECT 1003.710 960.430 1007.240 960.570 ;
        RECT 1003.710 960.000 1003.990 960.430 ;
        RECT 1007.100 30.930 1007.240 960.430 ;
        RECT 1007.040 30.610 1007.300 30.930 ;
        RECT 1114.680 30.610 1114.940 30.930 ;
        RECT 1114.740 2.400 1114.880 30.610 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1016.210 947.140 1016.530 947.200 ;
        RECT 1020.810 947.140 1021.130 947.200 ;
        RECT 1016.210 947.000 1021.130 947.140 ;
        RECT 1016.210 946.940 1016.530 947.000 ;
        RECT 1020.810 946.940 1021.130 947.000 ;
        RECT 1020.810 58.720 1021.130 58.780 ;
        RECT 1131.670 58.720 1131.990 58.780 ;
        RECT 1020.810 58.580 1131.990 58.720 ;
        RECT 1020.810 58.520 1021.130 58.580 ;
        RECT 1131.670 58.520 1131.990 58.580 ;
      LAYER via ;
        RECT 1016.240 946.940 1016.500 947.200 ;
        RECT 1020.840 946.940 1021.100 947.200 ;
        RECT 1020.840 58.520 1021.100 58.780 ;
        RECT 1131.700 58.520 1131.960 58.780 ;
      LAYER met2 ;
        RECT 1016.130 960.500 1016.410 964.000 ;
        RECT 1016.130 960.000 1016.440 960.500 ;
        RECT 1016.300 947.230 1016.440 960.000 ;
        RECT 1016.240 946.910 1016.500 947.230 ;
        RECT 1020.840 946.910 1021.100 947.230 ;
        RECT 1020.900 58.810 1021.040 946.910 ;
        RECT 1020.840 58.490 1021.100 58.810 ;
        RECT 1131.700 58.490 1131.960 58.810 ;
        RECT 1131.760 16.730 1131.900 58.490 ;
        RECT 1131.760 16.590 1132.820 16.730 ;
        RECT 1132.680 2.400 1132.820 16.590 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1028.630 946.460 1028.950 946.520 ;
        RECT 1034.610 946.460 1034.930 946.520 ;
        RECT 1028.630 946.320 1034.930 946.460 ;
        RECT 1028.630 946.260 1028.950 946.320 ;
        RECT 1034.610 946.260 1034.930 946.320 ;
        RECT 1034.610 51.580 1034.930 51.640 ;
        RECT 1145.470 51.580 1145.790 51.640 ;
        RECT 1034.610 51.440 1145.790 51.580 ;
        RECT 1034.610 51.380 1034.930 51.440 ;
        RECT 1145.470 51.380 1145.790 51.440 ;
      LAYER via ;
        RECT 1028.660 946.260 1028.920 946.520 ;
        RECT 1034.640 946.260 1034.900 946.520 ;
        RECT 1034.640 51.380 1034.900 51.640 ;
        RECT 1145.500 51.380 1145.760 51.640 ;
      LAYER met2 ;
        RECT 1028.550 960.500 1028.830 964.000 ;
        RECT 1028.550 960.000 1028.860 960.500 ;
        RECT 1028.720 946.550 1028.860 960.000 ;
        RECT 1028.660 946.230 1028.920 946.550 ;
        RECT 1034.640 946.230 1034.900 946.550 ;
        RECT 1034.700 51.670 1034.840 946.230 ;
        RECT 1034.640 51.350 1034.900 51.670 ;
        RECT 1145.500 51.350 1145.760 51.670 ;
        RECT 1145.560 17.410 1145.700 51.350 ;
        RECT 1145.560 17.270 1150.760 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 16.220 669.230 16.280 ;
        RECT 691.450 16.220 691.770 16.280 ;
        RECT 668.910 16.080 691.770 16.220 ;
        RECT 668.910 16.020 669.230 16.080 ;
        RECT 691.450 16.020 691.770 16.080 ;
      LAYER via ;
        RECT 668.940 16.020 669.200 16.280 ;
        RECT 691.480 16.020 691.740 16.280 ;
      LAYER met2 ;
        RECT 694.590 960.570 694.870 964.000 ;
        RECT 691.540 960.430 694.870 960.570 ;
        RECT 691.540 16.310 691.680 960.430 ;
        RECT 694.590 960.000 694.870 960.430 ;
        RECT 668.940 15.990 669.200 16.310 ;
        RECT 691.480 15.990 691.740 16.310 ;
        RECT 669.000 2.400 669.140 15.990 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.050 65.520 1041.370 65.580 ;
        RECT 1166.170 65.520 1166.490 65.580 ;
        RECT 1041.050 65.380 1166.490 65.520 ;
        RECT 1041.050 65.320 1041.370 65.380 ;
        RECT 1166.170 65.320 1166.490 65.380 ;
      LAYER via ;
        RECT 1041.080 65.320 1041.340 65.580 ;
        RECT 1166.200 65.320 1166.460 65.580 ;
      LAYER met2 ;
        RECT 1040.970 960.500 1041.250 964.000 ;
        RECT 1040.970 960.000 1041.280 960.500 ;
        RECT 1041.140 65.610 1041.280 960.000 ;
        RECT 1041.080 65.290 1041.340 65.610 ;
        RECT 1166.200 65.290 1166.460 65.610 ;
        RECT 1166.260 17.410 1166.400 65.290 ;
        RECT 1166.260 17.270 1168.700 17.410 ;
        RECT 1168.560 2.400 1168.700 17.270 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1054.850 44.780 1055.170 44.840 ;
        RECT 1185.950 44.780 1186.270 44.840 ;
        RECT 1054.850 44.640 1186.270 44.780 ;
        RECT 1054.850 44.580 1055.170 44.640 ;
        RECT 1185.950 44.580 1186.270 44.640 ;
      LAYER via ;
        RECT 1054.880 44.580 1055.140 44.840 ;
        RECT 1185.980 44.580 1186.240 44.840 ;
      LAYER met2 ;
        RECT 1053.390 960.570 1053.670 964.000 ;
        RECT 1053.390 960.430 1055.080 960.570 ;
        RECT 1053.390 960.000 1053.670 960.430 ;
        RECT 1054.940 44.870 1055.080 960.430 ;
        RECT 1054.880 44.550 1055.140 44.870 ;
        RECT 1185.980 44.550 1186.240 44.870 ;
        RECT 1186.040 2.400 1186.180 44.550 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1067.730 945.780 1068.050 945.840 ;
        RECT 1107.290 945.780 1107.610 945.840 ;
        RECT 1067.730 945.640 1107.610 945.780 ;
        RECT 1067.730 945.580 1068.050 945.640 ;
        RECT 1107.290 945.580 1107.610 945.640 ;
        RECT 1107.290 24.040 1107.610 24.100 ;
        RECT 1203.890 24.040 1204.210 24.100 ;
        RECT 1107.290 23.900 1204.210 24.040 ;
        RECT 1107.290 23.840 1107.610 23.900 ;
        RECT 1203.890 23.840 1204.210 23.900 ;
      LAYER via ;
        RECT 1067.760 945.580 1068.020 945.840 ;
        RECT 1107.320 945.580 1107.580 945.840 ;
        RECT 1107.320 23.840 1107.580 24.100 ;
        RECT 1203.920 23.840 1204.180 24.100 ;
      LAYER met2 ;
        RECT 1065.810 960.570 1066.090 964.000 ;
        RECT 1065.810 960.430 1067.960 960.570 ;
        RECT 1065.810 960.000 1066.090 960.430 ;
        RECT 1067.820 945.870 1067.960 960.430 ;
        RECT 1067.760 945.550 1068.020 945.870 ;
        RECT 1107.320 945.550 1107.580 945.870 ;
        RECT 1107.380 24.130 1107.520 945.550 ;
        RECT 1107.320 23.810 1107.580 24.130 ;
        RECT 1203.920 23.810 1204.180 24.130 ;
        RECT 1203.980 2.400 1204.120 23.810 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1078.310 945.440 1078.630 945.500 ;
        RECT 1082.910 945.440 1083.230 945.500 ;
        RECT 1078.310 945.300 1083.230 945.440 ;
        RECT 1078.310 945.240 1078.630 945.300 ;
        RECT 1082.910 945.240 1083.230 945.300 ;
        RECT 1082.910 72.320 1083.230 72.380 ;
        RECT 1221.830 72.320 1222.150 72.380 ;
        RECT 1082.910 72.180 1222.150 72.320 ;
        RECT 1082.910 72.120 1083.230 72.180 ;
        RECT 1221.830 72.120 1222.150 72.180 ;
      LAYER via ;
        RECT 1078.340 945.240 1078.600 945.500 ;
        RECT 1082.940 945.240 1083.200 945.500 ;
        RECT 1082.940 72.120 1083.200 72.380 ;
        RECT 1221.860 72.120 1222.120 72.380 ;
      LAYER met2 ;
        RECT 1078.230 960.500 1078.510 964.000 ;
        RECT 1078.230 960.000 1078.540 960.500 ;
        RECT 1078.400 945.530 1078.540 960.000 ;
        RECT 1078.340 945.210 1078.600 945.530 ;
        RECT 1082.940 945.210 1083.200 945.530 ;
        RECT 1083.000 72.410 1083.140 945.210 ;
        RECT 1082.940 72.090 1083.200 72.410 ;
        RECT 1221.860 72.090 1222.120 72.410 ;
        RECT 1221.920 2.400 1222.060 72.090 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 945.440 1091.050 945.500 ;
        RECT 1096.710 945.440 1097.030 945.500 ;
        RECT 1090.730 945.300 1097.030 945.440 ;
        RECT 1090.730 945.240 1091.050 945.300 ;
        RECT 1096.710 945.240 1097.030 945.300 ;
        RECT 1096.710 37.980 1097.030 38.040 ;
        RECT 1239.770 37.980 1240.090 38.040 ;
        RECT 1096.710 37.840 1240.090 37.980 ;
        RECT 1096.710 37.780 1097.030 37.840 ;
        RECT 1239.770 37.780 1240.090 37.840 ;
      LAYER via ;
        RECT 1090.760 945.240 1091.020 945.500 ;
        RECT 1096.740 945.240 1097.000 945.500 ;
        RECT 1096.740 37.780 1097.000 38.040 ;
        RECT 1239.800 37.780 1240.060 38.040 ;
      LAYER met2 ;
        RECT 1090.650 960.500 1090.930 964.000 ;
        RECT 1090.650 960.000 1090.960 960.500 ;
        RECT 1090.820 945.530 1090.960 960.000 ;
        RECT 1090.760 945.210 1091.020 945.530 ;
        RECT 1096.740 945.210 1097.000 945.530 ;
        RECT 1096.800 38.070 1096.940 945.210 ;
        RECT 1096.740 37.750 1097.000 38.070 ;
        RECT 1239.800 37.750 1240.060 38.070 ;
        RECT 1239.860 2.400 1240.000 37.750 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1103.610 941.700 1103.930 941.760 ;
        RECT 1255.870 941.700 1256.190 941.760 ;
        RECT 1103.610 941.560 1256.190 941.700 ;
        RECT 1103.610 941.500 1103.930 941.560 ;
        RECT 1255.870 941.500 1256.190 941.560 ;
      LAYER via ;
        RECT 1103.640 941.500 1103.900 941.760 ;
        RECT 1255.900 941.500 1256.160 941.760 ;
      LAYER met2 ;
        RECT 1103.070 960.570 1103.350 964.000 ;
        RECT 1103.070 960.430 1103.840 960.570 ;
        RECT 1103.070 960.000 1103.350 960.430 ;
        RECT 1103.700 941.790 1103.840 960.430 ;
        RECT 1103.640 941.470 1103.900 941.790 ;
        RECT 1255.900 941.470 1256.160 941.790 ;
        RECT 1255.960 17.410 1256.100 941.470 ;
        RECT 1255.960 17.270 1257.480 17.410 ;
        RECT 1257.340 2.400 1257.480 17.270 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1115.570 948.840 1115.890 948.900 ;
        RECT 1210.790 948.840 1211.110 948.900 ;
        RECT 1115.570 948.700 1211.110 948.840 ;
        RECT 1115.570 948.640 1115.890 948.700 ;
        RECT 1210.790 948.640 1211.110 948.700 ;
        RECT 1210.790 24.040 1211.110 24.100 ;
        RECT 1275.190 24.040 1275.510 24.100 ;
        RECT 1210.790 23.900 1275.510 24.040 ;
        RECT 1210.790 23.840 1211.110 23.900 ;
        RECT 1275.190 23.840 1275.510 23.900 ;
      LAYER via ;
        RECT 1115.600 948.640 1115.860 948.900 ;
        RECT 1210.820 948.640 1211.080 948.900 ;
        RECT 1210.820 23.840 1211.080 24.100 ;
        RECT 1275.220 23.840 1275.480 24.100 ;
      LAYER met2 ;
        RECT 1115.490 960.500 1115.770 964.000 ;
        RECT 1115.490 960.000 1115.800 960.500 ;
        RECT 1115.660 948.930 1115.800 960.000 ;
        RECT 1115.600 948.610 1115.860 948.930 ;
        RECT 1210.820 948.610 1211.080 948.930 ;
        RECT 1210.880 24.130 1211.020 948.610 ;
        RECT 1210.820 23.810 1211.080 24.130 ;
        RECT 1275.220 23.810 1275.480 24.130 ;
        RECT 1275.280 2.400 1275.420 23.810 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 30.840 1131.530 30.900 ;
        RECT 1293.130 30.840 1293.450 30.900 ;
        RECT 1131.210 30.700 1293.450 30.840 ;
        RECT 1131.210 30.640 1131.530 30.700 ;
        RECT 1293.130 30.640 1293.450 30.700 ;
      LAYER via ;
        RECT 1131.240 30.640 1131.500 30.900 ;
        RECT 1293.160 30.640 1293.420 30.900 ;
      LAYER met2 ;
        RECT 1127.450 960.570 1127.730 964.000 ;
        RECT 1127.450 960.430 1131.440 960.570 ;
        RECT 1127.450 960.000 1127.730 960.430 ;
        RECT 1131.300 30.930 1131.440 960.430 ;
        RECT 1131.240 30.610 1131.500 30.930 ;
        RECT 1293.160 30.610 1293.420 30.930 ;
        RECT 1293.220 2.400 1293.360 30.610 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1139.950 945.440 1140.270 945.500 ;
        RECT 1145.010 945.440 1145.330 945.500 ;
        RECT 1139.950 945.300 1145.330 945.440 ;
        RECT 1139.950 945.240 1140.270 945.300 ;
        RECT 1145.010 945.240 1145.330 945.300 ;
        RECT 1145.010 58.720 1145.330 58.780 ;
        RECT 1311.530 58.720 1311.850 58.780 ;
        RECT 1145.010 58.580 1311.850 58.720 ;
        RECT 1145.010 58.520 1145.330 58.580 ;
        RECT 1311.530 58.520 1311.850 58.580 ;
      LAYER via ;
        RECT 1139.980 945.240 1140.240 945.500 ;
        RECT 1145.040 945.240 1145.300 945.500 ;
        RECT 1145.040 58.520 1145.300 58.780 ;
        RECT 1311.560 58.520 1311.820 58.780 ;
      LAYER met2 ;
        RECT 1139.870 960.500 1140.150 964.000 ;
        RECT 1139.870 960.000 1140.180 960.500 ;
        RECT 1140.040 945.530 1140.180 960.000 ;
        RECT 1139.980 945.210 1140.240 945.530 ;
        RECT 1145.040 945.210 1145.300 945.530 ;
        RECT 1145.100 58.810 1145.240 945.210 ;
        RECT 1145.040 58.490 1145.300 58.810 ;
        RECT 1311.560 58.490 1311.820 58.810 ;
        RECT 1311.620 17.410 1311.760 58.490 ;
        RECT 1311.160 17.270 1311.760 17.410 ;
        RECT 1311.160 2.400 1311.300 17.270 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.370 946.460 1152.690 946.520 ;
        RECT 1158.810 946.460 1159.130 946.520 ;
        RECT 1152.370 946.320 1159.130 946.460 ;
        RECT 1152.370 946.260 1152.690 946.320 ;
        RECT 1158.810 946.260 1159.130 946.320 ;
        RECT 1158.810 51.580 1159.130 51.640 ;
        RECT 1324.870 51.580 1325.190 51.640 ;
        RECT 1158.810 51.440 1325.190 51.580 ;
        RECT 1158.810 51.380 1159.130 51.440 ;
        RECT 1324.870 51.380 1325.190 51.440 ;
      LAYER via ;
        RECT 1152.400 946.260 1152.660 946.520 ;
        RECT 1158.840 946.260 1159.100 946.520 ;
        RECT 1158.840 51.380 1159.100 51.640 ;
        RECT 1324.900 51.380 1325.160 51.640 ;
      LAYER met2 ;
        RECT 1152.290 960.500 1152.570 964.000 ;
        RECT 1152.290 960.000 1152.600 960.500 ;
        RECT 1152.460 946.550 1152.600 960.000 ;
        RECT 1152.400 946.230 1152.660 946.550 ;
        RECT 1158.840 946.230 1159.100 946.550 ;
        RECT 1158.900 51.670 1159.040 946.230 ;
        RECT 1158.840 51.350 1159.100 51.670 ;
        RECT 1324.900 51.350 1325.160 51.670 ;
        RECT 1324.960 17.410 1325.100 51.350 ;
        RECT 1324.960 17.270 1329.240 17.410 ;
        RECT 1329.100 2.400 1329.240 17.270 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 17.580 686.710 17.640 ;
        RECT 703.870 17.580 704.190 17.640 ;
        RECT 686.390 17.440 704.190 17.580 ;
        RECT 686.390 17.380 686.710 17.440 ;
        RECT 703.870 17.380 704.190 17.440 ;
      LAYER via ;
        RECT 686.420 17.380 686.680 17.640 ;
        RECT 703.900 17.380 704.160 17.640 ;
      LAYER met2 ;
        RECT 707.010 960.570 707.290 964.000 ;
        RECT 703.960 960.430 707.290 960.570 ;
        RECT 703.960 17.670 704.100 960.430 ;
        RECT 707.010 960.000 707.290 960.430 ;
        RECT 686.420 17.350 686.680 17.670 ;
        RECT 703.900 17.350 704.160 17.670 ;
        RECT 686.480 2.400 686.620 17.350 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 79.460 1166.030 79.520 ;
        RECT 1345.570 79.460 1345.890 79.520 ;
        RECT 1165.710 79.320 1345.890 79.460 ;
        RECT 1165.710 79.260 1166.030 79.320 ;
        RECT 1345.570 79.260 1345.890 79.320 ;
      LAYER via ;
        RECT 1165.740 79.260 1166.000 79.520 ;
        RECT 1345.600 79.260 1345.860 79.520 ;
      LAYER met2 ;
        RECT 1164.710 960.570 1164.990 964.000 ;
        RECT 1164.710 960.430 1165.940 960.570 ;
        RECT 1164.710 960.000 1164.990 960.430 ;
        RECT 1165.800 79.550 1165.940 960.430 ;
        RECT 1165.740 79.230 1166.000 79.550 ;
        RECT 1345.600 79.230 1345.860 79.550 ;
        RECT 1345.660 17.410 1345.800 79.230 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1177.210 934.900 1177.530 934.960 ;
        RECT 1359.370 934.900 1359.690 934.960 ;
        RECT 1177.210 934.760 1359.690 934.900 ;
        RECT 1177.210 934.700 1177.530 934.760 ;
        RECT 1359.370 934.700 1359.690 934.760 ;
      LAYER via ;
        RECT 1177.240 934.700 1177.500 934.960 ;
        RECT 1359.400 934.700 1359.660 934.960 ;
      LAYER met2 ;
        RECT 1177.130 960.500 1177.410 964.000 ;
        RECT 1177.130 960.000 1177.440 960.500 ;
        RECT 1177.300 934.990 1177.440 960.000 ;
        RECT 1177.240 934.670 1177.500 934.990 ;
        RECT 1359.400 934.670 1359.660 934.990 ;
        RECT 1359.460 17.410 1359.600 934.670 ;
        RECT 1359.460 17.270 1364.660 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1189.630 949.860 1189.950 949.920 ;
        RECT 1193.310 949.860 1193.630 949.920 ;
        RECT 1189.630 949.720 1193.630 949.860 ;
        RECT 1189.630 949.660 1189.950 949.720 ;
        RECT 1193.310 949.660 1193.630 949.720 ;
        RECT 1193.310 45.120 1193.630 45.180 ;
        RECT 1382.370 45.120 1382.690 45.180 ;
        RECT 1193.310 44.980 1382.690 45.120 ;
        RECT 1193.310 44.920 1193.630 44.980 ;
        RECT 1382.370 44.920 1382.690 44.980 ;
      LAYER via ;
        RECT 1189.660 949.660 1189.920 949.920 ;
        RECT 1193.340 949.660 1193.600 949.920 ;
        RECT 1193.340 44.920 1193.600 45.180 ;
        RECT 1382.400 44.920 1382.660 45.180 ;
      LAYER met2 ;
        RECT 1189.550 960.500 1189.830 964.000 ;
        RECT 1189.550 960.000 1189.860 960.500 ;
        RECT 1189.720 949.950 1189.860 960.000 ;
        RECT 1189.660 949.630 1189.920 949.950 ;
        RECT 1193.340 949.630 1193.600 949.950 ;
        RECT 1193.400 45.210 1193.540 949.630 ;
        RECT 1193.340 44.890 1193.600 45.210 ;
        RECT 1382.400 44.890 1382.660 45.210 ;
        RECT 1382.460 2.400 1382.600 44.890 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.050 949.180 1202.370 949.240 ;
        RECT 1279.790 949.180 1280.110 949.240 ;
        RECT 1202.050 949.040 1280.110 949.180 ;
        RECT 1202.050 948.980 1202.370 949.040 ;
        RECT 1279.790 948.980 1280.110 949.040 ;
        RECT 1279.790 24.040 1280.110 24.100 ;
        RECT 1400.310 24.040 1400.630 24.100 ;
        RECT 1279.790 23.900 1400.630 24.040 ;
        RECT 1279.790 23.840 1280.110 23.900 ;
        RECT 1400.310 23.840 1400.630 23.900 ;
      LAYER via ;
        RECT 1202.080 948.980 1202.340 949.240 ;
        RECT 1279.820 948.980 1280.080 949.240 ;
        RECT 1279.820 23.840 1280.080 24.100 ;
        RECT 1400.340 23.840 1400.600 24.100 ;
      LAYER met2 ;
        RECT 1201.970 960.500 1202.250 964.000 ;
        RECT 1201.970 960.000 1202.280 960.500 ;
        RECT 1202.140 949.270 1202.280 960.000 ;
        RECT 1202.080 948.950 1202.340 949.270 ;
        RECT 1279.820 948.950 1280.080 949.270 ;
        RECT 1279.880 24.130 1280.020 948.950 ;
        RECT 1279.820 23.810 1280.080 24.130 ;
        RECT 1400.340 23.810 1400.600 24.130 ;
        RECT 1400.400 2.400 1400.540 23.810 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.470 945.440 1214.790 945.500 ;
        RECT 1220.910 945.440 1221.230 945.500 ;
        RECT 1214.470 945.300 1221.230 945.440 ;
        RECT 1214.470 945.240 1214.790 945.300 ;
        RECT 1220.910 945.240 1221.230 945.300 ;
        RECT 1220.910 65.520 1221.230 65.580 ;
        RECT 1414.570 65.520 1414.890 65.580 ;
        RECT 1220.910 65.380 1414.890 65.520 ;
        RECT 1220.910 65.320 1221.230 65.380 ;
        RECT 1414.570 65.320 1414.890 65.380 ;
      LAYER via ;
        RECT 1214.500 945.240 1214.760 945.500 ;
        RECT 1220.940 945.240 1221.200 945.500 ;
        RECT 1220.940 65.320 1221.200 65.580 ;
        RECT 1414.600 65.320 1414.860 65.580 ;
      LAYER met2 ;
        RECT 1214.390 960.500 1214.670 964.000 ;
        RECT 1214.390 960.000 1214.700 960.500 ;
        RECT 1214.560 945.530 1214.700 960.000 ;
        RECT 1214.500 945.210 1214.760 945.530 ;
        RECT 1220.940 945.210 1221.200 945.530 ;
        RECT 1221.000 65.610 1221.140 945.210 ;
        RECT 1220.940 65.290 1221.200 65.610 ;
        RECT 1414.600 65.290 1414.860 65.610 ;
        RECT 1414.660 16.730 1414.800 65.290 ;
        RECT 1414.660 16.590 1418.480 16.730 ;
        RECT 1418.340 2.400 1418.480 16.590 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.810 72.320 1228.130 72.380 ;
        RECT 1435.730 72.320 1436.050 72.380 ;
        RECT 1227.810 72.180 1436.050 72.320 ;
        RECT 1227.810 72.120 1228.130 72.180 ;
        RECT 1435.730 72.120 1436.050 72.180 ;
      LAYER via ;
        RECT 1227.840 72.120 1228.100 72.380 ;
        RECT 1435.760 72.120 1436.020 72.380 ;
      LAYER met2 ;
        RECT 1226.810 960.570 1227.090 964.000 ;
        RECT 1226.810 960.430 1228.040 960.570 ;
        RECT 1226.810 960.000 1227.090 960.430 ;
        RECT 1227.900 72.410 1228.040 960.430 ;
        RECT 1227.840 72.090 1228.100 72.410 ;
        RECT 1435.760 72.090 1436.020 72.410 ;
        RECT 1435.820 2.400 1435.960 72.090 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 37.980 1241.930 38.040 ;
        RECT 1453.670 37.980 1453.990 38.040 ;
        RECT 1241.610 37.840 1453.990 37.980 ;
        RECT 1241.610 37.780 1241.930 37.840 ;
        RECT 1453.670 37.780 1453.990 37.840 ;
      LAYER via ;
        RECT 1241.640 37.780 1241.900 38.040 ;
        RECT 1453.700 37.780 1453.960 38.040 ;
      LAYER met2 ;
        RECT 1238.770 960.570 1239.050 964.000 ;
        RECT 1238.770 960.430 1241.840 960.570 ;
        RECT 1238.770 960.000 1239.050 960.430 ;
        RECT 1241.700 38.070 1241.840 960.430 ;
        RECT 1241.640 37.750 1241.900 38.070 ;
        RECT 1453.700 37.750 1453.960 38.070 ;
        RECT 1453.760 2.400 1453.900 37.750 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.270 947.480 1251.590 947.540 ;
        RECT 1255.410 947.480 1255.730 947.540 ;
        RECT 1251.270 947.340 1255.730 947.480 ;
        RECT 1251.270 947.280 1251.590 947.340 ;
        RECT 1255.410 947.280 1255.730 947.340 ;
        RECT 1255.410 86.600 1255.730 86.660 ;
        RECT 1469.770 86.600 1470.090 86.660 ;
        RECT 1255.410 86.460 1470.090 86.600 ;
        RECT 1255.410 86.400 1255.730 86.460 ;
        RECT 1469.770 86.400 1470.090 86.460 ;
      LAYER via ;
        RECT 1251.300 947.280 1251.560 947.540 ;
        RECT 1255.440 947.280 1255.700 947.540 ;
        RECT 1255.440 86.400 1255.700 86.660 ;
        RECT 1469.800 86.400 1470.060 86.660 ;
      LAYER met2 ;
        RECT 1251.190 960.500 1251.470 964.000 ;
        RECT 1251.190 960.000 1251.500 960.500 ;
        RECT 1251.360 947.570 1251.500 960.000 ;
        RECT 1251.300 947.250 1251.560 947.570 ;
        RECT 1255.440 947.250 1255.700 947.570 ;
        RECT 1255.500 86.690 1255.640 947.250 ;
        RECT 1255.440 86.370 1255.700 86.690 ;
        RECT 1469.800 86.370 1470.060 86.690 ;
        RECT 1469.860 17.410 1470.000 86.370 ;
        RECT 1469.860 17.270 1471.840 17.410 ;
        RECT 1471.700 2.400 1471.840 17.270 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1263.690 941.700 1264.010 941.760 ;
        RECT 1483.570 941.700 1483.890 941.760 ;
        RECT 1263.690 941.560 1483.890 941.700 ;
        RECT 1263.690 941.500 1264.010 941.560 ;
        RECT 1483.570 941.500 1483.890 941.560 ;
        RECT 1483.570 17.580 1483.890 17.640 ;
        RECT 1489.550 17.580 1489.870 17.640 ;
        RECT 1483.570 17.440 1489.870 17.580 ;
        RECT 1483.570 17.380 1483.890 17.440 ;
        RECT 1489.550 17.380 1489.870 17.440 ;
      LAYER via ;
        RECT 1263.720 941.500 1263.980 941.760 ;
        RECT 1483.600 941.500 1483.860 941.760 ;
        RECT 1483.600 17.380 1483.860 17.640 ;
        RECT 1489.580 17.380 1489.840 17.640 ;
      LAYER met2 ;
        RECT 1263.610 960.500 1263.890 964.000 ;
        RECT 1263.610 960.000 1263.920 960.500 ;
        RECT 1263.780 941.790 1263.920 960.000 ;
        RECT 1263.720 941.470 1263.980 941.790 ;
        RECT 1483.600 941.470 1483.860 941.790 ;
        RECT 1483.660 17.670 1483.800 941.470 ;
        RECT 1483.600 17.350 1483.860 17.670 ;
        RECT 1489.580 17.350 1489.840 17.670 ;
        RECT 1489.640 2.400 1489.780 17.350 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 93.060 1276.430 93.120 ;
        RECT 1504.270 93.060 1504.590 93.120 ;
        RECT 1276.110 92.920 1504.590 93.060 ;
        RECT 1276.110 92.860 1276.430 92.920 ;
        RECT 1504.270 92.860 1504.590 92.920 ;
      LAYER via ;
        RECT 1276.140 92.860 1276.400 93.120 ;
        RECT 1504.300 92.860 1504.560 93.120 ;
      LAYER met2 ;
        RECT 1276.030 960.500 1276.310 964.000 ;
        RECT 1276.030 960.000 1276.340 960.500 ;
        RECT 1276.200 93.150 1276.340 960.000 ;
        RECT 1276.140 92.830 1276.400 93.150 ;
        RECT 1504.300 92.830 1504.560 93.150 ;
        RECT 1504.360 17.410 1504.500 92.830 ;
        RECT 1504.360 17.270 1507.260 17.410 ;
        RECT 1507.120 2.400 1507.260 17.270 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 20.300 704.650 20.360 ;
        RECT 717.670 20.300 717.990 20.360 ;
        RECT 704.330 20.160 717.990 20.300 ;
        RECT 704.330 20.100 704.650 20.160 ;
        RECT 717.670 20.100 717.990 20.160 ;
      LAYER via ;
        RECT 704.360 20.100 704.620 20.360 ;
        RECT 717.700 20.100 717.960 20.360 ;
      LAYER met2 ;
        RECT 719.430 960.570 719.710 964.000 ;
        RECT 717.760 960.430 719.710 960.570 ;
        RECT 717.760 20.390 717.900 960.430 ;
        RECT 719.430 960.000 719.710 960.430 ;
        RECT 704.360 20.070 704.620 20.390 ;
        RECT 717.700 20.070 717.960 20.390 ;
        RECT 704.420 2.400 704.560 20.070 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1288.530 949.180 1288.850 949.240 ;
        RECT 1507.490 949.180 1507.810 949.240 ;
        RECT 1288.530 949.040 1507.810 949.180 ;
        RECT 1288.530 948.980 1288.850 949.040 ;
        RECT 1507.490 948.980 1507.810 949.040 ;
        RECT 1507.490 96.460 1507.810 96.520 ;
        RECT 1525.430 96.460 1525.750 96.520 ;
        RECT 1507.490 96.320 1525.750 96.460 ;
        RECT 1507.490 96.260 1507.810 96.320 ;
        RECT 1525.430 96.260 1525.750 96.320 ;
      LAYER via ;
        RECT 1288.560 948.980 1288.820 949.240 ;
        RECT 1507.520 948.980 1507.780 949.240 ;
        RECT 1507.520 96.260 1507.780 96.520 ;
        RECT 1525.460 96.260 1525.720 96.520 ;
      LAYER met2 ;
        RECT 1288.450 960.500 1288.730 964.000 ;
        RECT 1288.450 960.000 1288.760 960.500 ;
        RECT 1288.620 949.270 1288.760 960.000 ;
        RECT 1288.560 948.950 1288.820 949.270 ;
        RECT 1507.520 948.950 1507.780 949.270 ;
        RECT 1507.580 96.550 1507.720 948.950 ;
        RECT 1507.520 96.230 1507.780 96.550 ;
        RECT 1525.460 96.230 1525.720 96.550 ;
        RECT 1525.520 7.210 1525.660 96.230 ;
        RECT 1525.060 7.070 1525.660 7.210 ;
        RECT 1525.060 2.400 1525.200 7.070 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1303.710 30.840 1304.030 30.900 ;
        RECT 1542.910 30.840 1543.230 30.900 ;
        RECT 1303.710 30.700 1543.230 30.840 ;
        RECT 1303.710 30.640 1304.030 30.700 ;
        RECT 1542.910 30.640 1543.230 30.700 ;
      LAYER via ;
        RECT 1303.740 30.640 1304.000 30.900 ;
        RECT 1542.940 30.640 1543.200 30.900 ;
      LAYER met2 ;
        RECT 1300.870 960.570 1301.150 964.000 ;
        RECT 1300.870 960.430 1303.940 960.570 ;
        RECT 1300.870 960.000 1301.150 960.430 ;
        RECT 1303.800 30.930 1303.940 960.430 ;
        RECT 1303.740 30.610 1304.000 30.930 ;
        RECT 1542.940 30.610 1543.200 30.930 ;
        RECT 1543.000 2.400 1543.140 30.610 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.370 945.440 1313.690 945.500 ;
        RECT 1317.510 945.440 1317.830 945.500 ;
        RECT 1313.370 945.300 1317.830 945.440 ;
        RECT 1313.370 945.240 1313.690 945.300 ;
        RECT 1317.510 945.240 1317.830 945.300 ;
        RECT 1317.510 58.720 1317.830 58.780 ;
        RECT 1559.470 58.720 1559.790 58.780 ;
        RECT 1317.510 58.580 1559.790 58.720 ;
        RECT 1317.510 58.520 1317.830 58.580 ;
        RECT 1559.470 58.520 1559.790 58.580 ;
      LAYER via ;
        RECT 1313.400 945.240 1313.660 945.500 ;
        RECT 1317.540 945.240 1317.800 945.500 ;
        RECT 1317.540 58.520 1317.800 58.780 ;
        RECT 1559.500 58.520 1559.760 58.780 ;
      LAYER met2 ;
        RECT 1313.290 960.500 1313.570 964.000 ;
        RECT 1313.290 960.000 1313.600 960.500 ;
        RECT 1313.460 945.530 1313.600 960.000 ;
        RECT 1313.400 945.210 1313.660 945.530 ;
        RECT 1317.540 945.210 1317.800 945.530 ;
        RECT 1317.600 58.810 1317.740 945.210 ;
        RECT 1317.540 58.490 1317.800 58.810 ;
        RECT 1559.500 58.490 1559.760 58.810 ;
        RECT 1559.560 16.730 1559.700 58.490 ;
        RECT 1559.560 16.590 1561.080 16.730 ;
        RECT 1560.940 2.400 1561.080 16.590 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.790 946.460 1326.110 946.520 ;
        RECT 1331.310 946.460 1331.630 946.520 ;
        RECT 1325.790 946.320 1331.630 946.460 ;
        RECT 1325.790 946.260 1326.110 946.320 ;
        RECT 1331.310 946.260 1331.630 946.320 ;
        RECT 1331.310 99.860 1331.630 99.920 ;
        RECT 1573.270 99.860 1573.590 99.920 ;
        RECT 1331.310 99.720 1573.590 99.860 ;
        RECT 1331.310 99.660 1331.630 99.720 ;
        RECT 1573.270 99.660 1573.590 99.720 ;
      LAYER via ;
        RECT 1325.820 946.260 1326.080 946.520 ;
        RECT 1331.340 946.260 1331.600 946.520 ;
        RECT 1331.340 99.660 1331.600 99.920 ;
        RECT 1573.300 99.660 1573.560 99.920 ;
      LAYER met2 ;
        RECT 1325.710 960.500 1325.990 964.000 ;
        RECT 1325.710 960.000 1326.020 960.500 ;
        RECT 1325.880 946.550 1326.020 960.000 ;
        RECT 1325.820 946.230 1326.080 946.550 ;
        RECT 1331.340 946.230 1331.600 946.550 ;
        RECT 1331.400 99.950 1331.540 946.230 ;
        RECT 1331.340 99.630 1331.600 99.950 ;
        RECT 1573.300 99.630 1573.560 99.950 ;
        RECT 1573.360 16.730 1573.500 99.630 ;
        RECT 1573.360 16.590 1579.020 16.730 ;
        RECT 1578.880 2.400 1579.020 16.590 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1338.210 51.580 1338.530 51.640 ;
        RECT 1593.970 51.580 1594.290 51.640 ;
        RECT 1338.210 51.440 1594.290 51.580 ;
        RECT 1338.210 51.380 1338.530 51.440 ;
        RECT 1593.970 51.380 1594.290 51.440 ;
      LAYER via ;
        RECT 1338.240 51.380 1338.500 51.640 ;
        RECT 1594.000 51.380 1594.260 51.640 ;
      LAYER met2 ;
        RECT 1338.130 960.500 1338.410 964.000 ;
        RECT 1338.130 960.000 1338.440 960.500 ;
        RECT 1338.300 51.670 1338.440 960.000 ;
        RECT 1338.240 51.350 1338.500 51.670 ;
        RECT 1594.000 51.350 1594.260 51.670 ;
        RECT 1594.060 17.410 1594.200 51.350 ;
        RECT 1594.060 17.270 1596.500 17.410 ;
        RECT 1596.360 2.400 1596.500 17.270 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.010 79.460 1352.330 79.520 ;
        RECT 1608.230 79.460 1608.550 79.520 ;
        RECT 1352.010 79.320 1608.550 79.460 ;
        RECT 1352.010 79.260 1352.330 79.320 ;
        RECT 1608.230 79.260 1608.550 79.320 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1608.230 17.780 1614.530 17.920 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
      LAYER via ;
        RECT 1352.040 79.260 1352.300 79.520 ;
        RECT 1608.260 79.260 1608.520 79.520 ;
        RECT 1608.260 17.720 1608.520 17.980 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
      LAYER met2 ;
        RECT 1350.090 960.570 1350.370 964.000 ;
        RECT 1350.090 960.430 1352.240 960.570 ;
        RECT 1350.090 960.000 1350.370 960.430 ;
        RECT 1352.100 79.550 1352.240 960.430 ;
        RECT 1352.040 79.230 1352.300 79.550 ;
        RECT 1608.260 79.230 1608.520 79.550 ;
        RECT 1608.320 18.010 1608.460 79.230 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1614.300 2.400 1614.440 17.690 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 44.780 1366.130 44.840 ;
        RECT 1632.150 44.780 1632.470 44.840 ;
        RECT 1365.810 44.640 1632.470 44.780 ;
        RECT 1365.810 44.580 1366.130 44.640 ;
        RECT 1632.150 44.580 1632.470 44.640 ;
      LAYER via ;
        RECT 1365.840 44.580 1366.100 44.840 ;
        RECT 1632.180 44.580 1632.440 44.840 ;
      LAYER met2 ;
        RECT 1362.510 960.570 1362.790 964.000 ;
        RECT 1362.510 960.430 1366.040 960.570 ;
        RECT 1362.510 960.000 1362.790 960.430 ;
        RECT 1365.900 44.870 1366.040 960.430 ;
        RECT 1365.840 44.550 1366.100 44.870 ;
        RECT 1632.180 44.550 1632.440 44.870 ;
        RECT 1632.240 2.400 1632.380 44.550 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1375.010 948.840 1375.330 948.900 ;
        RECT 1403.990 948.840 1404.310 948.900 ;
        RECT 1375.010 948.700 1404.310 948.840 ;
        RECT 1375.010 948.640 1375.330 948.700 ;
        RECT 1403.990 948.640 1404.310 948.700 ;
        RECT 1403.990 24.720 1404.310 24.780 ;
        RECT 1403.990 24.580 1459.420 24.720 ;
        RECT 1403.990 24.520 1404.310 24.580 ;
        RECT 1459.280 24.380 1459.420 24.580 ;
        RECT 1650.090 24.380 1650.410 24.440 ;
        RECT 1459.280 24.240 1650.410 24.380 ;
        RECT 1650.090 24.180 1650.410 24.240 ;
      LAYER via ;
        RECT 1375.040 948.640 1375.300 948.900 ;
        RECT 1404.020 948.640 1404.280 948.900 ;
        RECT 1404.020 24.520 1404.280 24.780 ;
        RECT 1650.120 24.180 1650.380 24.440 ;
      LAYER met2 ;
        RECT 1374.930 960.500 1375.210 964.000 ;
        RECT 1374.930 960.000 1375.240 960.500 ;
        RECT 1375.100 948.930 1375.240 960.000 ;
        RECT 1375.040 948.610 1375.300 948.930 ;
        RECT 1404.020 948.610 1404.280 948.930 ;
        RECT 1404.080 24.810 1404.220 948.610 ;
        RECT 1404.020 24.490 1404.280 24.810 ;
        RECT 1650.120 24.150 1650.380 24.470 ;
        RECT 1650.180 2.400 1650.320 24.150 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1387.430 946.800 1387.750 946.860 ;
        RECT 1393.410 946.800 1393.730 946.860 ;
        RECT 1387.430 946.660 1393.730 946.800 ;
        RECT 1387.430 946.600 1387.750 946.660 ;
        RECT 1393.410 946.600 1393.730 946.660 ;
        RECT 1393.410 107.340 1393.730 107.400 ;
        RECT 1662.970 107.340 1663.290 107.400 ;
        RECT 1393.410 107.200 1663.290 107.340 ;
        RECT 1393.410 107.140 1393.730 107.200 ;
        RECT 1662.970 107.140 1663.290 107.200 ;
      LAYER via ;
        RECT 1387.460 946.600 1387.720 946.860 ;
        RECT 1393.440 946.600 1393.700 946.860 ;
        RECT 1393.440 107.140 1393.700 107.400 ;
        RECT 1663.000 107.140 1663.260 107.400 ;
      LAYER met2 ;
        RECT 1387.350 960.500 1387.630 964.000 ;
        RECT 1387.350 960.000 1387.660 960.500 ;
        RECT 1387.520 946.890 1387.660 960.000 ;
        RECT 1387.460 946.570 1387.720 946.890 ;
        RECT 1393.440 946.570 1393.700 946.890 ;
        RECT 1393.500 107.430 1393.640 946.570 ;
        RECT 1393.440 107.110 1393.700 107.430 ;
        RECT 1663.000 107.110 1663.260 107.430 ;
        RECT 1663.060 17.410 1663.200 107.110 ;
        RECT 1663.060 17.270 1668.260 17.410 ;
        RECT 1668.120 2.400 1668.260 17.270 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 113.800 1400.630 113.860 ;
        RECT 1683.670 113.800 1683.990 113.860 ;
        RECT 1400.310 113.660 1683.990 113.800 ;
        RECT 1400.310 113.600 1400.630 113.660 ;
        RECT 1683.670 113.600 1683.990 113.660 ;
      LAYER via ;
        RECT 1400.340 113.600 1400.600 113.860 ;
        RECT 1683.700 113.600 1683.960 113.860 ;
      LAYER met2 ;
        RECT 1399.770 960.570 1400.050 964.000 ;
        RECT 1399.770 960.430 1400.540 960.570 ;
        RECT 1399.770 960.000 1400.050 960.430 ;
        RECT 1400.400 113.890 1400.540 960.430 ;
        RECT 1400.340 113.570 1400.600 113.890 ;
        RECT 1683.700 113.570 1683.960 113.890 ;
        RECT 1683.760 17.410 1683.900 113.570 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 20.640 722.590 20.700 ;
        RECT 731.930 20.640 732.250 20.700 ;
        RECT 722.270 20.500 732.250 20.640 ;
        RECT 722.270 20.440 722.590 20.500 ;
        RECT 731.930 20.440 732.250 20.500 ;
      LAYER via ;
        RECT 722.300 20.440 722.560 20.700 ;
        RECT 731.960 20.440 732.220 20.700 ;
      LAYER met2 ;
        RECT 731.850 960.500 732.130 964.000 ;
        RECT 731.850 960.000 732.160 960.500 ;
        RECT 732.020 20.730 732.160 960.000 ;
        RECT 722.300 20.410 722.560 20.730 ;
        RECT 731.960 20.410 732.220 20.730 ;
        RECT 722.360 2.400 722.500 20.410 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 120.600 1414.430 120.660 ;
        RECT 1697.930 120.600 1698.250 120.660 ;
        RECT 1414.110 120.460 1698.250 120.600 ;
        RECT 1414.110 120.400 1414.430 120.460 ;
        RECT 1697.930 120.400 1698.250 120.460 ;
      LAYER via ;
        RECT 1414.140 120.400 1414.400 120.660 ;
        RECT 1697.960 120.400 1698.220 120.660 ;
      LAYER met2 ;
        RECT 1412.190 960.570 1412.470 964.000 ;
        RECT 1412.190 960.430 1414.340 960.570 ;
        RECT 1412.190 960.000 1412.470 960.430 ;
        RECT 1414.200 120.690 1414.340 960.430 ;
        RECT 1414.140 120.370 1414.400 120.690 ;
        RECT 1697.960 120.370 1698.220 120.690 ;
        RECT 1698.020 17.410 1698.160 120.370 ;
        RECT 1698.020 17.270 1703.680 17.410 ;
        RECT 1703.540 2.400 1703.680 17.270 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 65.520 1428.230 65.580 ;
        RECT 1718.170 65.520 1718.490 65.580 ;
        RECT 1427.910 65.380 1718.490 65.520 ;
        RECT 1427.910 65.320 1428.230 65.380 ;
        RECT 1718.170 65.320 1718.490 65.380 ;
      LAYER via ;
        RECT 1427.940 65.320 1428.200 65.580 ;
        RECT 1718.200 65.320 1718.460 65.580 ;
      LAYER met2 ;
        RECT 1424.610 960.570 1424.890 964.000 ;
        RECT 1424.610 960.430 1428.140 960.570 ;
        RECT 1424.610 960.000 1424.890 960.430 ;
        RECT 1428.000 65.610 1428.140 960.430 ;
        RECT 1427.940 65.290 1428.200 65.610 ;
        RECT 1718.200 65.290 1718.460 65.610 ;
        RECT 1718.260 17.410 1718.400 65.290 ;
        RECT 1718.260 17.270 1721.620 17.410 ;
        RECT 1721.480 2.400 1721.620 17.270 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.110 945.440 1437.430 945.500 ;
        RECT 1441.710 945.440 1442.030 945.500 ;
        RECT 1437.110 945.300 1442.030 945.440 ;
        RECT 1437.110 945.240 1437.430 945.300 ;
        RECT 1441.710 945.240 1442.030 945.300 ;
        RECT 1441.710 72.660 1442.030 72.720 ;
        RECT 1739.330 72.660 1739.650 72.720 ;
        RECT 1441.710 72.520 1739.650 72.660 ;
        RECT 1441.710 72.460 1442.030 72.520 ;
        RECT 1739.330 72.460 1739.650 72.520 ;
      LAYER via ;
        RECT 1437.140 945.240 1437.400 945.500 ;
        RECT 1441.740 945.240 1442.000 945.500 ;
        RECT 1441.740 72.460 1442.000 72.720 ;
        RECT 1739.360 72.460 1739.620 72.720 ;
      LAYER met2 ;
        RECT 1437.030 960.500 1437.310 964.000 ;
        RECT 1437.030 960.000 1437.340 960.500 ;
        RECT 1437.200 945.530 1437.340 960.000 ;
        RECT 1437.140 945.210 1437.400 945.530 ;
        RECT 1441.740 945.210 1442.000 945.530 ;
        RECT 1441.800 72.750 1441.940 945.210 ;
        RECT 1441.740 72.430 1442.000 72.750 ;
        RECT 1739.360 72.430 1739.620 72.750 ;
        RECT 1739.420 2.400 1739.560 72.430 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1449.530 945.440 1449.850 945.500 ;
        RECT 1455.510 945.440 1455.830 945.500 ;
        RECT 1449.530 945.300 1455.830 945.440 ;
        RECT 1449.530 945.240 1449.850 945.300 ;
        RECT 1455.510 945.240 1455.830 945.300 ;
        RECT 1455.510 37.980 1455.830 38.040 ;
        RECT 1756.810 37.980 1757.130 38.040 ;
        RECT 1455.510 37.840 1757.130 37.980 ;
        RECT 1455.510 37.780 1455.830 37.840 ;
        RECT 1756.810 37.780 1757.130 37.840 ;
      LAYER via ;
        RECT 1449.560 945.240 1449.820 945.500 ;
        RECT 1455.540 945.240 1455.800 945.500 ;
        RECT 1455.540 37.780 1455.800 38.040 ;
        RECT 1756.840 37.780 1757.100 38.040 ;
      LAYER met2 ;
        RECT 1449.450 960.500 1449.730 964.000 ;
        RECT 1449.450 960.000 1449.760 960.500 ;
        RECT 1449.620 945.530 1449.760 960.000 ;
        RECT 1449.560 945.210 1449.820 945.530 ;
        RECT 1455.540 945.210 1455.800 945.530 ;
        RECT 1455.600 38.070 1455.740 945.210 ;
        RECT 1455.540 37.750 1455.800 38.070 ;
        RECT 1756.840 37.750 1757.100 38.070 ;
        RECT 1756.900 2.400 1757.040 37.750 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 86.260 1462.730 86.320 ;
        RECT 1773.370 86.260 1773.690 86.320 ;
        RECT 1462.410 86.120 1773.690 86.260 ;
        RECT 1462.410 86.060 1462.730 86.120 ;
        RECT 1773.370 86.060 1773.690 86.120 ;
      LAYER via ;
        RECT 1462.440 86.060 1462.700 86.320 ;
        RECT 1773.400 86.060 1773.660 86.320 ;
      LAYER met2 ;
        RECT 1461.410 960.570 1461.690 964.000 ;
        RECT 1461.410 960.430 1462.640 960.570 ;
        RECT 1461.410 960.000 1461.690 960.430 ;
        RECT 1462.500 86.350 1462.640 960.430 ;
        RECT 1462.440 86.030 1462.700 86.350 ;
        RECT 1773.400 86.030 1773.660 86.350 ;
        RECT 1773.460 16.730 1773.600 86.030 ;
        RECT 1773.460 16.590 1774.980 16.730 ;
        RECT 1774.840 2.400 1774.980 16.590 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1473.910 948.840 1474.230 948.900 ;
        RECT 1762.790 948.840 1763.110 948.900 ;
        RECT 1473.910 948.700 1763.110 948.840 ;
        RECT 1473.910 948.640 1474.230 948.700 ;
        RECT 1762.790 948.640 1763.110 948.700 ;
        RECT 1762.790 24.380 1763.110 24.440 ;
        RECT 1792.690 24.380 1793.010 24.440 ;
        RECT 1762.790 24.240 1793.010 24.380 ;
        RECT 1762.790 24.180 1763.110 24.240 ;
        RECT 1792.690 24.180 1793.010 24.240 ;
      LAYER via ;
        RECT 1473.940 948.640 1474.200 948.900 ;
        RECT 1762.820 948.640 1763.080 948.900 ;
        RECT 1762.820 24.180 1763.080 24.440 ;
        RECT 1792.720 24.180 1792.980 24.440 ;
      LAYER met2 ;
        RECT 1473.830 960.500 1474.110 964.000 ;
        RECT 1473.830 960.000 1474.140 960.500 ;
        RECT 1474.000 948.930 1474.140 960.000 ;
        RECT 1473.940 948.610 1474.200 948.930 ;
        RECT 1762.820 948.610 1763.080 948.930 ;
        RECT 1762.880 24.470 1763.020 948.610 ;
        RECT 1762.820 24.150 1763.080 24.470 ;
        RECT 1792.720 24.150 1792.980 24.470 ;
        RECT 1792.780 2.400 1792.920 24.150 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 127.740 1490.330 127.800 ;
        RECT 1807.870 127.740 1808.190 127.800 ;
        RECT 1490.010 127.600 1808.190 127.740 ;
        RECT 1490.010 127.540 1490.330 127.600 ;
        RECT 1807.870 127.540 1808.190 127.600 ;
      LAYER via ;
        RECT 1490.040 127.540 1490.300 127.800 ;
        RECT 1807.900 127.540 1808.160 127.800 ;
      LAYER met2 ;
        RECT 1486.250 960.570 1486.530 964.000 ;
        RECT 1486.250 960.430 1490.240 960.570 ;
        RECT 1486.250 960.000 1486.530 960.430 ;
        RECT 1490.100 127.830 1490.240 960.430 ;
        RECT 1490.040 127.510 1490.300 127.830 ;
        RECT 1807.900 127.510 1808.160 127.830 ;
        RECT 1807.960 16.730 1808.100 127.510 ;
        RECT 1807.960 16.590 1810.860 16.730 ;
        RECT 1810.720 2.400 1810.860 16.590 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1498.750 946.800 1499.070 946.860 ;
        RECT 1503.810 946.800 1504.130 946.860 ;
        RECT 1498.750 946.660 1504.130 946.800 ;
        RECT 1498.750 946.600 1499.070 946.660 ;
        RECT 1503.810 946.600 1504.130 946.660 ;
        RECT 1503.810 134.540 1504.130 134.600 ;
        RECT 1829.030 134.540 1829.350 134.600 ;
        RECT 1503.810 134.400 1829.350 134.540 ;
        RECT 1503.810 134.340 1504.130 134.400 ;
        RECT 1829.030 134.340 1829.350 134.400 ;
      LAYER via ;
        RECT 1498.780 946.600 1499.040 946.860 ;
        RECT 1503.840 946.600 1504.100 946.860 ;
        RECT 1503.840 134.340 1504.100 134.600 ;
        RECT 1829.060 134.340 1829.320 134.600 ;
      LAYER met2 ;
        RECT 1498.670 960.500 1498.950 964.000 ;
        RECT 1498.670 960.000 1498.980 960.500 ;
        RECT 1498.840 946.890 1498.980 960.000 ;
        RECT 1498.780 946.570 1499.040 946.890 ;
        RECT 1503.840 946.570 1504.100 946.890 ;
        RECT 1503.900 134.630 1504.040 946.570 ;
        RECT 1503.840 134.310 1504.100 134.630 ;
        RECT 1829.060 134.310 1829.320 134.630 ;
        RECT 1829.120 17.410 1829.260 134.310 ;
        RECT 1828.660 17.270 1829.260 17.410 ;
        RECT 1828.660 2.400 1828.800 17.270 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1511.170 946.460 1511.490 946.520 ;
        RECT 1517.610 946.460 1517.930 946.520 ;
        RECT 1511.170 946.320 1517.930 946.460 ;
        RECT 1511.170 946.260 1511.490 946.320 ;
        RECT 1517.610 946.260 1517.930 946.320 ;
        RECT 1517.610 141.340 1517.930 141.400 ;
        RECT 1842.370 141.340 1842.690 141.400 ;
        RECT 1517.610 141.200 1842.690 141.340 ;
        RECT 1517.610 141.140 1517.930 141.200 ;
        RECT 1842.370 141.140 1842.690 141.200 ;
        RECT 1842.370 2.960 1842.690 3.020 ;
        RECT 1846.050 2.960 1846.370 3.020 ;
        RECT 1842.370 2.820 1846.370 2.960 ;
        RECT 1842.370 2.760 1842.690 2.820 ;
        RECT 1846.050 2.760 1846.370 2.820 ;
      LAYER via ;
        RECT 1511.200 946.260 1511.460 946.520 ;
        RECT 1517.640 946.260 1517.900 946.520 ;
        RECT 1517.640 141.140 1517.900 141.400 ;
        RECT 1842.400 141.140 1842.660 141.400 ;
        RECT 1842.400 2.760 1842.660 3.020 ;
        RECT 1846.080 2.760 1846.340 3.020 ;
      LAYER met2 ;
        RECT 1511.090 960.500 1511.370 964.000 ;
        RECT 1511.090 960.000 1511.400 960.500 ;
        RECT 1511.260 946.550 1511.400 960.000 ;
        RECT 1511.200 946.230 1511.460 946.550 ;
        RECT 1517.640 946.230 1517.900 946.550 ;
        RECT 1517.700 141.430 1517.840 946.230 ;
        RECT 1517.640 141.110 1517.900 141.430 ;
        RECT 1842.400 141.110 1842.660 141.430 ;
        RECT 1842.460 3.050 1842.600 141.110 ;
        RECT 1842.400 2.730 1842.660 3.050 ;
        RECT 1846.080 2.730 1846.340 3.050 ;
        RECT 1846.140 2.400 1846.280 2.730 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 148.140 1524.830 148.200 ;
        RECT 1863.070 148.140 1863.390 148.200 ;
        RECT 1524.510 148.000 1863.390 148.140 ;
        RECT 1524.510 147.940 1524.830 148.000 ;
        RECT 1863.070 147.940 1863.390 148.000 ;
        RECT 1863.070 2.960 1863.390 3.020 ;
        RECT 1863.990 2.960 1864.310 3.020 ;
        RECT 1863.070 2.820 1864.310 2.960 ;
        RECT 1863.070 2.760 1863.390 2.820 ;
        RECT 1863.990 2.760 1864.310 2.820 ;
      LAYER via ;
        RECT 1524.540 147.940 1524.800 148.200 ;
        RECT 1863.100 147.940 1863.360 148.200 ;
        RECT 1863.100 2.760 1863.360 3.020 ;
        RECT 1864.020 2.760 1864.280 3.020 ;
      LAYER met2 ;
        RECT 1523.510 960.570 1523.790 964.000 ;
        RECT 1523.510 960.430 1524.740 960.570 ;
        RECT 1523.510 960.000 1523.790 960.430 ;
        RECT 1524.600 148.230 1524.740 960.430 ;
        RECT 1524.540 147.910 1524.800 148.230 ;
        RECT 1863.100 147.910 1863.360 148.230 ;
        RECT 1863.160 3.050 1863.300 147.910 ;
        RECT 1863.100 2.730 1863.360 3.050 ;
        RECT 1864.020 2.730 1864.280 3.050 ;
        RECT 1864.080 2.400 1864.220 2.730 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 738.370 928.100 738.690 928.160 ;
        RECT 742.510 928.100 742.830 928.160 ;
        RECT 738.370 927.960 742.830 928.100 ;
        RECT 738.370 927.900 738.690 927.960 ;
        RECT 742.510 927.900 742.830 927.960 ;
      LAYER via ;
        RECT 738.400 927.900 738.660 928.160 ;
        RECT 742.540 927.900 742.800 928.160 ;
      LAYER met2 ;
        RECT 744.270 960.570 744.550 964.000 ;
        RECT 742.600 960.430 744.550 960.570 ;
        RECT 742.600 928.190 742.740 960.430 ;
        RECT 744.270 960.000 744.550 960.430 ;
        RECT 738.400 927.870 738.660 928.190 ;
        RECT 742.540 927.870 742.800 928.190 ;
        RECT 738.460 17.410 738.600 927.870 ;
        RECT 738.460 17.270 740.440 17.410 ;
        RECT 740.300 2.400 740.440 17.270 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1536.010 945.780 1536.330 945.840 ;
        RECT 1548.890 945.780 1549.210 945.840 ;
        RECT 1536.010 945.640 1549.210 945.780 ;
        RECT 1536.010 945.580 1536.330 945.640 ;
        RECT 1548.890 945.580 1549.210 945.640 ;
        RECT 1548.890 30.840 1549.210 30.900 ;
        RECT 1881.930 30.840 1882.250 30.900 ;
        RECT 1548.890 30.700 1882.250 30.840 ;
        RECT 1548.890 30.640 1549.210 30.700 ;
        RECT 1881.930 30.640 1882.250 30.700 ;
      LAYER via ;
        RECT 1536.040 945.580 1536.300 945.840 ;
        RECT 1548.920 945.580 1549.180 945.840 ;
        RECT 1548.920 30.640 1549.180 30.900 ;
        RECT 1881.960 30.640 1882.220 30.900 ;
      LAYER met2 ;
        RECT 1535.930 960.500 1536.210 964.000 ;
        RECT 1535.930 960.000 1536.240 960.500 ;
        RECT 1536.100 945.870 1536.240 960.000 ;
        RECT 1536.040 945.550 1536.300 945.870 ;
        RECT 1548.920 945.550 1549.180 945.870 ;
        RECT 1548.980 30.930 1549.120 945.550 ;
        RECT 1548.920 30.610 1549.180 30.930 ;
        RECT 1881.960 30.610 1882.220 30.930 ;
        RECT 1882.020 2.400 1882.160 30.610 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1548.430 948.500 1548.750 948.560 ;
        RECT 1552.110 948.500 1552.430 948.560 ;
        RECT 1548.430 948.360 1552.430 948.500 ;
        RECT 1548.430 948.300 1548.750 948.360 ;
        RECT 1552.110 948.300 1552.430 948.360 ;
        RECT 1552.110 93.060 1552.430 93.120 ;
        RECT 1897.570 93.060 1897.890 93.120 ;
        RECT 1552.110 92.920 1897.890 93.060 ;
        RECT 1552.110 92.860 1552.430 92.920 ;
        RECT 1897.570 92.860 1897.890 92.920 ;
        RECT 1897.570 2.960 1897.890 3.020 ;
        RECT 1899.870 2.960 1900.190 3.020 ;
        RECT 1897.570 2.820 1900.190 2.960 ;
        RECT 1897.570 2.760 1897.890 2.820 ;
        RECT 1899.870 2.760 1900.190 2.820 ;
      LAYER via ;
        RECT 1548.460 948.300 1548.720 948.560 ;
        RECT 1552.140 948.300 1552.400 948.560 ;
        RECT 1552.140 92.860 1552.400 93.120 ;
        RECT 1897.600 92.860 1897.860 93.120 ;
        RECT 1897.600 2.760 1897.860 3.020 ;
        RECT 1899.900 2.760 1900.160 3.020 ;
      LAYER met2 ;
        RECT 1548.350 960.500 1548.630 964.000 ;
        RECT 1548.350 960.000 1548.660 960.500 ;
        RECT 1548.520 948.590 1548.660 960.000 ;
        RECT 1548.460 948.270 1548.720 948.590 ;
        RECT 1552.140 948.270 1552.400 948.590 ;
        RECT 1552.200 93.150 1552.340 948.270 ;
        RECT 1552.140 92.830 1552.400 93.150 ;
        RECT 1897.600 92.830 1897.860 93.150 ;
        RECT 1897.660 3.050 1897.800 92.830 ;
        RECT 1897.600 2.730 1897.860 3.050 ;
        RECT 1899.900 2.730 1900.160 3.050 ;
        RECT 1899.960 2.400 1900.100 2.730 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.850 946.460 1561.170 946.520 ;
        RECT 1565.910 946.460 1566.230 946.520 ;
        RECT 1560.850 946.320 1566.230 946.460 ;
        RECT 1560.850 946.260 1561.170 946.320 ;
        RECT 1565.910 946.260 1566.230 946.320 ;
        RECT 1565.910 58.720 1566.230 58.780 ;
        RECT 1911.830 58.720 1912.150 58.780 ;
        RECT 1565.910 58.580 1912.150 58.720 ;
        RECT 1565.910 58.520 1566.230 58.580 ;
        RECT 1911.830 58.520 1912.150 58.580 ;
        RECT 1911.830 16.900 1912.150 16.960 ;
        RECT 1917.810 16.900 1918.130 16.960 ;
        RECT 1911.830 16.760 1918.130 16.900 ;
        RECT 1911.830 16.700 1912.150 16.760 ;
        RECT 1917.810 16.700 1918.130 16.760 ;
      LAYER via ;
        RECT 1560.880 946.260 1561.140 946.520 ;
        RECT 1565.940 946.260 1566.200 946.520 ;
        RECT 1565.940 58.520 1566.200 58.780 ;
        RECT 1911.860 58.520 1912.120 58.780 ;
        RECT 1911.860 16.700 1912.120 16.960 ;
        RECT 1917.840 16.700 1918.100 16.960 ;
      LAYER met2 ;
        RECT 1560.770 960.500 1561.050 964.000 ;
        RECT 1560.770 960.000 1561.080 960.500 ;
        RECT 1560.940 946.550 1561.080 960.000 ;
        RECT 1560.880 946.230 1561.140 946.550 ;
        RECT 1565.940 946.230 1566.200 946.550 ;
        RECT 1566.000 58.810 1566.140 946.230 ;
        RECT 1565.940 58.490 1566.200 58.810 ;
        RECT 1911.860 58.490 1912.120 58.810 ;
        RECT 1911.920 16.990 1912.060 58.490 ;
        RECT 1911.860 16.670 1912.120 16.990 ;
        RECT 1917.840 16.670 1918.100 16.990 ;
        RECT 1917.900 2.400 1918.040 16.670 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 162.080 1573.130 162.140 ;
        RECT 1932.070 162.080 1932.390 162.140 ;
        RECT 1572.810 161.940 1932.390 162.080 ;
        RECT 1572.810 161.880 1573.130 161.940 ;
        RECT 1932.070 161.880 1932.390 161.940 ;
      LAYER via ;
        RECT 1572.840 161.880 1573.100 162.140 ;
        RECT 1932.100 161.880 1932.360 162.140 ;
      LAYER met2 ;
        RECT 1572.730 960.500 1573.010 964.000 ;
        RECT 1572.730 960.000 1573.040 960.500 ;
        RECT 1572.900 162.170 1573.040 960.000 ;
        RECT 1572.840 161.850 1573.100 162.170 ;
        RECT 1932.100 161.850 1932.360 162.170 ;
        RECT 1932.160 17.410 1932.300 161.850 ;
        RECT 1932.160 17.270 1935.520 17.410 ;
        RECT 1935.380 2.400 1935.520 17.270 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1586.610 176.020 1586.930 176.080 ;
        RECT 1953.230 176.020 1953.550 176.080 ;
        RECT 1586.610 175.880 1953.550 176.020 ;
        RECT 1586.610 175.820 1586.930 175.880 ;
        RECT 1953.230 175.820 1953.550 175.880 ;
      LAYER via ;
        RECT 1586.640 175.820 1586.900 176.080 ;
        RECT 1953.260 175.820 1953.520 176.080 ;
      LAYER met2 ;
        RECT 1585.150 960.570 1585.430 964.000 ;
        RECT 1585.150 960.430 1586.840 960.570 ;
        RECT 1585.150 960.000 1585.430 960.430 ;
        RECT 1586.700 176.110 1586.840 960.430 ;
        RECT 1586.640 175.790 1586.900 176.110 ;
        RECT 1953.260 175.790 1953.520 176.110 ;
        RECT 1953.320 2.400 1953.460 175.790 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 51.580 1600.730 51.640 ;
        RECT 1966.570 51.580 1966.890 51.640 ;
        RECT 1600.410 51.440 1966.890 51.580 ;
        RECT 1600.410 51.380 1600.730 51.440 ;
        RECT 1966.570 51.380 1966.890 51.440 ;
      LAYER via ;
        RECT 1600.440 51.380 1600.700 51.640 ;
        RECT 1966.600 51.380 1966.860 51.640 ;
      LAYER met2 ;
        RECT 1597.570 960.570 1597.850 964.000 ;
        RECT 1597.570 960.430 1600.640 960.570 ;
        RECT 1597.570 960.000 1597.850 960.430 ;
        RECT 1600.500 51.670 1600.640 960.430 ;
        RECT 1600.440 51.350 1600.700 51.670 ;
        RECT 1966.600 51.350 1966.860 51.670 ;
        RECT 1966.660 17.410 1966.800 51.350 ;
        RECT 1966.660 17.270 1971.400 17.410 ;
        RECT 1971.260 2.400 1971.400 17.270 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1610.070 947.480 1610.390 947.540 ;
        RECT 1614.210 947.480 1614.530 947.540 ;
        RECT 1610.070 947.340 1614.530 947.480 ;
        RECT 1610.070 947.280 1610.390 947.340 ;
        RECT 1614.210 947.280 1614.530 947.340 ;
        RECT 1614.210 79.460 1614.530 79.520 ;
        RECT 1987.270 79.460 1987.590 79.520 ;
        RECT 1614.210 79.320 1987.590 79.460 ;
        RECT 1614.210 79.260 1614.530 79.320 ;
        RECT 1987.270 79.260 1987.590 79.320 ;
      LAYER via ;
        RECT 1610.100 947.280 1610.360 947.540 ;
        RECT 1614.240 947.280 1614.500 947.540 ;
        RECT 1614.240 79.260 1614.500 79.520 ;
        RECT 1987.300 79.260 1987.560 79.520 ;
      LAYER met2 ;
        RECT 1609.990 960.500 1610.270 964.000 ;
        RECT 1609.990 960.000 1610.300 960.500 ;
        RECT 1610.160 947.570 1610.300 960.000 ;
        RECT 1610.100 947.250 1610.360 947.570 ;
        RECT 1614.240 947.250 1614.500 947.570 ;
        RECT 1614.300 79.550 1614.440 947.250 ;
        RECT 1614.240 79.230 1614.500 79.550 ;
        RECT 1987.300 79.230 1987.560 79.550 ;
        RECT 1987.360 17.410 1987.500 79.230 ;
        RECT 1987.360 17.270 1989.340 17.410 ;
        RECT 1989.200 2.400 1989.340 17.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1622.490 945.440 1622.810 945.500 ;
        RECT 1638.590 945.440 1638.910 945.500 ;
        RECT 1622.490 945.300 1638.910 945.440 ;
        RECT 1622.490 945.240 1622.810 945.300 ;
        RECT 1638.590 945.240 1638.910 945.300 ;
        RECT 1638.590 44.780 1638.910 44.840 ;
        RECT 2006.590 44.780 2006.910 44.840 ;
        RECT 1638.590 44.640 2006.910 44.780 ;
        RECT 1638.590 44.580 1638.910 44.640 ;
        RECT 2006.590 44.580 2006.910 44.640 ;
      LAYER via ;
        RECT 1622.520 945.240 1622.780 945.500 ;
        RECT 1638.620 945.240 1638.880 945.500 ;
        RECT 1638.620 44.580 1638.880 44.840 ;
        RECT 2006.620 44.580 2006.880 44.840 ;
      LAYER met2 ;
        RECT 1622.410 960.500 1622.690 964.000 ;
        RECT 1622.410 960.000 1622.720 960.500 ;
        RECT 1622.580 945.530 1622.720 960.000 ;
        RECT 1622.520 945.210 1622.780 945.530 ;
        RECT 1638.620 945.210 1638.880 945.530 ;
        RECT 1638.680 44.870 1638.820 945.210 ;
        RECT 1638.620 44.550 1638.880 44.870 ;
        RECT 2006.620 44.550 2006.880 44.870 ;
        RECT 2006.680 2.400 2006.820 44.550 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.910 99.860 1635.230 99.920 ;
        RECT 2021.770 99.860 2022.090 99.920 ;
        RECT 1634.910 99.720 2022.090 99.860 ;
        RECT 1634.910 99.660 1635.230 99.720 ;
        RECT 2021.770 99.660 2022.090 99.720 ;
      LAYER via ;
        RECT 1634.940 99.660 1635.200 99.920 ;
        RECT 2021.800 99.660 2022.060 99.920 ;
      LAYER met2 ;
        RECT 1634.830 960.500 1635.110 964.000 ;
        RECT 1634.830 960.000 1635.140 960.500 ;
        RECT 1635.000 99.950 1635.140 960.000 ;
        RECT 1634.940 99.630 1635.200 99.950 ;
        RECT 2021.800 99.630 2022.060 99.950 ;
        RECT 2021.860 17.410 2022.000 99.630 ;
        RECT 2021.860 17.270 2024.760 17.410 ;
        RECT 2024.620 2.400 2024.760 17.270 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1647.330 949.860 1647.650 949.920 ;
        RECT 1659.290 949.860 1659.610 949.920 ;
        RECT 1647.330 949.720 1659.610 949.860 ;
        RECT 1647.330 949.660 1647.650 949.720 ;
        RECT 1659.290 949.660 1659.610 949.720 ;
        RECT 1659.290 520.780 1659.610 520.840 ;
        RECT 2042.470 520.780 2042.790 520.840 ;
        RECT 1659.290 520.640 2042.790 520.780 ;
        RECT 1659.290 520.580 1659.610 520.640 ;
        RECT 2042.470 520.580 2042.790 520.640 ;
      LAYER via ;
        RECT 1647.360 949.660 1647.620 949.920 ;
        RECT 1659.320 949.660 1659.580 949.920 ;
        RECT 1659.320 520.580 1659.580 520.840 ;
        RECT 2042.500 520.580 2042.760 520.840 ;
      LAYER met2 ;
        RECT 1647.250 960.500 1647.530 964.000 ;
        RECT 1647.250 960.000 1647.560 960.500 ;
        RECT 1647.420 949.950 1647.560 960.000 ;
        RECT 1647.360 949.630 1647.620 949.950 ;
        RECT 1659.320 949.630 1659.580 949.950 ;
        RECT 1659.380 520.870 1659.520 949.630 ;
        RECT 1659.320 520.550 1659.580 520.870 ;
        RECT 2042.500 520.550 2042.760 520.870 ;
        RECT 2042.560 2.400 2042.700 520.550 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.170 928.100 752.490 928.160 ;
        RECT 755.390 928.100 755.710 928.160 ;
        RECT 752.170 927.960 755.710 928.100 ;
        RECT 752.170 927.900 752.490 927.960 ;
        RECT 755.390 927.900 755.710 927.960 ;
        RECT 752.170 17.920 752.490 17.980 ;
        RECT 757.690 17.920 758.010 17.980 ;
        RECT 752.170 17.780 758.010 17.920 ;
        RECT 752.170 17.720 752.490 17.780 ;
        RECT 757.690 17.720 758.010 17.780 ;
      LAYER via ;
        RECT 752.200 927.900 752.460 928.160 ;
        RECT 755.420 927.900 755.680 928.160 ;
        RECT 752.200 17.720 752.460 17.980 ;
        RECT 757.720 17.720 757.980 17.980 ;
      LAYER met2 ;
        RECT 756.690 960.570 756.970 964.000 ;
        RECT 755.480 960.430 756.970 960.570 ;
        RECT 755.480 928.190 755.620 960.430 ;
        RECT 756.690 960.000 756.970 960.430 ;
        RECT 752.200 927.870 752.460 928.190 ;
        RECT 755.420 927.870 755.680 928.190 ;
        RECT 752.260 18.010 752.400 927.870 ;
        RECT 752.200 17.690 752.460 18.010 ;
        RECT 757.720 17.690 757.980 18.010 ;
        RECT 757.780 2.400 757.920 17.690 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 107.000 1662.830 107.060 ;
        RECT 2056.270 107.000 2056.590 107.060 ;
        RECT 1662.510 106.860 2056.590 107.000 ;
        RECT 1662.510 106.800 1662.830 106.860 ;
        RECT 2056.270 106.800 2056.590 106.860 ;
      LAYER via ;
        RECT 1662.540 106.800 1662.800 107.060 ;
        RECT 2056.300 106.800 2056.560 107.060 ;
      LAYER met2 ;
        RECT 1659.670 960.570 1659.950 964.000 ;
        RECT 1659.670 960.430 1662.740 960.570 ;
        RECT 1659.670 960.000 1659.950 960.430 ;
        RECT 1662.600 107.090 1662.740 960.430 ;
        RECT 1662.540 106.770 1662.800 107.090 ;
        RECT 2056.300 106.770 2056.560 107.090 ;
        RECT 2056.360 17.410 2056.500 106.770 ;
        RECT 2056.360 17.270 2060.640 17.410 ;
        RECT 2060.500 2.400 2060.640 17.270 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1675.850 886.620 1676.170 886.680 ;
        RECT 2076.970 886.620 2077.290 886.680 ;
        RECT 1675.850 886.480 2077.290 886.620 ;
        RECT 1675.850 886.420 1676.170 886.480 ;
        RECT 2076.970 886.420 2077.290 886.480 ;
      LAYER via ;
        RECT 1675.880 886.420 1676.140 886.680 ;
        RECT 2077.000 886.420 2077.260 886.680 ;
      LAYER met2 ;
        RECT 1672.090 960.570 1672.370 964.000 ;
        RECT 1672.090 960.430 1676.080 960.570 ;
        RECT 1672.090 960.000 1672.370 960.430 ;
        RECT 1675.940 886.710 1676.080 960.430 ;
        RECT 1675.880 886.390 1676.140 886.710 ;
        RECT 2077.000 886.390 2077.260 886.710 ;
        RECT 2077.060 17.410 2077.200 886.390 ;
        RECT 2077.060 17.270 2078.580 17.410 ;
        RECT 2078.440 2.400 2078.580 17.270 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1684.590 946.460 1684.910 946.520 ;
        RECT 1690.110 946.460 1690.430 946.520 ;
        RECT 1684.590 946.320 1690.430 946.460 ;
        RECT 1684.590 946.260 1684.910 946.320 ;
        RECT 1690.110 946.260 1690.430 946.320 ;
        RECT 1690.110 113.800 1690.430 113.860 ;
        RECT 2090.770 113.800 2091.090 113.860 ;
        RECT 1690.110 113.660 2091.090 113.800 ;
        RECT 1690.110 113.600 1690.430 113.660 ;
        RECT 2090.770 113.600 2091.090 113.660 ;
      LAYER via ;
        RECT 1684.620 946.260 1684.880 946.520 ;
        RECT 1690.140 946.260 1690.400 946.520 ;
        RECT 1690.140 113.600 1690.400 113.860 ;
        RECT 2090.800 113.600 2091.060 113.860 ;
      LAYER met2 ;
        RECT 1684.510 960.500 1684.790 964.000 ;
        RECT 1684.510 960.000 1684.820 960.500 ;
        RECT 1684.680 946.550 1684.820 960.000 ;
        RECT 1684.620 946.230 1684.880 946.550 ;
        RECT 1690.140 946.230 1690.400 946.550 ;
        RECT 1690.200 113.890 1690.340 946.230 ;
        RECT 1690.140 113.570 1690.400 113.890 ;
        RECT 2090.800 113.570 2091.060 113.890 ;
        RECT 2090.860 17.410 2091.000 113.570 ;
        RECT 2090.860 17.270 2096.060 17.410 ;
        RECT 2095.920 2.400 2096.060 17.270 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.010 120.940 1697.330 121.000 ;
        RECT 2111.470 120.940 2111.790 121.000 ;
        RECT 1697.010 120.800 2111.790 120.940 ;
        RECT 1697.010 120.740 1697.330 120.800 ;
        RECT 2111.470 120.740 2111.790 120.800 ;
      LAYER via ;
        RECT 1697.040 120.740 1697.300 121.000 ;
        RECT 2111.500 120.740 2111.760 121.000 ;
      LAYER met2 ;
        RECT 1696.470 960.570 1696.750 964.000 ;
        RECT 1696.470 960.430 1697.240 960.570 ;
        RECT 1696.470 960.000 1696.750 960.430 ;
        RECT 1697.100 121.030 1697.240 960.430 ;
        RECT 1697.040 120.710 1697.300 121.030 ;
        RECT 2111.500 120.710 2111.760 121.030 ;
        RECT 2111.560 17.410 2111.700 120.710 ;
        RECT 2111.560 17.270 2114.000 17.410 ;
        RECT 2113.860 2.400 2114.000 17.270 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 189.620 1711.130 189.680 ;
        RECT 2125.730 189.620 2126.050 189.680 ;
        RECT 1710.810 189.480 2126.050 189.620 ;
        RECT 1710.810 189.420 1711.130 189.480 ;
        RECT 2125.730 189.420 2126.050 189.480 ;
        RECT 2125.730 20.980 2126.050 21.040 ;
        RECT 2131.710 20.980 2132.030 21.040 ;
        RECT 2125.730 20.840 2132.030 20.980 ;
        RECT 2125.730 20.780 2126.050 20.840 ;
        RECT 2131.710 20.780 2132.030 20.840 ;
      LAYER via ;
        RECT 1710.840 189.420 1711.100 189.680 ;
        RECT 2125.760 189.420 2126.020 189.680 ;
        RECT 2125.760 20.780 2126.020 21.040 ;
        RECT 2131.740 20.780 2132.000 21.040 ;
      LAYER met2 ;
        RECT 1708.890 960.570 1709.170 964.000 ;
        RECT 1708.890 960.430 1711.040 960.570 ;
        RECT 1708.890 960.000 1709.170 960.430 ;
        RECT 1710.900 189.710 1711.040 960.430 ;
        RECT 1710.840 189.390 1711.100 189.710 ;
        RECT 2125.760 189.390 2126.020 189.710 ;
        RECT 2125.820 21.070 2125.960 189.390 ;
        RECT 2125.760 20.750 2126.020 21.070 ;
        RECT 2131.740 20.750 2132.000 21.070 ;
        RECT 2131.800 2.400 2131.940 20.750 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 72.320 1724.930 72.380 ;
        RECT 2145.970 72.320 2146.290 72.380 ;
        RECT 1724.610 72.180 2146.290 72.320 ;
        RECT 1724.610 72.120 1724.930 72.180 ;
        RECT 2145.970 72.120 2146.290 72.180 ;
      LAYER via ;
        RECT 1724.640 72.120 1724.900 72.380 ;
        RECT 2146.000 72.120 2146.260 72.380 ;
      LAYER met2 ;
        RECT 1721.310 960.570 1721.590 964.000 ;
        RECT 1721.310 960.430 1724.840 960.570 ;
        RECT 1721.310 960.000 1721.590 960.430 ;
        RECT 1724.700 72.410 1724.840 960.430 ;
        RECT 1724.640 72.090 1724.900 72.410 ;
        RECT 2146.000 72.090 2146.260 72.410 ;
        RECT 2146.060 17.410 2146.200 72.090 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1733.810 945.440 1734.130 945.500 ;
        RECT 1742.090 945.440 1742.410 945.500 ;
        RECT 1733.810 945.300 1742.410 945.440 ;
        RECT 1733.810 945.240 1734.130 945.300 ;
        RECT 1742.090 945.240 1742.410 945.300 ;
        RECT 1742.090 155.280 1742.410 155.340 ;
        RECT 2167.130 155.280 2167.450 155.340 ;
        RECT 1742.090 155.140 2167.450 155.280 ;
        RECT 1742.090 155.080 1742.410 155.140 ;
        RECT 2167.130 155.080 2167.450 155.140 ;
      LAYER via ;
        RECT 1733.840 945.240 1734.100 945.500 ;
        RECT 1742.120 945.240 1742.380 945.500 ;
        RECT 1742.120 155.080 1742.380 155.340 ;
        RECT 2167.160 155.080 2167.420 155.340 ;
      LAYER met2 ;
        RECT 1733.730 960.500 1734.010 964.000 ;
        RECT 1733.730 960.000 1734.040 960.500 ;
        RECT 1733.900 945.530 1734.040 960.000 ;
        RECT 1733.840 945.210 1734.100 945.530 ;
        RECT 1742.120 945.210 1742.380 945.530 ;
        RECT 1742.180 155.370 1742.320 945.210 ;
        RECT 1742.120 155.050 1742.380 155.370 ;
        RECT 2167.160 155.050 2167.420 155.370 ;
        RECT 2167.220 17.410 2167.360 155.050 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1746.230 949.180 1746.550 949.240 ;
        RECT 1921.490 949.180 1921.810 949.240 ;
        RECT 1746.230 949.040 1921.810 949.180 ;
        RECT 1746.230 948.980 1746.550 949.040 ;
        RECT 1921.490 948.980 1921.810 949.040 ;
        RECT 1921.490 86.260 1921.810 86.320 ;
        RECT 2180.470 86.260 2180.790 86.320 ;
        RECT 1921.490 86.120 2180.790 86.260 ;
        RECT 1921.490 86.060 1921.810 86.120 ;
        RECT 2180.470 86.060 2180.790 86.120 ;
      LAYER via ;
        RECT 1746.260 948.980 1746.520 949.240 ;
        RECT 1921.520 948.980 1921.780 949.240 ;
        RECT 1921.520 86.060 1921.780 86.320 ;
        RECT 2180.500 86.060 2180.760 86.320 ;
      LAYER met2 ;
        RECT 1746.150 960.500 1746.430 964.000 ;
        RECT 1746.150 960.000 1746.460 960.500 ;
        RECT 1746.320 949.270 1746.460 960.000 ;
        RECT 1746.260 948.950 1746.520 949.270 ;
        RECT 1921.520 948.950 1921.780 949.270 ;
        RECT 1921.580 86.350 1921.720 948.950 ;
        RECT 1921.520 86.030 1921.780 86.350 ;
        RECT 2180.500 86.030 2180.760 86.350 ;
        RECT 2180.560 17.410 2180.700 86.030 ;
        RECT 2180.560 17.270 2185.300 17.410 ;
        RECT 2185.160 2.400 2185.300 17.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 168.880 1759.430 168.940 ;
        RECT 2201.170 168.880 2201.490 168.940 ;
        RECT 1759.110 168.740 2201.490 168.880 ;
        RECT 1759.110 168.680 1759.430 168.740 ;
        RECT 2201.170 168.680 2201.490 168.740 ;
      LAYER via ;
        RECT 1759.140 168.680 1759.400 168.940 ;
        RECT 2201.200 168.680 2201.460 168.940 ;
      LAYER met2 ;
        RECT 1758.570 960.570 1758.850 964.000 ;
        RECT 1758.570 960.430 1759.340 960.570 ;
        RECT 1758.570 960.000 1758.850 960.430 ;
        RECT 1759.200 168.970 1759.340 960.430 ;
        RECT 1759.140 168.650 1759.400 168.970 ;
        RECT 2201.200 168.650 2201.460 168.970 ;
        RECT 2201.260 17.410 2201.400 168.650 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 203.560 1773.230 203.620 ;
        RECT 2215.430 203.560 2215.750 203.620 ;
        RECT 1772.910 203.420 2215.750 203.560 ;
        RECT 1772.910 203.360 1773.230 203.420 ;
        RECT 2215.430 203.360 2215.750 203.420 ;
      LAYER via ;
        RECT 1772.940 203.360 1773.200 203.620 ;
        RECT 2215.460 203.360 2215.720 203.620 ;
      LAYER met2 ;
        RECT 1770.990 960.570 1771.270 964.000 ;
        RECT 1770.990 960.430 1773.140 960.570 ;
        RECT 1770.990 960.000 1771.270 960.430 ;
        RECT 1773.000 203.650 1773.140 960.430 ;
        RECT 1772.940 203.330 1773.200 203.650 ;
        RECT 2215.460 203.330 2215.720 203.650 ;
        RECT 2215.520 16.730 2215.660 203.330 ;
        RECT 2215.520 16.590 2221.180 16.730 ;
        RECT 2221.040 2.400 2221.180 16.590 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 17.240 772.730 17.300 ;
        RECT 775.630 17.240 775.950 17.300 ;
        RECT 772.410 17.100 775.950 17.240 ;
        RECT 772.410 17.040 772.730 17.100 ;
        RECT 775.630 17.040 775.950 17.100 ;
      LAYER via ;
        RECT 772.440 17.040 772.700 17.300 ;
        RECT 775.660 17.040 775.920 17.300 ;
      LAYER met2 ;
        RECT 769.110 960.570 769.390 964.000 ;
        RECT 769.110 960.430 772.640 960.570 ;
        RECT 769.110 960.000 769.390 960.430 ;
        RECT 772.500 17.330 772.640 960.430 ;
        RECT 772.440 17.010 772.700 17.330 ;
        RECT 775.660 17.010 775.920 17.330 ;
        RECT 775.720 2.400 775.860 17.010 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 182.820 1787.030 182.880 ;
        RECT 2235.670 182.820 2235.990 182.880 ;
        RECT 1786.710 182.680 2235.990 182.820 ;
        RECT 1786.710 182.620 1787.030 182.680 ;
        RECT 2235.670 182.620 2235.990 182.680 ;
      LAYER via ;
        RECT 1786.740 182.620 1787.000 182.880 ;
        RECT 2235.700 182.620 2235.960 182.880 ;
      LAYER met2 ;
        RECT 1783.410 960.570 1783.690 964.000 ;
        RECT 1783.410 960.430 1786.940 960.570 ;
        RECT 1783.410 960.000 1783.690 960.430 ;
        RECT 1786.800 182.910 1786.940 960.430 ;
        RECT 1786.740 182.590 1787.000 182.910 ;
        RECT 2235.700 182.590 2235.960 182.910 ;
        RECT 2235.760 16.730 2235.900 182.590 ;
        RECT 2235.760 16.590 2239.120 16.730 ;
        RECT 2238.980 2.400 2239.120 16.590 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1795.910 945.440 1796.230 945.500 ;
        RECT 1800.510 945.440 1800.830 945.500 ;
        RECT 1795.910 945.300 1800.830 945.440 ;
        RECT 1795.910 945.240 1796.230 945.300 ;
        RECT 1800.510 945.240 1800.830 945.300 ;
        RECT 1800.510 217.160 1800.830 217.220 ;
        RECT 2256.830 217.160 2257.150 217.220 ;
        RECT 1800.510 217.020 2257.150 217.160 ;
        RECT 1800.510 216.960 1800.830 217.020 ;
        RECT 2256.830 216.960 2257.150 217.020 ;
      LAYER via ;
        RECT 1795.940 945.240 1796.200 945.500 ;
        RECT 1800.540 945.240 1800.800 945.500 ;
        RECT 1800.540 216.960 1800.800 217.220 ;
        RECT 2256.860 216.960 2257.120 217.220 ;
      LAYER met2 ;
        RECT 1795.830 960.500 1796.110 964.000 ;
        RECT 1795.830 960.000 1796.140 960.500 ;
        RECT 1796.000 945.530 1796.140 960.000 ;
        RECT 1795.940 945.210 1796.200 945.530 ;
        RECT 1800.540 945.210 1800.800 945.530 ;
        RECT 1800.600 217.250 1800.740 945.210 ;
        RECT 1800.540 216.930 1800.800 217.250 ;
        RECT 2256.860 216.930 2257.120 217.250 ;
        RECT 2256.920 17.410 2257.060 216.930 ;
        RECT 2256.460 17.270 2257.060 17.410 ;
        RECT 2256.460 2.400 2256.600 17.270 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.870 945.440 1808.190 945.500 ;
        RECT 1814.310 945.440 1814.630 945.500 ;
        RECT 1807.870 945.300 1814.630 945.440 ;
        RECT 1807.870 945.240 1808.190 945.300 ;
        RECT 1814.310 945.240 1814.630 945.300 ;
        RECT 1814.310 196.760 1814.630 196.820 ;
        RECT 2270.170 196.760 2270.490 196.820 ;
        RECT 1814.310 196.620 2270.490 196.760 ;
        RECT 1814.310 196.560 1814.630 196.620 ;
        RECT 2270.170 196.560 2270.490 196.620 ;
      LAYER via ;
        RECT 1807.900 945.240 1808.160 945.500 ;
        RECT 1814.340 945.240 1814.600 945.500 ;
        RECT 1814.340 196.560 1814.600 196.820 ;
        RECT 2270.200 196.560 2270.460 196.820 ;
      LAYER met2 ;
        RECT 1807.790 960.500 1808.070 964.000 ;
        RECT 1807.790 960.000 1808.100 960.500 ;
        RECT 1807.960 945.530 1808.100 960.000 ;
        RECT 1807.900 945.210 1808.160 945.530 ;
        RECT 1814.340 945.210 1814.600 945.530 ;
        RECT 1814.400 196.850 1814.540 945.210 ;
        RECT 1814.340 196.530 1814.600 196.850 ;
        RECT 2270.200 196.530 2270.460 196.850 ;
        RECT 2270.260 17.410 2270.400 196.530 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1820.750 817.600 1821.070 817.660 ;
        RECT 2290.870 817.600 2291.190 817.660 ;
        RECT 1820.750 817.460 2291.190 817.600 ;
        RECT 1820.750 817.400 1821.070 817.460 ;
        RECT 2290.870 817.400 2291.190 817.460 ;
      LAYER via ;
        RECT 1820.780 817.400 1821.040 817.660 ;
        RECT 2290.900 817.400 2291.160 817.660 ;
      LAYER met2 ;
        RECT 1820.210 960.570 1820.490 964.000 ;
        RECT 1820.210 960.430 1820.980 960.570 ;
        RECT 1820.210 960.000 1820.490 960.430 ;
        RECT 1820.840 817.690 1820.980 960.430 ;
        RECT 1820.780 817.370 1821.040 817.690 ;
        RECT 2290.900 817.370 2291.160 817.690 ;
        RECT 2290.960 17.410 2291.100 817.370 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1834.550 810.800 1834.870 810.860 ;
        RECT 2304.670 810.800 2304.990 810.860 ;
        RECT 1834.550 810.660 2304.990 810.800 ;
        RECT 1834.550 810.600 1834.870 810.660 ;
        RECT 2304.670 810.600 2304.990 810.660 ;
      LAYER via ;
        RECT 1834.580 810.600 1834.840 810.860 ;
        RECT 2304.700 810.600 2304.960 810.860 ;
      LAYER met2 ;
        RECT 1832.630 960.570 1832.910 964.000 ;
        RECT 1832.630 960.430 1834.780 960.570 ;
        RECT 1832.630 960.000 1832.910 960.430 ;
        RECT 1834.640 810.890 1834.780 960.430 ;
        RECT 1834.580 810.570 1834.840 810.890 ;
        RECT 2304.700 810.570 2304.960 810.890 ;
        RECT 2304.760 17.410 2304.900 810.570 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.810 141.340 1849.130 141.400 ;
        RECT 2325.370 141.340 2325.690 141.400 ;
        RECT 1848.810 141.200 2325.690 141.340 ;
        RECT 1848.810 141.140 1849.130 141.200 ;
        RECT 2325.370 141.140 2325.690 141.200 ;
      LAYER via ;
        RECT 1848.840 141.140 1849.100 141.400 ;
        RECT 2325.400 141.140 2325.660 141.400 ;
      LAYER met2 ;
        RECT 1845.050 960.570 1845.330 964.000 ;
        RECT 1845.050 960.430 1849.040 960.570 ;
        RECT 1845.050 960.000 1845.330 960.430 ;
        RECT 1848.900 141.430 1849.040 960.430 ;
        RECT 1848.840 141.110 1849.100 141.430 ;
        RECT 2325.400 141.110 2325.660 141.430 ;
        RECT 2325.460 17.410 2325.600 141.110 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1857.550 946.800 1857.870 946.860 ;
        RECT 1862.610 946.800 1862.930 946.860 ;
        RECT 1857.550 946.660 1862.930 946.800 ;
        RECT 1857.550 946.600 1857.870 946.660 ;
        RECT 1862.610 946.600 1862.930 946.660 ;
        RECT 1862.610 134.540 1862.930 134.600 ;
        RECT 2339.630 134.540 2339.950 134.600 ;
        RECT 1862.610 134.400 2339.950 134.540 ;
        RECT 1862.610 134.340 1862.930 134.400 ;
        RECT 2339.630 134.340 2339.950 134.400 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.610 16.900 2345.930 16.960 ;
        RECT 2339.630 16.760 2345.930 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.610 16.700 2345.930 16.760 ;
      LAYER via ;
        RECT 1857.580 946.600 1857.840 946.860 ;
        RECT 1862.640 946.600 1862.900 946.860 ;
        RECT 1862.640 134.340 1862.900 134.600 ;
        RECT 2339.660 134.340 2339.920 134.600 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.640 16.700 2345.900 16.960 ;
      LAYER met2 ;
        RECT 1857.470 960.500 1857.750 964.000 ;
        RECT 1857.470 960.000 1857.780 960.500 ;
        RECT 1857.640 946.890 1857.780 960.000 ;
        RECT 1857.580 946.570 1857.840 946.890 ;
        RECT 1862.640 946.570 1862.900 946.890 ;
        RECT 1862.700 134.630 1862.840 946.570 ;
        RECT 1862.640 134.310 1862.900 134.630 ;
        RECT 2339.660 134.310 2339.920 134.630 ;
        RECT 2339.720 16.990 2339.860 134.310 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.640 16.670 2345.900 16.990 ;
        RECT 2345.700 2.400 2345.840 16.670 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.970 946.460 1870.290 946.520 ;
        RECT 1876.410 946.460 1876.730 946.520 ;
        RECT 1869.970 946.320 1876.730 946.460 ;
        RECT 1869.970 946.260 1870.290 946.320 ;
        RECT 1876.410 946.260 1876.730 946.320 ;
        RECT 1876.410 231.100 1876.730 231.160 ;
        RECT 2359.870 231.100 2360.190 231.160 ;
        RECT 1876.410 230.960 2360.190 231.100 ;
        RECT 1876.410 230.900 1876.730 230.960 ;
        RECT 2359.870 230.900 2360.190 230.960 ;
      LAYER via ;
        RECT 1870.000 946.260 1870.260 946.520 ;
        RECT 1876.440 946.260 1876.700 946.520 ;
        RECT 1876.440 230.900 1876.700 231.160 ;
        RECT 2359.900 230.900 2360.160 231.160 ;
      LAYER met2 ;
        RECT 1869.890 960.500 1870.170 964.000 ;
        RECT 1869.890 960.000 1870.200 960.500 ;
        RECT 1870.060 946.550 1870.200 960.000 ;
        RECT 1870.000 946.230 1870.260 946.550 ;
        RECT 1876.440 946.230 1876.700 946.550 ;
        RECT 1876.500 231.190 1876.640 946.230 ;
        RECT 1876.440 230.870 1876.700 231.190 ;
        RECT 2359.900 230.870 2360.160 231.190 ;
        RECT 2359.960 17.410 2360.100 230.870 ;
        RECT 2359.960 17.270 2363.780 17.410 ;
        RECT 2363.640 2.400 2363.780 17.270 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1882.850 803.660 1883.170 803.720 ;
        RECT 2380.570 803.660 2380.890 803.720 ;
        RECT 1882.850 803.520 2380.890 803.660 ;
        RECT 1882.850 803.460 1883.170 803.520 ;
        RECT 2380.570 803.460 2380.890 803.520 ;
      LAYER via ;
        RECT 1882.880 803.460 1883.140 803.720 ;
        RECT 2380.600 803.460 2380.860 803.720 ;
      LAYER met2 ;
        RECT 1882.310 960.570 1882.590 964.000 ;
        RECT 1882.310 960.430 1883.080 960.570 ;
        RECT 1882.310 960.000 1882.590 960.430 ;
        RECT 1882.940 803.750 1883.080 960.430 ;
        RECT 1882.880 803.430 1883.140 803.750 ;
        RECT 2380.600 803.430 2380.860 803.750 ;
        RECT 2380.660 17.410 2380.800 803.430 ;
        RECT 2380.660 17.270 2381.720 17.410 ;
        RECT 2381.580 2.400 2381.720 17.270 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1894.810 945.780 1895.130 945.840 ;
        RECT 1907.690 945.780 1908.010 945.840 ;
        RECT 1894.810 945.640 1908.010 945.780 ;
        RECT 1894.810 945.580 1895.130 945.640 ;
        RECT 1907.690 945.580 1908.010 945.640 ;
        RECT 1907.690 796.860 1908.010 796.920 ;
        RECT 2394.370 796.860 2394.690 796.920 ;
        RECT 1907.690 796.720 2394.690 796.860 ;
        RECT 1907.690 796.660 1908.010 796.720 ;
        RECT 2394.370 796.660 2394.690 796.720 ;
      LAYER via ;
        RECT 1894.840 945.580 1895.100 945.840 ;
        RECT 1907.720 945.580 1907.980 945.840 ;
        RECT 1907.720 796.660 1907.980 796.920 ;
        RECT 2394.400 796.660 2394.660 796.920 ;
      LAYER met2 ;
        RECT 1894.730 960.500 1895.010 964.000 ;
        RECT 1894.730 960.000 1895.040 960.500 ;
        RECT 1894.900 945.870 1895.040 960.000 ;
        RECT 1894.840 945.550 1895.100 945.870 ;
        RECT 1907.720 945.550 1907.980 945.870 ;
        RECT 1907.780 796.950 1907.920 945.550 ;
        RECT 1907.720 796.630 1907.980 796.950 ;
        RECT 2394.400 796.630 2394.660 796.950 ;
        RECT 2394.460 17.410 2394.600 796.630 ;
        RECT 2394.460 17.270 2399.660 17.410 ;
        RECT 2399.520 2.400 2399.660 17.270 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 781.150 946.800 781.470 946.860 ;
        RECT 786.210 946.800 786.530 946.860 ;
        RECT 781.150 946.660 786.530 946.800 ;
        RECT 781.150 946.600 781.470 946.660 ;
        RECT 786.210 946.600 786.530 946.660 ;
        RECT 786.210 17.580 786.530 17.640 ;
        RECT 793.570 17.580 793.890 17.640 ;
        RECT 786.210 17.440 793.890 17.580 ;
        RECT 786.210 17.380 786.530 17.440 ;
        RECT 793.570 17.380 793.890 17.440 ;
      LAYER via ;
        RECT 781.180 946.600 781.440 946.860 ;
        RECT 786.240 946.600 786.500 946.860 ;
        RECT 786.240 17.380 786.500 17.640 ;
        RECT 793.600 17.380 793.860 17.640 ;
      LAYER met2 ;
        RECT 781.070 960.500 781.350 964.000 ;
        RECT 781.070 960.000 781.380 960.500 ;
        RECT 781.240 946.890 781.380 960.000 ;
        RECT 781.180 946.570 781.440 946.890 ;
        RECT 786.240 946.570 786.500 946.890 ;
        RECT 786.300 17.670 786.440 946.570 ;
        RECT 786.240 17.350 786.500 17.670 ;
        RECT 793.600 17.350 793.860 17.670 ;
        RECT 793.660 2.400 793.800 17.350 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 20.640 639.330 20.700 ;
        RECT 670.750 20.640 671.070 20.700 ;
        RECT 639.010 20.500 671.070 20.640 ;
        RECT 639.010 20.440 639.330 20.500 ;
        RECT 670.750 20.440 671.070 20.500 ;
      LAYER via ;
        RECT 639.040 20.440 639.300 20.700 ;
        RECT 670.780 20.440 671.040 20.700 ;
      LAYER met2 ;
        RECT 673.890 960.570 674.170 964.000 ;
        RECT 670.840 960.430 674.170 960.570 ;
        RECT 670.840 20.730 670.980 960.430 ;
        RECT 673.890 960.000 674.170 960.430 ;
        RECT 639.040 20.410 639.300 20.730 ;
        RECT 670.780 20.410 671.040 20.730 ;
        RECT 639.100 2.400 639.240 20.410 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1911.370 949.520 1911.690 949.580 ;
        RECT 1935.290 949.520 1935.610 949.580 ;
        RECT 1911.370 949.380 1935.610 949.520 ;
        RECT 1911.370 949.320 1911.690 949.380 ;
        RECT 1935.290 949.320 1935.610 949.380 ;
        RECT 1935.290 783.260 1935.610 783.320 ;
        RECT 2421.970 783.260 2422.290 783.320 ;
        RECT 1935.290 783.120 2422.290 783.260 ;
        RECT 1935.290 783.060 1935.610 783.120 ;
        RECT 2421.970 783.060 2422.290 783.120 ;
      LAYER via ;
        RECT 1911.400 949.320 1911.660 949.580 ;
        RECT 1935.320 949.320 1935.580 949.580 ;
        RECT 1935.320 783.060 1935.580 783.320 ;
        RECT 2422.000 783.060 2422.260 783.320 ;
      LAYER met2 ;
        RECT 1911.290 960.500 1911.570 964.000 ;
        RECT 1911.290 960.000 1911.600 960.500 ;
        RECT 1911.460 949.610 1911.600 960.000 ;
        RECT 1911.400 949.290 1911.660 949.610 ;
        RECT 1935.320 949.290 1935.580 949.610 ;
        RECT 1935.380 783.350 1935.520 949.290 ;
        RECT 1935.320 783.030 1935.580 783.350 ;
        RECT 2422.000 783.030 2422.260 783.350 ;
        RECT 2422.060 17.410 2422.200 783.030 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 776.120 1925.030 776.180 ;
        RECT 2435.770 776.120 2436.090 776.180 ;
        RECT 1924.710 775.980 2436.090 776.120 ;
        RECT 1924.710 775.920 1925.030 775.980 ;
        RECT 2435.770 775.920 2436.090 775.980 ;
      LAYER via ;
        RECT 1924.740 775.920 1925.000 776.180 ;
        RECT 2435.800 775.920 2436.060 776.180 ;
      LAYER met2 ;
        RECT 1923.250 960.570 1923.530 964.000 ;
        RECT 1923.250 960.430 1924.940 960.570 ;
        RECT 1923.250 960.000 1923.530 960.430 ;
        RECT 1924.800 776.210 1924.940 960.430 ;
        RECT 1924.740 775.890 1925.000 776.210 ;
        RECT 2435.800 775.890 2436.060 776.210 ;
        RECT 2435.860 17.410 2436.000 775.890 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1938.510 162.080 1938.830 162.140 ;
        RECT 2456.470 162.080 2456.790 162.140 ;
        RECT 1938.510 161.940 2456.790 162.080 ;
        RECT 1938.510 161.880 1938.830 161.940 ;
        RECT 2456.470 161.880 2456.790 161.940 ;
      LAYER via ;
        RECT 1938.540 161.880 1938.800 162.140 ;
        RECT 2456.500 161.880 2456.760 162.140 ;
      LAYER met2 ;
        RECT 1935.670 960.570 1935.950 964.000 ;
        RECT 1935.670 960.430 1938.740 960.570 ;
        RECT 1935.670 960.000 1935.950 960.430 ;
        RECT 1938.600 162.170 1938.740 960.430 ;
        RECT 1938.540 161.850 1938.800 162.170 ;
        RECT 2456.500 161.850 2456.760 162.170 ;
        RECT 2456.560 6.530 2456.700 161.850 ;
        RECT 2456.560 6.390 2459.000 6.530 ;
        RECT 2458.860 2.400 2459.000 6.390 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1948.170 947.140 1948.490 947.200 ;
        RECT 1952.310 947.140 1952.630 947.200 ;
        RECT 1948.170 947.000 1952.630 947.140 ;
        RECT 1948.170 946.940 1948.490 947.000 ;
        RECT 1952.310 946.940 1952.630 947.000 ;
        RECT 1952.310 93.060 1952.630 93.120 ;
        RECT 2470.730 93.060 2471.050 93.120 ;
        RECT 1952.310 92.920 2471.050 93.060 ;
        RECT 1952.310 92.860 1952.630 92.920 ;
        RECT 2470.730 92.860 2471.050 92.920 ;
        RECT 2470.730 17.920 2471.050 17.980 ;
        RECT 2476.710 17.920 2477.030 17.980 ;
        RECT 2470.730 17.780 2477.030 17.920 ;
        RECT 2470.730 17.720 2471.050 17.780 ;
        RECT 2476.710 17.720 2477.030 17.780 ;
      LAYER via ;
        RECT 1948.200 946.940 1948.460 947.200 ;
        RECT 1952.340 946.940 1952.600 947.200 ;
        RECT 1952.340 92.860 1952.600 93.120 ;
        RECT 2470.760 92.860 2471.020 93.120 ;
        RECT 2470.760 17.720 2471.020 17.980 ;
        RECT 2476.740 17.720 2477.000 17.980 ;
      LAYER met2 ;
        RECT 1948.090 960.500 1948.370 964.000 ;
        RECT 1948.090 960.000 1948.400 960.500 ;
        RECT 1948.260 947.230 1948.400 960.000 ;
        RECT 1948.200 946.910 1948.460 947.230 ;
        RECT 1952.340 946.910 1952.600 947.230 ;
        RECT 1952.400 93.150 1952.540 946.910 ;
        RECT 1952.340 92.830 1952.600 93.150 ;
        RECT 2470.760 92.830 2471.020 93.150 ;
        RECT 2470.820 18.010 2470.960 92.830 ;
        RECT 2470.760 17.690 2471.020 18.010 ;
        RECT 2476.740 17.690 2477.000 18.010 ;
        RECT 2476.800 2.400 2476.940 17.690 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1960.590 951.220 1960.910 951.280 ;
        RECT 1965.650 951.220 1965.970 951.280 ;
        RECT 1960.590 951.080 1965.970 951.220 ;
        RECT 1960.590 951.020 1960.910 951.080 ;
        RECT 1965.650 951.020 1965.970 951.080 ;
        RECT 1965.650 769.320 1965.970 769.380 ;
        RECT 2490.970 769.320 2491.290 769.380 ;
        RECT 1965.650 769.180 2491.290 769.320 ;
        RECT 1965.650 769.120 1965.970 769.180 ;
        RECT 2490.970 769.120 2491.290 769.180 ;
      LAYER via ;
        RECT 1960.620 951.020 1960.880 951.280 ;
        RECT 1965.680 951.020 1965.940 951.280 ;
        RECT 1965.680 769.120 1965.940 769.380 ;
        RECT 2491.000 769.120 2491.260 769.380 ;
      LAYER met2 ;
        RECT 1960.510 960.500 1960.790 964.000 ;
        RECT 1960.510 960.000 1960.820 960.500 ;
        RECT 1960.680 951.310 1960.820 960.000 ;
        RECT 1960.620 950.990 1960.880 951.310 ;
        RECT 1965.680 950.990 1965.940 951.310 ;
        RECT 1965.740 769.410 1965.880 950.990 ;
        RECT 1965.680 769.090 1965.940 769.410 ;
        RECT 2491.000 769.090 2491.260 769.410 ;
        RECT 2491.060 17.410 2491.200 769.090 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 176.020 1973.330 176.080 ;
        RECT 2512.130 176.020 2512.450 176.080 ;
        RECT 1973.010 175.880 2512.450 176.020 ;
        RECT 1973.010 175.820 1973.330 175.880 ;
        RECT 2512.130 175.820 2512.450 175.880 ;
      LAYER via ;
        RECT 1973.040 175.820 1973.300 176.080 ;
        RECT 2512.160 175.820 2512.420 176.080 ;
      LAYER met2 ;
        RECT 1972.930 960.500 1973.210 964.000 ;
        RECT 1972.930 960.000 1973.240 960.500 ;
        RECT 1973.100 176.110 1973.240 960.000 ;
        RECT 1973.040 175.790 1973.300 176.110 ;
        RECT 2512.160 175.790 2512.420 176.110 ;
        RECT 2512.220 2.400 2512.360 175.790 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1986.810 762.520 1987.130 762.580 ;
        RECT 2525.470 762.520 2525.790 762.580 ;
        RECT 1986.810 762.380 2525.790 762.520 ;
        RECT 1986.810 762.320 1987.130 762.380 ;
        RECT 2525.470 762.320 2525.790 762.380 ;
        RECT 2525.470 2.960 2525.790 3.020 ;
        RECT 2530.070 2.960 2530.390 3.020 ;
        RECT 2525.470 2.820 2530.390 2.960 ;
        RECT 2525.470 2.760 2525.790 2.820 ;
        RECT 2530.070 2.760 2530.390 2.820 ;
      LAYER via ;
        RECT 1986.840 762.320 1987.100 762.580 ;
        RECT 2525.500 762.320 2525.760 762.580 ;
        RECT 2525.500 2.760 2525.760 3.020 ;
        RECT 2530.100 2.760 2530.360 3.020 ;
      LAYER met2 ;
        RECT 1985.350 960.570 1985.630 964.000 ;
        RECT 1985.350 960.430 1987.040 960.570 ;
        RECT 1985.350 960.000 1985.630 960.430 ;
        RECT 1986.900 762.610 1987.040 960.430 ;
        RECT 1986.840 762.290 1987.100 762.610 ;
        RECT 2525.500 762.290 2525.760 762.610 ;
        RECT 2525.560 3.050 2525.700 762.290 ;
        RECT 2525.500 2.730 2525.760 3.050 ;
        RECT 2530.100 2.730 2530.360 3.050 ;
        RECT 2530.160 2.400 2530.300 2.730 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2000.610 79.460 2000.930 79.520 ;
        RECT 2546.170 79.460 2546.490 79.520 ;
        RECT 2000.610 79.320 2546.490 79.460 ;
        RECT 2000.610 79.260 2000.930 79.320 ;
        RECT 2546.170 79.260 2546.490 79.320 ;
      LAYER via ;
        RECT 2000.640 79.260 2000.900 79.520 ;
        RECT 2546.200 79.260 2546.460 79.520 ;
      LAYER met2 ;
        RECT 1997.770 960.570 1998.050 964.000 ;
        RECT 1997.770 960.430 2000.840 960.570 ;
        RECT 1997.770 960.000 1998.050 960.430 ;
        RECT 2000.700 79.550 2000.840 960.430 ;
        RECT 2000.640 79.230 2000.900 79.550 ;
        RECT 2546.200 79.230 2546.460 79.550 ;
        RECT 2546.260 17.410 2546.400 79.230 ;
        RECT 2546.260 17.270 2548.240 17.410 ;
        RECT 2548.100 2.400 2548.240 17.270 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2010.270 945.440 2010.590 945.500 ;
        RECT 2014.410 945.440 2014.730 945.500 ;
        RECT 2010.270 945.300 2014.730 945.440 ;
        RECT 2010.270 945.240 2010.590 945.300 ;
        RECT 2014.410 945.240 2014.730 945.300 ;
        RECT 2014.410 210.360 2014.730 210.420 ;
        RECT 2560.430 210.360 2560.750 210.420 ;
        RECT 2014.410 210.220 2560.750 210.360 ;
        RECT 2014.410 210.160 2014.730 210.220 ;
        RECT 2560.430 210.160 2560.750 210.220 ;
      LAYER via ;
        RECT 2010.300 945.240 2010.560 945.500 ;
        RECT 2014.440 945.240 2014.700 945.500 ;
        RECT 2014.440 210.160 2014.700 210.420 ;
        RECT 2560.460 210.160 2560.720 210.420 ;
      LAYER met2 ;
        RECT 2010.190 960.500 2010.470 964.000 ;
        RECT 2010.190 960.000 2010.500 960.500 ;
        RECT 2010.360 945.530 2010.500 960.000 ;
        RECT 2010.300 945.210 2010.560 945.530 ;
        RECT 2014.440 945.210 2014.700 945.530 ;
        RECT 2014.500 210.450 2014.640 945.210 ;
        RECT 2014.440 210.130 2014.700 210.450 ;
        RECT 2560.460 210.130 2560.720 210.450 ;
        RECT 2560.520 17.410 2560.660 210.130 ;
        RECT 2560.520 17.270 2566.180 17.410 ;
        RECT 2566.040 2.400 2566.180 17.270 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2022.690 945.440 2023.010 945.500 ;
        RECT 2027.750 945.440 2028.070 945.500 ;
        RECT 2022.690 945.300 2028.070 945.440 ;
        RECT 2022.690 945.240 2023.010 945.300 ;
        RECT 2027.750 945.240 2028.070 945.300 ;
        RECT 2027.750 755.380 2028.070 755.440 ;
        RECT 2580.670 755.380 2580.990 755.440 ;
        RECT 2027.750 755.240 2580.990 755.380 ;
        RECT 2027.750 755.180 2028.070 755.240 ;
        RECT 2580.670 755.180 2580.990 755.240 ;
      LAYER via ;
        RECT 2022.720 945.240 2022.980 945.500 ;
        RECT 2027.780 945.240 2028.040 945.500 ;
        RECT 2027.780 755.180 2028.040 755.440 ;
        RECT 2580.700 755.180 2580.960 755.440 ;
      LAYER met2 ;
        RECT 2022.610 960.500 2022.890 964.000 ;
        RECT 2022.610 960.000 2022.920 960.500 ;
        RECT 2022.780 945.530 2022.920 960.000 ;
        RECT 2022.720 945.210 2022.980 945.530 ;
        RECT 2027.780 945.210 2028.040 945.530 ;
        RECT 2027.840 755.470 2027.980 945.210 ;
        RECT 2027.780 755.150 2028.040 755.470 ;
        RECT 2580.700 755.150 2580.960 755.470 ;
        RECT 2580.760 17.410 2580.900 755.150 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 20.640 800.330 20.700 ;
        RECT 817.490 20.640 817.810 20.700 ;
        RECT 800.010 20.500 817.810 20.640 ;
        RECT 800.010 20.440 800.330 20.500 ;
        RECT 817.490 20.440 817.810 20.500 ;
      LAYER via ;
        RECT 800.040 20.440 800.300 20.700 ;
        RECT 817.520 20.440 817.780 20.700 ;
      LAYER met2 ;
        RECT 797.630 960.570 797.910 964.000 ;
        RECT 797.630 960.430 800.240 960.570 ;
        RECT 797.630 960.000 797.910 960.430 ;
        RECT 800.100 20.730 800.240 960.430 ;
        RECT 800.040 20.410 800.300 20.730 ;
        RECT 817.520 20.410 817.780 20.730 ;
        RECT 817.580 2.400 817.720 20.410 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2035.110 237.900 2035.430 237.960 ;
        RECT 2601.830 237.900 2602.150 237.960 ;
        RECT 2035.110 237.760 2602.150 237.900 ;
        RECT 2035.110 237.700 2035.430 237.760 ;
        RECT 2601.830 237.700 2602.150 237.760 ;
      LAYER via ;
        RECT 2035.140 237.700 2035.400 237.960 ;
        RECT 2601.860 237.700 2602.120 237.960 ;
      LAYER met2 ;
        RECT 2034.570 960.570 2034.850 964.000 ;
        RECT 2034.570 960.430 2035.340 960.570 ;
        RECT 2034.570 960.000 2034.850 960.430 ;
        RECT 2035.200 237.990 2035.340 960.430 ;
        RECT 2035.140 237.670 2035.400 237.990 ;
        RECT 2601.860 237.670 2602.120 237.990 ;
        RECT 2601.920 7.890 2602.060 237.670 ;
        RECT 2601.460 7.750 2602.060 7.890 ;
        RECT 2601.460 2.400 2601.600 7.750 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2048.910 245.040 2049.230 245.100 ;
        RECT 2615.170 245.040 2615.490 245.100 ;
        RECT 2048.910 244.900 2615.490 245.040 ;
        RECT 2048.910 244.840 2049.230 244.900 ;
        RECT 2615.170 244.840 2615.490 244.900 ;
      LAYER via ;
        RECT 2048.940 244.840 2049.200 245.100 ;
        RECT 2615.200 244.840 2615.460 245.100 ;
      LAYER met2 ;
        RECT 2046.990 960.570 2047.270 964.000 ;
        RECT 2046.990 960.430 2049.140 960.570 ;
        RECT 2046.990 960.000 2047.270 960.430 ;
        RECT 2049.000 245.130 2049.140 960.430 ;
        RECT 2048.940 244.810 2049.200 245.130 ;
        RECT 2615.200 244.810 2615.460 245.130 ;
        RECT 2615.260 17.410 2615.400 244.810 ;
        RECT 2615.260 17.270 2619.540 17.410 ;
        RECT 2619.400 2.400 2619.540 17.270 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.710 107.000 2063.030 107.060 ;
        RECT 2635.870 107.000 2636.190 107.060 ;
        RECT 2062.710 106.860 2636.190 107.000 ;
        RECT 2062.710 106.800 2063.030 106.860 ;
        RECT 2635.870 106.800 2636.190 106.860 ;
      LAYER via ;
        RECT 2062.740 106.800 2063.000 107.060 ;
        RECT 2635.900 106.800 2636.160 107.060 ;
      LAYER met2 ;
        RECT 2059.410 960.570 2059.690 964.000 ;
        RECT 2059.410 960.430 2062.940 960.570 ;
        RECT 2059.410 960.000 2059.690 960.430 ;
        RECT 2062.800 107.090 2062.940 960.430 ;
        RECT 2062.740 106.770 2063.000 107.090 ;
        RECT 2635.900 106.770 2636.160 107.090 ;
        RECT 2635.960 17.410 2636.100 106.770 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2071.910 945.440 2072.230 945.500 ;
        RECT 2080.190 945.440 2080.510 945.500 ;
        RECT 2071.910 945.300 2080.510 945.440 ;
        RECT 2071.910 945.240 2072.230 945.300 ;
        RECT 2080.190 945.240 2080.510 945.300 ;
        RECT 2080.190 748.580 2080.510 748.640 ;
        RECT 2649.670 748.580 2649.990 748.640 ;
        RECT 2080.190 748.440 2649.990 748.580 ;
        RECT 2080.190 748.380 2080.510 748.440 ;
        RECT 2649.670 748.380 2649.990 748.440 ;
      LAYER via ;
        RECT 2071.940 945.240 2072.200 945.500 ;
        RECT 2080.220 945.240 2080.480 945.500 ;
        RECT 2080.220 748.380 2080.480 748.640 ;
        RECT 2649.700 748.380 2649.960 748.640 ;
      LAYER met2 ;
        RECT 2071.830 960.500 2072.110 964.000 ;
        RECT 2071.830 960.000 2072.140 960.500 ;
        RECT 2072.000 945.530 2072.140 960.000 ;
        RECT 2071.940 945.210 2072.200 945.530 ;
        RECT 2080.220 945.210 2080.480 945.530 ;
        RECT 2080.280 748.670 2080.420 945.210 ;
        RECT 2080.220 748.350 2080.480 748.670 ;
        RECT 2649.700 748.350 2649.960 748.670 ;
        RECT 2649.760 17.410 2649.900 748.350 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2084.330 951.220 2084.650 951.280 ;
        RECT 2089.850 951.220 2090.170 951.280 ;
        RECT 2084.330 951.080 2090.170 951.220 ;
        RECT 2084.330 951.020 2084.650 951.080 ;
        RECT 2089.850 951.020 2090.170 951.080 ;
        RECT 2089.850 741.780 2090.170 741.840 ;
        RECT 2670.370 741.780 2670.690 741.840 ;
        RECT 2089.850 741.640 2670.690 741.780 ;
        RECT 2089.850 741.580 2090.170 741.640 ;
        RECT 2670.370 741.580 2670.690 741.640 ;
      LAYER via ;
        RECT 2084.360 951.020 2084.620 951.280 ;
        RECT 2089.880 951.020 2090.140 951.280 ;
        RECT 2089.880 741.580 2090.140 741.840 ;
        RECT 2670.400 741.580 2670.660 741.840 ;
      LAYER met2 ;
        RECT 2084.250 960.500 2084.530 964.000 ;
        RECT 2084.250 960.000 2084.560 960.500 ;
        RECT 2084.420 951.310 2084.560 960.000 ;
        RECT 2084.360 950.990 2084.620 951.310 ;
        RECT 2089.880 950.990 2090.140 951.310 ;
        RECT 2089.940 741.870 2090.080 950.990 ;
        RECT 2089.880 741.550 2090.140 741.870 ;
        RECT 2670.400 741.550 2670.660 741.870 ;
        RECT 2670.460 17.410 2670.600 741.550 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2097.210 113.800 2097.530 113.860 ;
        RECT 2684.630 113.800 2684.950 113.860 ;
        RECT 2097.210 113.660 2684.950 113.800 ;
        RECT 2097.210 113.600 2097.530 113.660 ;
        RECT 2684.630 113.600 2684.950 113.660 ;
        RECT 2684.630 17.920 2684.950 17.980 ;
        RECT 2690.610 17.920 2690.930 17.980 ;
        RECT 2684.630 17.780 2690.930 17.920 ;
        RECT 2684.630 17.720 2684.950 17.780 ;
        RECT 2690.610 17.720 2690.930 17.780 ;
      LAYER via ;
        RECT 2097.240 113.600 2097.500 113.860 ;
        RECT 2684.660 113.600 2684.920 113.860 ;
        RECT 2684.660 17.720 2684.920 17.980 ;
        RECT 2690.640 17.720 2690.900 17.980 ;
      LAYER met2 ;
        RECT 2096.670 960.570 2096.950 964.000 ;
        RECT 2096.670 960.430 2097.440 960.570 ;
        RECT 2096.670 960.000 2096.950 960.430 ;
        RECT 2097.300 113.890 2097.440 960.430 ;
        RECT 2097.240 113.570 2097.500 113.890 ;
        RECT 2684.660 113.570 2684.920 113.890 ;
        RECT 2684.720 18.010 2684.860 113.570 ;
        RECT 2684.660 17.690 2684.920 18.010 ;
        RECT 2690.640 17.690 2690.900 18.010 ;
        RECT 2690.700 2.400 2690.840 17.690 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2111.010 120.600 2111.330 120.660 ;
        RECT 2704.870 120.600 2705.190 120.660 ;
        RECT 2111.010 120.460 2705.190 120.600 ;
        RECT 2111.010 120.400 2111.330 120.460 ;
        RECT 2704.870 120.400 2705.190 120.460 ;
      LAYER via ;
        RECT 2111.040 120.400 2111.300 120.660 ;
        RECT 2704.900 120.400 2705.160 120.660 ;
      LAYER met2 ;
        RECT 2109.090 960.570 2109.370 964.000 ;
        RECT 2109.090 960.430 2111.240 960.570 ;
        RECT 2109.090 960.000 2109.370 960.430 ;
        RECT 2111.100 120.690 2111.240 960.430 ;
        RECT 2111.040 120.370 2111.300 120.690 ;
        RECT 2704.900 120.370 2705.160 120.690 ;
        RECT 2704.960 17.410 2705.100 120.370 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 224.300 2125.130 224.360 ;
        RECT 2725.570 224.300 2725.890 224.360 ;
        RECT 2124.810 224.160 2725.890 224.300 ;
        RECT 2124.810 224.100 2125.130 224.160 ;
        RECT 2725.570 224.100 2725.890 224.160 ;
      LAYER via ;
        RECT 2124.840 224.100 2125.100 224.360 ;
        RECT 2725.600 224.100 2725.860 224.360 ;
      LAYER met2 ;
        RECT 2121.510 960.570 2121.790 964.000 ;
        RECT 2121.510 960.430 2125.040 960.570 ;
        RECT 2121.510 960.000 2121.790 960.430 ;
        RECT 2124.900 224.390 2125.040 960.430 ;
        RECT 2124.840 224.070 2125.100 224.390 ;
        RECT 2725.600 224.070 2725.860 224.390 ;
        RECT 2725.660 17.410 2725.800 224.070 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2134.010 945.440 2134.330 945.500 ;
        RECT 2138.150 945.440 2138.470 945.500 ;
        RECT 2134.010 945.300 2138.470 945.440 ;
        RECT 2134.010 945.240 2134.330 945.300 ;
        RECT 2138.150 945.240 2138.470 945.300 ;
        RECT 2138.150 734.640 2138.470 734.700 ;
        RECT 2739.370 734.640 2739.690 734.700 ;
        RECT 2138.150 734.500 2739.690 734.640 ;
        RECT 2138.150 734.440 2138.470 734.500 ;
        RECT 2739.370 734.440 2739.690 734.500 ;
      LAYER via ;
        RECT 2134.040 945.240 2134.300 945.500 ;
        RECT 2138.180 945.240 2138.440 945.500 ;
        RECT 2138.180 734.440 2138.440 734.700 ;
        RECT 2739.400 734.440 2739.660 734.700 ;
      LAYER met2 ;
        RECT 2133.930 960.500 2134.210 964.000 ;
        RECT 2133.930 960.000 2134.240 960.500 ;
        RECT 2134.100 945.530 2134.240 960.000 ;
        RECT 2134.040 945.210 2134.300 945.530 ;
        RECT 2138.180 945.210 2138.440 945.530 ;
        RECT 2138.240 734.730 2138.380 945.210 ;
        RECT 2138.180 734.410 2138.440 734.730 ;
        RECT 2739.400 734.410 2739.660 734.730 ;
        RECT 2739.460 17.410 2739.600 734.410 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.970 949.860 2146.290 949.920 ;
        RECT 2151.950 949.860 2152.270 949.920 ;
        RECT 2145.970 949.720 2152.270 949.860 ;
        RECT 2145.970 949.660 2146.290 949.720 ;
        RECT 2151.950 949.660 2152.270 949.720 ;
        RECT 2151.950 727.840 2152.270 727.900 ;
        RECT 2760.070 727.840 2760.390 727.900 ;
        RECT 2151.950 727.700 2760.390 727.840 ;
        RECT 2151.950 727.640 2152.270 727.700 ;
        RECT 2760.070 727.640 2760.390 727.700 ;
      LAYER via ;
        RECT 2146.000 949.660 2146.260 949.920 ;
        RECT 2151.980 949.660 2152.240 949.920 ;
        RECT 2151.980 727.640 2152.240 727.900 ;
        RECT 2760.100 727.640 2760.360 727.900 ;
      LAYER met2 ;
        RECT 2145.890 960.500 2146.170 964.000 ;
        RECT 2145.890 960.000 2146.200 960.500 ;
        RECT 2146.060 949.950 2146.200 960.000 ;
        RECT 2146.000 949.630 2146.260 949.950 ;
        RECT 2151.980 949.630 2152.240 949.950 ;
        RECT 2152.040 727.930 2152.180 949.630 ;
        RECT 2151.980 727.610 2152.240 727.930 ;
        RECT 2760.100 727.610 2760.360 727.930 ;
        RECT 2760.160 17.410 2760.300 727.610 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.810 17.580 814.130 17.640 ;
        RECT 835.430 17.580 835.750 17.640 ;
        RECT 813.810 17.440 835.750 17.580 ;
        RECT 813.810 17.380 814.130 17.440 ;
        RECT 835.430 17.380 835.750 17.440 ;
      LAYER via ;
        RECT 813.840 17.380 814.100 17.640 ;
        RECT 835.460 17.380 835.720 17.640 ;
      LAYER met2 ;
        RECT 810.050 960.570 810.330 964.000 ;
        RECT 810.050 960.430 814.040 960.570 ;
        RECT 810.050 960.000 810.330 960.430 ;
        RECT 813.900 17.670 814.040 960.430 ;
        RECT 813.840 17.350 814.100 17.670 ;
        RECT 835.460 17.350 835.720 17.670 ;
        RECT 835.520 2.400 835.660 17.350 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2159.310 189.620 2159.630 189.680 ;
        RECT 2774.330 189.620 2774.650 189.680 ;
        RECT 2159.310 189.480 2774.650 189.620 ;
        RECT 2159.310 189.420 2159.630 189.480 ;
        RECT 2774.330 189.420 2774.650 189.480 ;
      LAYER via ;
        RECT 2159.340 189.420 2159.600 189.680 ;
        RECT 2774.360 189.420 2774.620 189.680 ;
      LAYER met2 ;
        RECT 2158.310 960.570 2158.590 964.000 ;
        RECT 2158.310 960.430 2159.540 960.570 ;
        RECT 2158.310 960.000 2158.590 960.430 ;
        RECT 2159.400 189.710 2159.540 960.430 ;
        RECT 2159.340 189.390 2159.600 189.710 ;
        RECT 2774.360 189.390 2774.620 189.710 ;
        RECT 2774.420 17.410 2774.560 189.390 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2173.110 251.840 2173.430 251.900 ;
        RECT 2794.570 251.840 2794.890 251.900 ;
        RECT 2173.110 251.700 2794.890 251.840 ;
        RECT 2173.110 251.640 2173.430 251.700 ;
        RECT 2794.570 251.640 2794.890 251.700 ;
      LAYER via ;
        RECT 2173.140 251.640 2173.400 251.900 ;
        RECT 2794.600 251.640 2794.860 251.900 ;
      LAYER met2 ;
        RECT 2170.730 960.570 2171.010 964.000 ;
        RECT 2170.730 960.430 2173.340 960.570 ;
        RECT 2170.730 960.000 2171.010 960.430 ;
        RECT 2173.200 251.930 2173.340 960.430 ;
        RECT 2173.140 251.610 2173.400 251.930 ;
        RECT 2794.600 251.610 2794.860 251.930 ;
        RECT 2794.660 17.410 2794.800 251.610 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2183.230 945.440 2183.550 945.500 ;
        RECT 2186.910 945.440 2187.230 945.500 ;
        RECT 2183.230 945.300 2187.230 945.440 ;
        RECT 2183.230 945.240 2183.550 945.300 ;
        RECT 2186.910 945.240 2187.230 945.300 ;
        RECT 2186.910 721.040 2187.230 721.100 ;
        RECT 2815.270 721.040 2815.590 721.100 ;
        RECT 2186.910 720.900 2815.590 721.040 ;
        RECT 2186.910 720.840 2187.230 720.900 ;
        RECT 2815.270 720.840 2815.590 720.900 ;
      LAYER via ;
        RECT 2183.260 945.240 2183.520 945.500 ;
        RECT 2186.940 945.240 2187.200 945.500 ;
        RECT 2186.940 720.840 2187.200 721.100 ;
        RECT 2815.300 720.840 2815.560 721.100 ;
      LAYER met2 ;
        RECT 2183.150 960.500 2183.430 964.000 ;
        RECT 2183.150 960.000 2183.460 960.500 ;
        RECT 2183.320 945.530 2183.460 960.000 ;
        RECT 2183.260 945.210 2183.520 945.530 ;
        RECT 2186.940 945.210 2187.200 945.530 ;
        RECT 2187.000 721.130 2187.140 945.210 ;
        RECT 2186.940 720.810 2187.200 721.130 ;
        RECT 2815.300 720.810 2815.560 721.130 ;
        RECT 2815.360 17.410 2815.500 720.810 ;
        RECT 2815.360 17.270 2815.960 17.410 ;
        RECT 2815.820 2.400 2815.960 17.270 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2195.650 946.460 2195.970 946.520 ;
        RECT 2200.250 946.460 2200.570 946.520 ;
        RECT 2195.650 946.320 2200.570 946.460 ;
        RECT 2195.650 946.260 2195.970 946.320 ;
        RECT 2200.250 946.260 2200.570 946.320 ;
        RECT 2200.250 714.240 2200.570 714.300 ;
        RECT 2829.070 714.240 2829.390 714.300 ;
        RECT 2200.250 714.100 2829.390 714.240 ;
        RECT 2200.250 714.040 2200.570 714.100 ;
        RECT 2829.070 714.040 2829.390 714.100 ;
      LAYER via ;
        RECT 2195.680 946.260 2195.940 946.520 ;
        RECT 2200.280 946.260 2200.540 946.520 ;
        RECT 2200.280 714.040 2200.540 714.300 ;
        RECT 2829.100 714.040 2829.360 714.300 ;
      LAYER met2 ;
        RECT 2195.570 960.500 2195.850 964.000 ;
        RECT 2195.570 960.000 2195.880 960.500 ;
        RECT 2195.740 946.550 2195.880 960.000 ;
        RECT 2195.680 946.230 2195.940 946.550 ;
        RECT 2200.280 946.230 2200.540 946.550 ;
        RECT 2200.340 714.330 2200.480 946.230 ;
        RECT 2200.280 714.010 2200.540 714.330 ;
        RECT 2829.100 714.010 2829.360 714.330 ;
        RECT 2829.160 17.410 2829.300 714.010 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2208.070 950.880 2208.390 950.940 ;
        RECT 2214.050 950.880 2214.370 950.940 ;
        RECT 2208.070 950.740 2214.370 950.880 ;
        RECT 2208.070 950.680 2208.390 950.740 ;
        RECT 2214.050 950.680 2214.370 950.740 ;
        RECT 2214.050 707.100 2214.370 707.160 ;
        RECT 2849.770 707.100 2850.090 707.160 ;
        RECT 2214.050 706.960 2850.090 707.100 ;
        RECT 2214.050 706.900 2214.370 706.960 ;
        RECT 2849.770 706.900 2850.090 706.960 ;
      LAYER via ;
        RECT 2208.100 950.680 2208.360 950.940 ;
        RECT 2214.080 950.680 2214.340 950.940 ;
        RECT 2214.080 706.900 2214.340 707.160 ;
        RECT 2849.800 706.900 2850.060 707.160 ;
      LAYER met2 ;
        RECT 2207.990 960.500 2208.270 964.000 ;
        RECT 2207.990 960.000 2208.300 960.500 ;
        RECT 2208.160 950.970 2208.300 960.000 ;
        RECT 2208.100 950.650 2208.360 950.970 ;
        RECT 2214.080 950.650 2214.340 950.970 ;
        RECT 2214.140 707.190 2214.280 950.650 ;
        RECT 2214.080 706.870 2214.340 707.190 ;
        RECT 2849.800 706.870 2850.060 707.190 ;
        RECT 2849.860 17.410 2850.000 706.870 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2221.410 258.640 2221.730 258.700 ;
        RECT 2863.570 258.640 2863.890 258.700 ;
        RECT 2221.410 258.500 2863.890 258.640 ;
        RECT 2221.410 258.440 2221.730 258.500 ;
        RECT 2863.570 258.440 2863.890 258.500 ;
      LAYER via ;
        RECT 2221.440 258.440 2221.700 258.700 ;
        RECT 2863.600 258.440 2863.860 258.700 ;
      LAYER met2 ;
        RECT 2220.410 960.570 2220.690 964.000 ;
        RECT 2220.410 960.430 2221.640 960.570 ;
        RECT 2220.410 960.000 2220.690 960.430 ;
        RECT 2221.500 258.730 2221.640 960.430 ;
        RECT 2221.440 258.410 2221.700 258.730 ;
        RECT 2863.600 258.410 2863.860 258.730 ;
        RECT 2863.660 17.410 2863.800 258.410 ;
        RECT 2863.660 17.270 2869.320 17.410 ;
        RECT 2869.180 2.400 2869.320 17.270 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2235.210 168.880 2235.530 168.940 ;
        RECT 2884.270 168.880 2884.590 168.940 ;
        RECT 2235.210 168.740 2884.590 168.880 ;
        RECT 2235.210 168.680 2235.530 168.740 ;
        RECT 2884.270 168.680 2884.590 168.740 ;
        RECT 2884.270 2.960 2884.590 3.020 ;
        RECT 2887.030 2.960 2887.350 3.020 ;
        RECT 2884.270 2.820 2887.350 2.960 ;
        RECT 2884.270 2.760 2884.590 2.820 ;
        RECT 2887.030 2.760 2887.350 2.820 ;
      LAYER via ;
        RECT 2235.240 168.680 2235.500 168.940 ;
        RECT 2884.300 168.680 2884.560 168.940 ;
        RECT 2884.300 2.760 2884.560 3.020 ;
        RECT 2887.060 2.760 2887.320 3.020 ;
      LAYER met2 ;
        RECT 2232.830 960.570 2233.110 964.000 ;
        RECT 2232.830 960.430 2235.440 960.570 ;
        RECT 2232.830 960.000 2233.110 960.430 ;
        RECT 2235.300 168.970 2235.440 960.430 ;
        RECT 2235.240 168.650 2235.500 168.970 ;
        RECT 2884.300 168.650 2884.560 168.970 ;
        RECT 2884.360 3.050 2884.500 168.650 ;
        RECT 2884.300 2.730 2884.560 3.050 ;
        RECT 2887.060 2.730 2887.320 3.050 ;
        RECT 2887.120 2.400 2887.260 2.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2249.010 182.820 2249.330 182.880 ;
        RECT 2894.850 182.820 2895.170 182.880 ;
        RECT 2249.010 182.680 2895.170 182.820 ;
        RECT 2249.010 182.620 2249.330 182.680 ;
        RECT 2894.850 182.620 2895.170 182.680 ;
        RECT 2894.850 17.580 2895.170 17.640 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2894.850 17.440 2905.290 17.580 ;
        RECT 2894.850 17.380 2895.170 17.440 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
      LAYER via ;
        RECT 2249.040 182.620 2249.300 182.880 ;
        RECT 2894.880 182.620 2895.140 182.880 ;
        RECT 2894.880 17.380 2895.140 17.640 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
      LAYER met2 ;
        RECT 2245.250 960.570 2245.530 964.000 ;
        RECT 2245.250 960.430 2249.240 960.570 ;
        RECT 2245.250 960.000 2245.530 960.430 ;
        RECT 2249.100 182.910 2249.240 960.430 ;
        RECT 2249.040 182.590 2249.300 182.910 ;
        RECT 2894.880 182.590 2895.140 182.910 ;
        RECT 2894.940 17.670 2895.080 182.590 ;
        RECT 2894.880 17.350 2895.140 17.670 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2905.060 2.400 2905.200 17.350 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 822.550 950.540 822.870 950.600 ;
        RECT 827.150 950.540 827.470 950.600 ;
        RECT 822.550 950.400 827.470 950.540 ;
        RECT 822.550 950.340 822.870 950.400 ;
        RECT 827.150 950.340 827.470 950.400 ;
        RECT 827.150 17.920 827.470 17.980 ;
        RECT 852.910 17.920 853.230 17.980 ;
        RECT 827.150 17.780 853.230 17.920 ;
        RECT 827.150 17.720 827.470 17.780 ;
        RECT 852.910 17.720 853.230 17.780 ;
      LAYER via ;
        RECT 822.580 950.340 822.840 950.600 ;
        RECT 827.180 950.340 827.440 950.600 ;
        RECT 827.180 17.720 827.440 17.980 ;
        RECT 852.940 17.720 853.200 17.980 ;
      LAYER met2 ;
        RECT 822.470 960.500 822.750 964.000 ;
        RECT 822.470 960.000 822.780 960.500 ;
        RECT 822.640 950.630 822.780 960.000 ;
        RECT 822.580 950.310 822.840 950.630 ;
        RECT 827.180 950.310 827.440 950.630 ;
        RECT 827.240 18.010 827.380 950.310 ;
        RECT 827.180 17.690 827.440 18.010 ;
        RECT 852.940 17.690 853.200 18.010 ;
        RECT 853.000 2.400 853.140 17.690 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 834.970 945.440 835.290 945.500 ;
        RECT 840.950 945.440 841.270 945.500 ;
        RECT 834.970 945.300 841.270 945.440 ;
        RECT 834.970 945.240 835.290 945.300 ;
        RECT 840.950 945.240 841.270 945.300 ;
        RECT 840.950 18.260 841.270 18.320 ;
        RECT 870.850 18.260 871.170 18.320 ;
        RECT 840.950 18.120 871.170 18.260 ;
        RECT 840.950 18.060 841.270 18.120 ;
        RECT 870.850 18.060 871.170 18.120 ;
      LAYER via ;
        RECT 835.000 945.240 835.260 945.500 ;
        RECT 840.980 945.240 841.240 945.500 ;
        RECT 840.980 18.060 841.240 18.320 ;
        RECT 870.880 18.060 871.140 18.320 ;
      LAYER met2 ;
        RECT 834.890 960.500 835.170 964.000 ;
        RECT 834.890 960.000 835.200 960.500 ;
        RECT 835.060 945.530 835.200 960.000 ;
        RECT 835.000 945.210 835.260 945.530 ;
        RECT 840.980 945.210 841.240 945.530 ;
        RECT 841.040 18.350 841.180 945.210 ;
        RECT 840.980 18.030 841.240 18.350 ;
        RECT 870.880 18.030 871.140 18.350 ;
        RECT 870.940 2.400 871.080 18.030 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 848.310 19.280 848.630 19.340 ;
        RECT 888.790 19.280 889.110 19.340 ;
        RECT 848.310 19.140 889.110 19.280 ;
        RECT 848.310 19.080 848.630 19.140 ;
        RECT 888.790 19.080 889.110 19.140 ;
      LAYER via ;
        RECT 848.340 19.080 848.600 19.340 ;
        RECT 888.820 19.080 889.080 19.340 ;
      LAYER met2 ;
        RECT 847.310 960.570 847.590 964.000 ;
        RECT 847.310 960.430 848.540 960.570 ;
        RECT 847.310 960.000 847.590 960.430 ;
        RECT 848.400 19.370 848.540 960.430 ;
        RECT 848.340 19.050 848.600 19.370 ;
        RECT 888.820 19.050 889.080 19.370 ;
        RECT 888.880 2.400 889.020 19.050 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 861.650 17.920 861.970 17.980 ;
        RECT 906.730 17.920 907.050 17.980 ;
        RECT 861.650 17.780 907.050 17.920 ;
        RECT 861.650 17.720 861.970 17.780 ;
        RECT 906.730 17.720 907.050 17.780 ;
      LAYER via ;
        RECT 861.680 17.720 861.940 17.980 ;
        RECT 906.760 17.720 907.020 17.980 ;
      LAYER met2 ;
        RECT 859.730 960.570 860.010 964.000 ;
        RECT 859.730 960.430 861.880 960.570 ;
        RECT 859.730 960.000 860.010 960.430 ;
        RECT 861.740 18.010 861.880 960.430 ;
        RECT 861.680 17.690 861.940 18.010 ;
        RECT 906.760 17.690 907.020 18.010 ;
        RECT 906.820 2.400 906.960 17.690 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 872.230 945.440 872.550 945.500 ;
        RECT 875.910 945.440 876.230 945.500 ;
        RECT 872.230 945.300 876.230 945.440 ;
        RECT 872.230 945.240 872.550 945.300 ;
        RECT 875.910 945.240 876.230 945.300 ;
        RECT 875.910 18.260 876.230 18.320 ;
        RECT 924.210 18.260 924.530 18.320 ;
        RECT 875.910 18.120 924.530 18.260 ;
        RECT 875.910 18.060 876.230 18.120 ;
        RECT 924.210 18.060 924.530 18.120 ;
      LAYER via ;
        RECT 872.260 945.240 872.520 945.500 ;
        RECT 875.940 945.240 876.200 945.500 ;
        RECT 875.940 18.060 876.200 18.320 ;
        RECT 924.240 18.060 924.500 18.320 ;
      LAYER met2 ;
        RECT 872.150 960.500 872.430 964.000 ;
        RECT 872.150 960.000 872.460 960.500 ;
        RECT 872.320 945.530 872.460 960.000 ;
        RECT 872.260 945.210 872.520 945.530 ;
        RECT 875.940 945.210 876.200 945.530 ;
        RECT 876.000 18.350 876.140 945.210 ;
        RECT 875.940 18.030 876.200 18.350 ;
        RECT 924.240 18.030 924.500 18.350 ;
        RECT 924.300 2.400 924.440 18.030 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 884.650 945.440 884.970 945.500 ;
        RECT 889.250 945.440 889.570 945.500 ;
        RECT 884.650 945.300 889.570 945.440 ;
        RECT 884.650 945.240 884.970 945.300 ;
        RECT 889.250 945.240 889.570 945.300 ;
        RECT 889.250 19.620 889.570 19.680 ;
        RECT 942.150 19.620 942.470 19.680 ;
        RECT 889.250 19.480 942.470 19.620 ;
        RECT 889.250 19.420 889.570 19.480 ;
        RECT 942.150 19.420 942.470 19.480 ;
      LAYER via ;
        RECT 884.680 945.240 884.940 945.500 ;
        RECT 889.280 945.240 889.540 945.500 ;
        RECT 889.280 19.420 889.540 19.680 ;
        RECT 942.180 19.420 942.440 19.680 ;
      LAYER met2 ;
        RECT 884.570 960.500 884.850 964.000 ;
        RECT 884.570 960.000 884.880 960.500 ;
        RECT 884.740 945.530 884.880 960.000 ;
        RECT 884.680 945.210 884.940 945.530 ;
        RECT 889.280 945.210 889.540 945.530 ;
        RECT 889.340 19.710 889.480 945.210 ;
        RECT 889.280 19.390 889.540 19.710 ;
        RECT 942.180 19.390 942.440 19.710 ;
        RECT 942.240 2.400 942.380 19.390 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 896.610 17.240 896.930 17.300 ;
        RECT 960.090 17.240 960.410 17.300 ;
        RECT 896.610 17.100 960.410 17.240 ;
        RECT 896.610 17.040 896.930 17.100 ;
        RECT 960.090 17.040 960.410 17.100 ;
      LAYER via ;
        RECT 896.640 17.040 896.900 17.300 ;
        RECT 960.120 17.040 960.380 17.300 ;
      LAYER met2 ;
        RECT 896.530 960.500 896.810 964.000 ;
        RECT 896.530 960.000 896.840 960.500 ;
        RECT 896.700 17.330 896.840 960.000 ;
        RECT 896.640 17.010 896.900 17.330 ;
        RECT 960.120 17.010 960.380 17.330 ;
        RECT 960.180 2.400 960.320 17.010 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.410 19.280 910.730 19.340 ;
        RECT 978.030 19.280 978.350 19.340 ;
        RECT 910.410 19.140 978.350 19.280 ;
        RECT 910.410 19.080 910.730 19.140 ;
        RECT 978.030 19.080 978.350 19.140 ;
      LAYER via ;
        RECT 910.440 19.080 910.700 19.340 ;
        RECT 978.060 19.080 978.320 19.340 ;
      LAYER met2 ;
        RECT 908.950 960.570 909.230 964.000 ;
        RECT 908.950 960.430 910.640 960.570 ;
        RECT 908.950 960.000 909.230 960.430 ;
        RECT 910.500 19.370 910.640 960.430 ;
        RECT 910.440 19.050 910.700 19.370 ;
        RECT 978.060 19.050 978.320 19.370 ;
        RECT 978.120 2.400 978.260 19.050 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 15.200 657.270 15.260 ;
        RECT 683.170 15.200 683.490 15.260 ;
        RECT 656.950 15.060 683.490 15.200 ;
        RECT 656.950 15.000 657.270 15.060 ;
        RECT 683.170 15.000 683.490 15.060 ;
      LAYER via ;
        RECT 656.980 15.000 657.240 15.260 ;
        RECT 683.200 15.000 683.460 15.260 ;
      LAYER met2 ;
        RECT 686.310 960.570 686.590 964.000 ;
        RECT 683.260 960.430 686.590 960.570 ;
        RECT 683.260 15.290 683.400 960.430 ;
        RECT 686.310 960.000 686.590 960.430 ;
        RECT 656.980 14.970 657.240 15.290 ;
        RECT 683.200 14.970 683.460 15.290 ;
        RECT 657.040 2.400 657.180 14.970 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 58.720 924.530 58.780 ;
        RECT 993.670 58.720 993.990 58.780 ;
        RECT 924.210 58.580 993.990 58.720 ;
        RECT 924.210 58.520 924.530 58.580 ;
        RECT 993.670 58.520 993.990 58.580 ;
      LAYER via ;
        RECT 924.240 58.520 924.500 58.780 ;
        RECT 993.700 58.520 993.960 58.780 ;
      LAYER met2 ;
        RECT 921.370 960.570 921.650 964.000 ;
        RECT 921.370 960.430 924.440 960.570 ;
        RECT 921.370 960.000 921.650 960.430 ;
        RECT 924.300 58.810 924.440 960.430 ;
        RECT 924.240 58.490 924.500 58.810 ;
        RECT 993.700 58.490 993.960 58.810 ;
        RECT 993.760 16.730 993.900 58.490 ;
        RECT 993.760 16.590 996.200 16.730 ;
        RECT 996.060 2.400 996.200 16.590 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 933.870 945.440 934.190 945.500 ;
        RECT 937.550 945.440 937.870 945.500 ;
        RECT 933.870 945.300 937.870 945.440 ;
        RECT 933.870 945.240 934.190 945.300 ;
        RECT 937.550 945.240 937.870 945.300 ;
        RECT 937.550 65.520 937.870 65.580 ;
        RECT 1007.470 65.520 1007.790 65.580 ;
        RECT 937.550 65.380 1007.790 65.520 ;
        RECT 937.550 65.320 937.870 65.380 ;
        RECT 1007.470 65.320 1007.790 65.380 ;
        RECT 1007.470 17.580 1007.790 17.640 ;
        RECT 1013.450 17.580 1013.770 17.640 ;
        RECT 1007.470 17.440 1013.770 17.580 ;
        RECT 1007.470 17.380 1007.790 17.440 ;
        RECT 1013.450 17.380 1013.770 17.440 ;
      LAYER via ;
        RECT 933.900 945.240 934.160 945.500 ;
        RECT 937.580 945.240 937.840 945.500 ;
        RECT 937.580 65.320 937.840 65.580 ;
        RECT 1007.500 65.320 1007.760 65.580 ;
        RECT 1007.500 17.380 1007.760 17.640 ;
        RECT 1013.480 17.380 1013.740 17.640 ;
      LAYER met2 ;
        RECT 933.790 960.500 934.070 964.000 ;
        RECT 933.790 960.000 934.100 960.500 ;
        RECT 933.960 945.530 934.100 960.000 ;
        RECT 933.900 945.210 934.160 945.530 ;
        RECT 937.580 945.210 937.840 945.530 ;
        RECT 937.640 65.610 937.780 945.210 ;
        RECT 937.580 65.290 937.840 65.610 ;
        RECT 1007.500 65.290 1007.760 65.610 ;
        RECT 1007.560 17.670 1007.700 65.290 ;
        RECT 1007.500 17.350 1007.760 17.670 ;
        RECT 1013.480 17.350 1013.740 17.670 ;
        RECT 1013.540 2.400 1013.680 17.350 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 946.290 945.440 946.610 945.500 ;
        RECT 951.350 945.440 951.670 945.500 ;
        RECT 946.290 945.300 951.670 945.440 ;
        RECT 946.290 945.240 946.610 945.300 ;
        RECT 951.350 945.240 951.670 945.300 ;
        RECT 951.350 72.320 951.670 72.380 ;
        RECT 1028.170 72.320 1028.490 72.380 ;
        RECT 951.350 72.180 1028.490 72.320 ;
        RECT 951.350 72.120 951.670 72.180 ;
        RECT 1028.170 72.120 1028.490 72.180 ;
      LAYER via ;
        RECT 946.320 945.240 946.580 945.500 ;
        RECT 951.380 945.240 951.640 945.500 ;
        RECT 951.380 72.120 951.640 72.380 ;
        RECT 1028.200 72.120 1028.460 72.380 ;
      LAYER met2 ;
        RECT 946.210 960.500 946.490 964.000 ;
        RECT 946.210 960.000 946.520 960.500 ;
        RECT 946.380 945.530 946.520 960.000 ;
        RECT 946.320 945.210 946.580 945.530 ;
        RECT 951.380 945.210 951.640 945.530 ;
        RECT 951.440 72.410 951.580 945.210 ;
        RECT 951.380 72.090 951.640 72.410 ;
        RECT 1028.200 72.090 1028.460 72.410 ;
        RECT 1028.260 16.730 1028.400 72.090 ;
        RECT 1028.260 16.590 1031.620 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 958.250 79.460 958.570 79.520 ;
        RECT 1049.330 79.460 1049.650 79.520 ;
        RECT 958.250 79.320 1049.650 79.460 ;
        RECT 958.250 79.260 958.570 79.320 ;
        RECT 1049.330 79.260 1049.650 79.320 ;
      LAYER via ;
        RECT 958.280 79.260 958.540 79.520 ;
        RECT 1049.360 79.260 1049.620 79.520 ;
      LAYER met2 ;
        RECT 958.630 960.570 958.910 964.000 ;
        RECT 958.340 960.430 958.910 960.570 ;
        RECT 958.340 79.550 958.480 960.430 ;
        RECT 958.630 960.000 958.910 960.430 ;
        RECT 958.280 79.230 958.540 79.550 ;
        RECT 1049.360 79.230 1049.620 79.550 ;
        RECT 1049.420 2.400 1049.560 79.230 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 972.050 86.260 972.370 86.320 ;
        RECT 1062.670 86.260 1062.990 86.320 ;
        RECT 972.050 86.120 1062.990 86.260 ;
        RECT 972.050 86.060 972.370 86.120 ;
        RECT 1062.670 86.060 1062.990 86.120 ;
      LAYER via ;
        RECT 972.080 86.060 972.340 86.320 ;
        RECT 1062.700 86.060 1062.960 86.320 ;
      LAYER met2 ;
        RECT 971.050 960.570 971.330 964.000 ;
        RECT 971.050 960.430 972.280 960.570 ;
        RECT 971.050 960.000 971.330 960.430 ;
        RECT 972.140 86.350 972.280 960.430 ;
        RECT 972.080 86.030 972.340 86.350 ;
        RECT 1062.700 86.030 1062.960 86.350 ;
        RECT 1062.760 18.090 1062.900 86.030 ;
        RECT 1062.760 17.950 1067.500 18.090 ;
        RECT 1067.360 2.400 1067.500 17.950 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 986.310 93.400 986.630 93.460 ;
        RECT 1083.370 93.400 1083.690 93.460 ;
        RECT 986.310 93.260 1083.690 93.400 ;
        RECT 986.310 93.200 986.630 93.260 ;
        RECT 1083.370 93.200 1083.690 93.260 ;
      LAYER via ;
        RECT 986.340 93.200 986.600 93.460 ;
        RECT 1083.400 93.200 1083.660 93.460 ;
      LAYER met2 ;
        RECT 983.470 960.570 983.750 964.000 ;
        RECT 983.470 960.430 986.540 960.570 ;
        RECT 983.470 960.000 983.750 960.430 ;
        RECT 986.400 93.490 986.540 960.430 ;
        RECT 986.340 93.170 986.600 93.490 ;
        RECT 1083.400 93.170 1083.660 93.490 ;
        RECT 1083.460 17.410 1083.600 93.170 ;
        RECT 1083.460 17.270 1085.440 17.410 ;
        RECT 1085.300 2.400 1085.440 17.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 995.970 945.440 996.290 945.500 ;
        RECT 1003.790 945.440 1004.110 945.500 ;
        RECT 995.970 945.300 1004.110 945.440 ;
        RECT 995.970 945.240 996.290 945.300 ;
        RECT 1003.790 945.240 1004.110 945.300 ;
        RECT 1003.790 100.200 1004.110 100.260 ;
        RECT 1097.170 100.200 1097.490 100.260 ;
        RECT 1003.790 100.060 1097.490 100.200 ;
        RECT 1003.790 100.000 1004.110 100.060 ;
        RECT 1097.170 100.000 1097.490 100.060 ;
      LAYER via ;
        RECT 996.000 945.240 996.260 945.500 ;
        RECT 1003.820 945.240 1004.080 945.500 ;
        RECT 1003.820 100.000 1004.080 100.260 ;
        RECT 1097.200 100.000 1097.460 100.260 ;
      LAYER met2 ;
        RECT 995.890 960.500 996.170 964.000 ;
        RECT 995.890 960.000 996.200 960.500 ;
        RECT 996.060 945.530 996.200 960.000 ;
        RECT 996.000 945.210 996.260 945.530 ;
        RECT 1003.820 945.210 1004.080 945.530 ;
        RECT 1003.880 100.290 1004.020 945.210 ;
        RECT 1003.820 99.970 1004.080 100.290 ;
        RECT 1097.200 99.970 1097.460 100.290 ;
        RECT 1097.260 16.730 1097.400 99.970 ;
        RECT 1097.260 16.590 1102.920 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1007.930 951.220 1008.250 951.280 ;
        RECT 1024.490 951.220 1024.810 951.280 ;
        RECT 1007.930 951.080 1024.810 951.220 ;
        RECT 1007.930 951.020 1008.250 951.080 ;
        RECT 1024.490 951.020 1024.810 951.080 ;
        RECT 1024.490 107.340 1024.810 107.400 ;
        RECT 1117.870 107.340 1118.190 107.400 ;
        RECT 1024.490 107.200 1118.190 107.340 ;
        RECT 1024.490 107.140 1024.810 107.200 ;
        RECT 1117.870 107.140 1118.190 107.200 ;
      LAYER via ;
        RECT 1007.960 951.020 1008.220 951.280 ;
        RECT 1024.520 951.020 1024.780 951.280 ;
        RECT 1024.520 107.140 1024.780 107.400 ;
        RECT 1117.900 107.140 1118.160 107.400 ;
      LAYER met2 ;
        RECT 1007.850 960.500 1008.130 964.000 ;
        RECT 1007.850 960.000 1008.160 960.500 ;
        RECT 1008.020 951.310 1008.160 960.000 ;
        RECT 1007.960 950.990 1008.220 951.310 ;
        RECT 1024.520 950.990 1024.780 951.310 ;
        RECT 1024.580 107.430 1024.720 950.990 ;
        RECT 1024.520 107.110 1024.780 107.430 ;
        RECT 1117.900 107.110 1118.160 107.430 ;
        RECT 1117.960 16.730 1118.100 107.110 ;
        RECT 1117.960 16.590 1120.860 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1020.350 113.800 1020.670 113.860 ;
        RECT 1139.030 113.800 1139.350 113.860 ;
        RECT 1020.350 113.660 1139.350 113.800 ;
        RECT 1020.350 113.600 1020.670 113.660 ;
        RECT 1139.030 113.600 1139.350 113.660 ;
      LAYER via ;
        RECT 1020.380 113.600 1020.640 113.860 ;
        RECT 1139.060 113.600 1139.320 113.860 ;
      LAYER met2 ;
        RECT 1020.270 960.500 1020.550 964.000 ;
        RECT 1020.270 960.000 1020.580 960.500 ;
        RECT 1020.440 113.890 1020.580 960.000 ;
        RECT 1020.380 113.570 1020.640 113.890 ;
        RECT 1139.060 113.570 1139.320 113.890 ;
        RECT 1139.120 7.210 1139.260 113.570 ;
        RECT 1138.660 7.070 1139.260 7.210 ;
        RECT 1138.660 2.400 1138.800 7.070 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.150 120.600 1034.470 120.660 ;
        RECT 1152.370 120.600 1152.690 120.660 ;
        RECT 1034.150 120.460 1152.690 120.600 ;
        RECT 1034.150 120.400 1034.470 120.460 ;
        RECT 1152.370 120.400 1152.690 120.460 ;
      LAYER via ;
        RECT 1034.180 120.400 1034.440 120.660 ;
        RECT 1152.400 120.400 1152.660 120.660 ;
      LAYER met2 ;
        RECT 1032.690 960.570 1032.970 964.000 ;
        RECT 1032.690 960.430 1034.380 960.570 ;
        RECT 1032.690 960.000 1032.970 960.430 ;
        RECT 1034.240 120.690 1034.380 960.430 ;
        RECT 1034.180 120.370 1034.440 120.690 ;
        RECT 1152.400 120.370 1152.660 120.690 ;
        RECT 1152.460 17.410 1152.600 120.370 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 17.240 674.750 17.300 ;
        RECT 696.970 17.240 697.290 17.300 ;
        RECT 674.430 17.100 697.290 17.240 ;
        RECT 674.430 17.040 674.750 17.100 ;
        RECT 696.970 17.040 697.290 17.100 ;
      LAYER via ;
        RECT 674.460 17.040 674.720 17.300 ;
        RECT 697.000 17.040 697.260 17.300 ;
      LAYER met2 ;
        RECT 698.730 960.570 699.010 964.000 ;
        RECT 697.060 960.430 699.010 960.570 ;
        RECT 697.060 17.330 697.200 960.430 ;
        RECT 698.730 960.000 699.010 960.430 ;
        RECT 674.460 17.010 674.720 17.330 ;
        RECT 697.000 17.010 697.260 17.330 ;
        RECT 674.520 2.400 674.660 17.010 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1048.410 79.800 1048.730 79.860 ;
        RECT 1173.070 79.800 1173.390 79.860 ;
        RECT 1048.410 79.660 1173.390 79.800 ;
        RECT 1048.410 79.600 1048.730 79.660 ;
        RECT 1173.070 79.600 1173.390 79.660 ;
      LAYER via ;
        RECT 1048.440 79.600 1048.700 79.860 ;
        RECT 1173.100 79.600 1173.360 79.860 ;
      LAYER met2 ;
        RECT 1045.110 960.570 1045.390 964.000 ;
        RECT 1045.110 960.430 1048.640 960.570 ;
        RECT 1045.110 960.000 1045.390 960.430 ;
        RECT 1048.500 79.890 1048.640 960.430 ;
        RECT 1048.440 79.570 1048.700 79.890 ;
        RECT 1173.100 79.570 1173.360 79.890 ;
        RECT 1173.160 17.410 1173.300 79.570 ;
        RECT 1173.160 17.270 1174.220 17.410 ;
        RECT 1174.080 2.400 1174.220 17.270 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1057.610 945.440 1057.930 945.500 ;
        RECT 1061.750 945.440 1062.070 945.500 ;
        RECT 1057.610 945.300 1062.070 945.440 ;
        RECT 1057.610 945.240 1057.930 945.300 ;
        RECT 1061.750 945.240 1062.070 945.300 ;
        RECT 1061.750 128.080 1062.070 128.140 ;
        RECT 1186.870 128.080 1187.190 128.140 ;
        RECT 1061.750 127.940 1187.190 128.080 ;
        RECT 1061.750 127.880 1062.070 127.940 ;
        RECT 1186.870 127.880 1187.190 127.940 ;
      LAYER via ;
        RECT 1057.640 945.240 1057.900 945.500 ;
        RECT 1061.780 945.240 1062.040 945.500 ;
        RECT 1061.780 127.880 1062.040 128.140 ;
        RECT 1186.900 127.880 1187.160 128.140 ;
      LAYER met2 ;
        RECT 1057.530 960.500 1057.810 964.000 ;
        RECT 1057.530 960.000 1057.840 960.500 ;
        RECT 1057.700 945.530 1057.840 960.000 ;
        RECT 1057.640 945.210 1057.900 945.530 ;
        RECT 1061.780 945.210 1062.040 945.530 ;
        RECT 1061.840 128.170 1061.980 945.210 ;
        RECT 1061.780 127.850 1062.040 128.170 ;
        RECT 1186.900 127.850 1187.160 128.170 ;
        RECT 1186.960 17.410 1187.100 127.850 ;
        RECT 1186.960 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1070.030 946.800 1070.350 946.860 ;
        RECT 1076.010 946.800 1076.330 946.860 ;
        RECT 1070.030 946.660 1076.330 946.800 ;
        RECT 1070.030 946.600 1070.350 946.660 ;
        RECT 1076.010 946.600 1076.330 946.660 ;
        RECT 1076.010 86.260 1076.330 86.320 ;
        RECT 1207.570 86.260 1207.890 86.320 ;
        RECT 1076.010 86.120 1207.890 86.260 ;
        RECT 1076.010 86.060 1076.330 86.120 ;
        RECT 1207.570 86.060 1207.890 86.120 ;
      LAYER via ;
        RECT 1070.060 946.600 1070.320 946.860 ;
        RECT 1076.040 946.600 1076.300 946.860 ;
        RECT 1076.040 86.060 1076.300 86.320 ;
        RECT 1207.600 86.060 1207.860 86.320 ;
      LAYER met2 ;
        RECT 1069.950 960.500 1070.230 964.000 ;
        RECT 1069.950 960.000 1070.260 960.500 ;
        RECT 1070.120 946.890 1070.260 960.000 ;
        RECT 1070.060 946.570 1070.320 946.890 ;
        RECT 1076.040 946.570 1076.300 946.890 ;
        RECT 1076.100 86.350 1076.240 946.570 ;
        RECT 1076.040 86.030 1076.300 86.350 ;
        RECT 1207.600 86.030 1207.860 86.350 ;
        RECT 1207.660 17.410 1207.800 86.030 ;
        RECT 1207.660 17.270 1210.100 17.410 ;
        RECT 1209.960 2.400 1210.100 17.270 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1082.450 93.060 1082.770 93.120 ;
        RECT 1221.370 93.060 1221.690 93.120 ;
        RECT 1082.450 92.920 1221.690 93.060 ;
        RECT 1082.450 92.860 1082.770 92.920 ;
        RECT 1221.370 92.860 1221.690 92.920 ;
        RECT 1221.370 17.580 1221.690 17.640 ;
        RECT 1227.810 17.580 1228.130 17.640 ;
        RECT 1221.370 17.440 1228.130 17.580 ;
        RECT 1221.370 17.380 1221.690 17.440 ;
        RECT 1227.810 17.380 1228.130 17.440 ;
      LAYER via ;
        RECT 1082.480 92.860 1082.740 93.120 ;
        RECT 1221.400 92.860 1221.660 93.120 ;
        RECT 1221.400 17.380 1221.660 17.640 ;
        RECT 1227.840 17.380 1228.100 17.640 ;
      LAYER met2 ;
        RECT 1082.370 960.500 1082.650 964.000 ;
        RECT 1082.370 960.000 1082.680 960.500 ;
        RECT 1082.540 93.150 1082.680 960.000 ;
        RECT 1082.480 92.830 1082.740 93.150 ;
        RECT 1221.400 92.830 1221.660 93.150 ;
        RECT 1221.460 17.670 1221.600 92.830 ;
        RECT 1221.400 17.350 1221.660 17.670 ;
        RECT 1227.840 17.350 1228.100 17.670 ;
        RECT 1227.900 2.400 1228.040 17.350 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1096.250 99.860 1096.570 99.920 ;
        RECT 1242.070 99.860 1242.390 99.920 ;
        RECT 1096.250 99.720 1242.390 99.860 ;
        RECT 1096.250 99.660 1096.570 99.720 ;
        RECT 1242.070 99.660 1242.390 99.720 ;
      LAYER via ;
        RECT 1096.280 99.660 1096.540 99.920 ;
        RECT 1242.100 99.660 1242.360 99.920 ;
      LAYER met2 ;
        RECT 1094.790 960.570 1095.070 964.000 ;
        RECT 1094.790 960.430 1096.480 960.570 ;
        RECT 1094.790 960.000 1095.070 960.430 ;
        RECT 1096.340 99.950 1096.480 960.430 ;
        RECT 1096.280 99.630 1096.540 99.950 ;
        RECT 1242.100 99.630 1242.360 99.950 ;
        RECT 1242.160 17.410 1242.300 99.630 ;
        RECT 1242.160 17.270 1245.980 17.410 ;
        RECT 1245.840 2.400 1245.980 17.270 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1107.290 946.460 1107.610 946.520 ;
        RECT 1114.190 946.460 1114.510 946.520 ;
        RECT 1107.290 946.320 1114.510 946.460 ;
        RECT 1107.290 946.260 1107.610 946.320 ;
        RECT 1114.190 946.260 1114.510 946.320 ;
        RECT 1114.190 107.000 1114.510 107.060 ;
        RECT 1263.230 107.000 1263.550 107.060 ;
        RECT 1114.190 106.860 1263.550 107.000 ;
        RECT 1114.190 106.800 1114.510 106.860 ;
        RECT 1263.230 106.800 1263.550 106.860 ;
      LAYER via ;
        RECT 1107.320 946.260 1107.580 946.520 ;
        RECT 1114.220 946.260 1114.480 946.520 ;
        RECT 1114.220 106.800 1114.480 107.060 ;
        RECT 1263.260 106.800 1263.520 107.060 ;
      LAYER met2 ;
        RECT 1107.210 960.500 1107.490 964.000 ;
        RECT 1107.210 960.000 1107.520 960.500 ;
        RECT 1107.380 946.550 1107.520 960.000 ;
        RECT 1107.320 946.230 1107.580 946.550 ;
        RECT 1114.220 946.230 1114.480 946.550 ;
        RECT 1114.280 107.090 1114.420 946.230 ;
        RECT 1114.220 106.770 1114.480 107.090 ;
        RECT 1263.260 106.770 1263.520 107.090 ;
        RECT 1263.320 2.400 1263.460 106.770 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1119.250 946.460 1119.570 946.520 ;
        RECT 1124.310 946.460 1124.630 946.520 ;
        RECT 1119.250 946.320 1124.630 946.460 ;
        RECT 1119.250 946.260 1119.570 946.320 ;
        RECT 1124.310 946.260 1124.630 946.320 ;
        RECT 1124.310 134.540 1124.630 134.600 ;
        RECT 1276.570 134.540 1276.890 134.600 ;
        RECT 1124.310 134.400 1276.890 134.540 ;
        RECT 1124.310 134.340 1124.630 134.400 ;
        RECT 1276.570 134.340 1276.890 134.400 ;
      LAYER via ;
        RECT 1119.280 946.260 1119.540 946.520 ;
        RECT 1124.340 946.260 1124.600 946.520 ;
        RECT 1124.340 134.340 1124.600 134.600 ;
        RECT 1276.600 134.340 1276.860 134.600 ;
      LAYER met2 ;
        RECT 1119.170 960.500 1119.450 964.000 ;
        RECT 1119.170 960.000 1119.480 960.500 ;
        RECT 1119.340 946.550 1119.480 960.000 ;
        RECT 1119.280 946.230 1119.540 946.550 ;
        RECT 1124.340 946.230 1124.600 946.550 ;
        RECT 1124.400 134.630 1124.540 946.230 ;
        RECT 1124.340 134.310 1124.600 134.630 ;
        RECT 1276.600 134.310 1276.860 134.630 ;
        RECT 1276.660 18.090 1276.800 134.310 ;
        RECT 1276.660 17.950 1281.400 18.090 ;
        RECT 1281.260 2.400 1281.400 17.950 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1131.670 950.200 1131.990 950.260 ;
        RECT 1137.650 950.200 1137.970 950.260 ;
        RECT 1131.670 950.060 1137.970 950.200 ;
        RECT 1131.670 950.000 1131.990 950.060 ;
        RECT 1137.650 950.000 1137.970 950.060 ;
        RECT 1137.650 886.620 1137.970 886.680 ;
        RECT 1297.270 886.620 1297.590 886.680 ;
        RECT 1137.650 886.480 1297.590 886.620 ;
        RECT 1137.650 886.420 1137.970 886.480 ;
        RECT 1297.270 886.420 1297.590 886.480 ;
      LAYER via ;
        RECT 1131.700 950.000 1131.960 950.260 ;
        RECT 1137.680 950.000 1137.940 950.260 ;
        RECT 1137.680 886.420 1137.940 886.680 ;
        RECT 1297.300 886.420 1297.560 886.680 ;
      LAYER met2 ;
        RECT 1131.590 960.500 1131.870 964.000 ;
        RECT 1131.590 960.000 1131.900 960.500 ;
        RECT 1131.760 950.290 1131.900 960.000 ;
        RECT 1131.700 949.970 1131.960 950.290 ;
        RECT 1137.680 949.970 1137.940 950.290 ;
        RECT 1137.740 886.710 1137.880 949.970 ;
        RECT 1137.680 886.390 1137.940 886.710 ;
        RECT 1297.300 886.390 1297.560 886.710 ;
        RECT 1297.360 17.410 1297.500 886.390 ;
        RECT 1297.360 17.270 1299.340 17.410 ;
        RECT 1299.200 2.400 1299.340 17.270 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1144.550 113.800 1144.870 113.860 ;
        RECT 1311.070 113.800 1311.390 113.860 ;
        RECT 1144.550 113.660 1311.390 113.800 ;
        RECT 1144.550 113.600 1144.870 113.660 ;
        RECT 1311.070 113.600 1311.390 113.660 ;
        RECT 1311.070 17.920 1311.390 17.980 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1311.070 17.780 1317.370 17.920 ;
        RECT 1311.070 17.720 1311.390 17.780 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
      LAYER via ;
        RECT 1144.580 113.600 1144.840 113.860 ;
        RECT 1311.100 113.600 1311.360 113.860 ;
        RECT 1311.100 17.720 1311.360 17.980 ;
        RECT 1317.080 17.720 1317.340 17.980 ;
      LAYER met2 ;
        RECT 1144.010 960.570 1144.290 964.000 ;
        RECT 1144.010 960.430 1144.780 960.570 ;
        RECT 1144.010 960.000 1144.290 960.430 ;
        RECT 1144.640 113.890 1144.780 960.430 ;
        RECT 1144.580 113.570 1144.840 113.890 ;
        RECT 1311.100 113.570 1311.360 113.890 ;
        RECT 1311.160 18.010 1311.300 113.570 ;
        RECT 1311.100 17.690 1311.360 18.010 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1317.140 2.400 1317.280 17.690 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.350 120.600 1158.670 120.660 ;
        RECT 1331.770 120.600 1332.090 120.660 ;
        RECT 1158.350 120.460 1332.090 120.600 ;
        RECT 1158.350 120.400 1158.670 120.460 ;
        RECT 1331.770 120.400 1332.090 120.460 ;
      LAYER via ;
        RECT 1158.380 120.400 1158.640 120.660 ;
        RECT 1331.800 120.400 1332.060 120.660 ;
      LAYER met2 ;
        RECT 1156.430 960.570 1156.710 964.000 ;
        RECT 1156.430 960.430 1158.580 960.570 ;
        RECT 1156.430 960.000 1156.710 960.430 ;
        RECT 1158.440 120.690 1158.580 960.430 ;
        RECT 1158.380 120.370 1158.640 120.690 ;
        RECT 1331.800 120.370 1332.060 120.690 ;
        RECT 1331.860 17.410 1332.000 120.370 ;
        RECT 1331.860 17.270 1335.220 17.410 ;
        RECT 1335.080 2.400 1335.220 17.270 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 17.920 692.690 17.980 ;
        RECT 711.230 17.920 711.550 17.980 ;
        RECT 692.370 17.780 711.550 17.920 ;
        RECT 692.370 17.720 692.690 17.780 ;
        RECT 711.230 17.720 711.550 17.780 ;
      LAYER via ;
        RECT 692.400 17.720 692.660 17.980 ;
        RECT 711.260 17.720 711.520 17.980 ;
      LAYER met2 ;
        RECT 711.150 960.500 711.430 964.000 ;
        RECT 711.150 960.000 711.460 960.500 ;
        RECT 711.320 18.010 711.460 960.000 ;
        RECT 692.400 17.690 692.660 18.010 ;
        RECT 711.260 17.690 711.520 18.010 ;
        RECT 692.460 2.400 692.600 17.690 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 141.340 1172.930 141.400 ;
        RECT 1352.930 141.340 1353.250 141.400 ;
        RECT 1172.610 141.200 1353.250 141.340 ;
        RECT 1172.610 141.140 1172.930 141.200 ;
        RECT 1352.930 141.140 1353.250 141.200 ;
      LAYER via ;
        RECT 1172.640 141.140 1172.900 141.400 ;
        RECT 1352.960 141.140 1353.220 141.400 ;
      LAYER met2 ;
        RECT 1168.850 960.570 1169.130 964.000 ;
        RECT 1168.850 960.430 1172.840 960.570 ;
        RECT 1168.850 960.000 1169.130 960.430 ;
        RECT 1172.700 141.430 1172.840 960.430 ;
        RECT 1172.640 141.110 1172.900 141.430 ;
        RECT 1352.960 141.110 1353.220 141.430 ;
        RECT 1353.020 17.410 1353.160 141.110 ;
        RECT 1352.560 17.270 1353.160 17.410 ;
        RECT 1352.560 2.400 1352.700 17.270 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 946.800 1181.670 946.860 ;
        RECT 1186.410 946.800 1186.730 946.860 ;
        RECT 1181.350 946.660 1186.730 946.800 ;
        RECT 1181.350 946.600 1181.670 946.660 ;
        RECT 1186.410 946.600 1186.730 946.660 ;
        RECT 1186.410 127.740 1186.730 127.800 ;
        RECT 1366.270 127.740 1366.590 127.800 ;
        RECT 1186.410 127.600 1366.590 127.740 ;
        RECT 1186.410 127.540 1186.730 127.600 ;
        RECT 1366.270 127.540 1366.590 127.600 ;
      LAYER via ;
        RECT 1181.380 946.600 1181.640 946.860 ;
        RECT 1186.440 946.600 1186.700 946.860 ;
        RECT 1186.440 127.540 1186.700 127.800 ;
        RECT 1366.300 127.540 1366.560 127.800 ;
      LAYER met2 ;
        RECT 1181.270 960.500 1181.550 964.000 ;
        RECT 1181.270 960.000 1181.580 960.500 ;
        RECT 1181.440 946.890 1181.580 960.000 ;
        RECT 1181.380 946.570 1181.640 946.890 ;
        RECT 1186.440 946.570 1186.700 946.890 ;
        RECT 1186.500 127.830 1186.640 946.570 ;
        RECT 1186.440 127.510 1186.700 127.830 ;
        RECT 1366.300 127.510 1366.560 127.830 ;
        RECT 1366.360 17.410 1366.500 127.510 ;
        RECT 1366.360 17.270 1370.640 17.410 ;
        RECT 1370.500 2.400 1370.640 17.270 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.770 946.460 1194.090 946.520 ;
        RECT 1200.210 946.460 1200.530 946.520 ;
        RECT 1193.770 946.320 1200.530 946.460 ;
        RECT 1193.770 946.260 1194.090 946.320 ;
        RECT 1200.210 946.260 1200.530 946.320 ;
        RECT 1200.210 148.140 1200.530 148.200 ;
        RECT 1386.970 148.140 1387.290 148.200 ;
        RECT 1200.210 148.000 1387.290 148.140 ;
        RECT 1200.210 147.940 1200.530 148.000 ;
        RECT 1386.970 147.940 1387.290 148.000 ;
      LAYER via ;
        RECT 1193.800 946.260 1194.060 946.520 ;
        RECT 1200.240 946.260 1200.500 946.520 ;
        RECT 1200.240 147.940 1200.500 148.200 ;
        RECT 1387.000 147.940 1387.260 148.200 ;
      LAYER met2 ;
        RECT 1193.690 960.500 1193.970 964.000 ;
        RECT 1193.690 960.000 1194.000 960.500 ;
        RECT 1193.860 946.550 1194.000 960.000 ;
        RECT 1193.800 946.230 1194.060 946.550 ;
        RECT 1200.240 946.230 1200.500 946.550 ;
        RECT 1200.300 148.230 1200.440 946.230 ;
        RECT 1200.240 147.910 1200.500 148.230 ;
        RECT 1387.000 147.910 1387.260 148.230 ;
        RECT 1387.060 16.730 1387.200 147.910 ;
        RECT 1387.060 16.590 1388.580 16.730 ;
        RECT 1388.440 2.400 1388.580 16.590 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.110 155.280 1207.430 155.340 ;
        RECT 1400.770 155.280 1401.090 155.340 ;
        RECT 1207.110 155.140 1401.090 155.280 ;
        RECT 1207.110 155.080 1207.430 155.140 ;
        RECT 1400.770 155.080 1401.090 155.140 ;
      LAYER via ;
        RECT 1207.140 155.080 1207.400 155.340 ;
        RECT 1400.800 155.080 1401.060 155.340 ;
      LAYER met2 ;
        RECT 1206.110 960.570 1206.390 964.000 ;
        RECT 1206.110 960.430 1207.340 960.570 ;
        RECT 1206.110 960.000 1206.390 960.430 ;
        RECT 1207.200 155.370 1207.340 960.430 ;
        RECT 1207.140 155.050 1207.400 155.370 ;
        RECT 1400.800 155.050 1401.060 155.370 ;
        RECT 1400.860 16.730 1401.000 155.050 ;
        RECT 1400.860 16.590 1406.520 16.730 ;
        RECT 1406.380 2.400 1406.520 16.590 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.450 162.080 1220.770 162.140 ;
        RECT 1421.470 162.080 1421.790 162.140 ;
        RECT 1220.450 161.940 1421.790 162.080 ;
        RECT 1220.450 161.880 1220.770 161.940 ;
        RECT 1421.470 161.880 1421.790 161.940 ;
      LAYER via ;
        RECT 1220.480 161.880 1220.740 162.140 ;
        RECT 1421.500 161.880 1421.760 162.140 ;
      LAYER met2 ;
        RECT 1218.530 960.570 1218.810 964.000 ;
        RECT 1218.530 960.430 1220.680 960.570 ;
        RECT 1218.530 960.000 1218.810 960.430 ;
        RECT 1220.540 162.170 1220.680 960.430 ;
        RECT 1220.480 161.850 1220.740 162.170 ;
        RECT 1421.500 161.850 1421.760 162.170 ;
        RECT 1421.560 16.730 1421.700 161.850 ;
        RECT 1421.560 16.590 1424.000 16.730 ;
        RECT 1423.860 2.400 1424.000 16.590 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1230.570 945.440 1230.890 945.500 ;
        RECT 1234.710 945.440 1235.030 945.500 ;
        RECT 1230.570 945.300 1235.030 945.440 ;
        RECT 1230.570 945.240 1230.890 945.300 ;
        RECT 1234.710 945.240 1235.030 945.300 ;
        RECT 1234.710 169.220 1235.030 169.280 ;
        RECT 1435.270 169.220 1435.590 169.280 ;
        RECT 1234.710 169.080 1435.590 169.220 ;
        RECT 1234.710 169.020 1235.030 169.080 ;
        RECT 1435.270 169.020 1435.590 169.080 ;
        RECT 1435.270 17.580 1435.590 17.640 ;
        RECT 1441.710 17.580 1442.030 17.640 ;
        RECT 1435.270 17.440 1442.030 17.580 ;
        RECT 1435.270 17.380 1435.590 17.440 ;
        RECT 1441.710 17.380 1442.030 17.440 ;
      LAYER via ;
        RECT 1230.600 945.240 1230.860 945.500 ;
        RECT 1234.740 945.240 1235.000 945.500 ;
        RECT 1234.740 169.020 1235.000 169.280 ;
        RECT 1435.300 169.020 1435.560 169.280 ;
        RECT 1435.300 17.380 1435.560 17.640 ;
        RECT 1441.740 17.380 1442.000 17.640 ;
      LAYER met2 ;
        RECT 1230.490 960.500 1230.770 964.000 ;
        RECT 1230.490 960.000 1230.800 960.500 ;
        RECT 1230.660 945.530 1230.800 960.000 ;
        RECT 1230.600 945.210 1230.860 945.530 ;
        RECT 1234.740 945.210 1235.000 945.530 ;
        RECT 1234.800 169.310 1234.940 945.210 ;
        RECT 1234.740 168.990 1235.000 169.310 ;
        RECT 1435.300 168.990 1435.560 169.310 ;
        RECT 1435.360 17.670 1435.500 168.990 ;
        RECT 1435.300 17.350 1435.560 17.670 ;
        RECT 1441.740 17.350 1442.000 17.670 ;
        RECT 1441.800 2.400 1441.940 17.350 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1242.990 946.460 1243.310 946.520 ;
        RECT 1248.510 946.460 1248.830 946.520 ;
        RECT 1242.990 946.320 1248.830 946.460 ;
        RECT 1242.990 946.260 1243.310 946.320 ;
        RECT 1248.510 946.260 1248.830 946.320 ;
        RECT 1248.510 176.020 1248.830 176.080 ;
        RECT 1455.970 176.020 1456.290 176.080 ;
        RECT 1248.510 175.880 1456.290 176.020 ;
        RECT 1248.510 175.820 1248.830 175.880 ;
        RECT 1455.970 175.820 1456.290 175.880 ;
      LAYER via ;
        RECT 1243.020 946.260 1243.280 946.520 ;
        RECT 1248.540 946.260 1248.800 946.520 ;
        RECT 1248.540 175.820 1248.800 176.080 ;
        RECT 1456.000 175.820 1456.260 176.080 ;
      LAYER met2 ;
        RECT 1242.910 960.500 1243.190 964.000 ;
        RECT 1242.910 960.000 1243.220 960.500 ;
        RECT 1243.080 946.550 1243.220 960.000 ;
        RECT 1243.020 946.230 1243.280 946.550 ;
        RECT 1248.540 946.230 1248.800 946.550 ;
        RECT 1248.600 176.110 1248.740 946.230 ;
        RECT 1248.540 175.790 1248.800 176.110 ;
        RECT 1456.000 175.790 1456.260 176.110 ;
        RECT 1456.060 17.410 1456.200 175.790 ;
        RECT 1456.060 17.270 1459.880 17.410 ;
        RECT 1459.740 2.400 1459.880 17.270 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1254.950 182.820 1255.270 182.880 ;
        RECT 1476.670 182.820 1476.990 182.880 ;
        RECT 1254.950 182.680 1476.990 182.820 ;
        RECT 1254.950 182.620 1255.270 182.680 ;
        RECT 1476.670 182.620 1476.990 182.680 ;
      LAYER via ;
        RECT 1254.980 182.620 1255.240 182.880 ;
        RECT 1476.700 182.620 1476.960 182.880 ;
      LAYER met2 ;
        RECT 1255.330 960.570 1255.610 964.000 ;
        RECT 1255.040 960.430 1255.610 960.570 ;
        RECT 1255.040 182.910 1255.180 960.430 ;
        RECT 1255.330 960.000 1255.610 960.430 ;
        RECT 1254.980 182.590 1255.240 182.910 ;
        RECT 1476.700 182.590 1476.960 182.910 ;
        RECT 1476.760 17.410 1476.900 182.590 ;
        RECT 1476.760 17.270 1477.820 17.410 ;
        RECT 1477.680 2.400 1477.820 17.270 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1267.830 950.540 1268.150 950.600 ;
        RECT 1286.690 950.540 1287.010 950.600 ;
        RECT 1267.830 950.400 1287.010 950.540 ;
        RECT 1267.830 950.340 1268.150 950.400 ;
        RECT 1286.690 950.340 1287.010 950.400 ;
        RECT 1286.690 134.540 1287.010 134.600 ;
        RECT 1490.470 134.540 1490.790 134.600 ;
        RECT 1286.690 134.400 1490.790 134.540 ;
        RECT 1286.690 134.340 1287.010 134.400 ;
        RECT 1490.470 134.340 1490.790 134.400 ;
      LAYER via ;
        RECT 1267.860 950.340 1268.120 950.600 ;
        RECT 1286.720 950.340 1286.980 950.600 ;
        RECT 1286.720 134.340 1286.980 134.600 ;
        RECT 1490.500 134.340 1490.760 134.600 ;
      LAYER met2 ;
        RECT 1267.750 960.500 1268.030 964.000 ;
        RECT 1267.750 960.000 1268.060 960.500 ;
        RECT 1267.920 950.630 1268.060 960.000 ;
        RECT 1267.860 950.310 1268.120 950.630 ;
        RECT 1286.720 950.310 1286.980 950.630 ;
        RECT 1286.780 134.630 1286.920 950.310 ;
        RECT 1286.720 134.310 1286.980 134.630 ;
        RECT 1490.500 134.310 1490.760 134.630 ;
        RECT 1490.560 17.410 1490.700 134.310 ;
        RECT 1490.560 17.270 1495.760 17.410 ;
        RECT 1495.620 2.400 1495.760 17.270 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 189.620 1283.330 189.680 ;
        RECT 1511.170 189.620 1511.490 189.680 ;
        RECT 1283.010 189.480 1511.490 189.620 ;
        RECT 1283.010 189.420 1283.330 189.480 ;
        RECT 1511.170 189.420 1511.490 189.480 ;
      LAYER via ;
        RECT 1283.040 189.420 1283.300 189.680 ;
        RECT 1511.200 189.420 1511.460 189.680 ;
      LAYER met2 ;
        RECT 1280.170 960.570 1280.450 964.000 ;
        RECT 1280.170 960.430 1283.240 960.570 ;
        RECT 1280.170 960.000 1280.450 960.430 ;
        RECT 1283.100 189.710 1283.240 960.430 ;
        RECT 1283.040 189.390 1283.300 189.710 ;
        RECT 1511.200 189.390 1511.460 189.710 ;
        RECT 1511.260 17.410 1511.400 189.390 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 719.125 641.325 719.295 717.655 ;
        RECT 718.205 386.325 718.375 434.775 ;
        RECT 718.665 241.485 718.835 289.595 ;
      LAYER mcon ;
        RECT 719.125 717.485 719.295 717.655 ;
        RECT 718.205 434.605 718.375 434.775 ;
        RECT 718.665 289.425 718.835 289.595 ;
      LAYER met1 ;
        RECT 719.510 869.620 719.830 869.680 ;
        RECT 720.890 869.620 721.210 869.680 ;
        RECT 719.510 869.480 721.210 869.620 ;
        RECT 719.510 869.420 719.830 869.480 ;
        RECT 720.890 869.420 721.210 869.480 ;
        RECT 718.130 821.000 718.450 821.060 ;
        RECT 719.050 821.000 719.370 821.060 ;
        RECT 718.130 820.860 719.370 821.000 ;
        RECT 718.130 820.800 718.450 820.860 ;
        RECT 719.050 820.800 719.370 820.860 ;
        RECT 719.050 717.640 719.370 717.700 ;
        RECT 718.855 717.500 719.370 717.640 ;
        RECT 719.050 717.440 719.370 717.500 ;
        RECT 719.050 641.480 719.370 641.540 ;
        RECT 718.855 641.340 719.370 641.480 ;
        RECT 719.050 641.280 719.370 641.340 ;
        RECT 718.145 434.760 718.435 434.805 ;
        RECT 718.590 434.760 718.910 434.820 ;
        RECT 718.145 434.620 718.910 434.760 ;
        RECT 718.145 434.575 718.435 434.620 ;
        RECT 718.590 434.560 718.910 434.620 ;
        RECT 718.130 386.480 718.450 386.540 ;
        RECT 717.935 386.340 718.450 386.480 ;
        RECT 718.130 386.280 718.450 386.340 ;
        RECT 718.590 303.520 718.910 303.580 ;
        RECT 719.510 303.520 719.830 303.580 ;
        RECT 718.590 303.380 719.830 303.520 ;
        RECT 718.590 303.320 718.910 303.380 ;
        RECT 719.510 303.320 719.830 303.380 ;
        RECT 718.605 289.580 718.895 289.625 ;
        RECT 719.510 289.580 719.830 289.640 ;
        RECT 718.605 289.440 719.830 289.580 ;
        RECT 718.605 289.395 718.895 289.440 ;
        RECT 719.510 289.380 719.830 289.440 ;
        RECT 718.590 241.640 718.910 241.700 ;
        RECT 718.395 241.500 718.910 241.640 ;
        RECT 718.590 241.440 718.910 241.500 ;
        RECT 718.590 193.360 718.910 193.420 ;
        RECT 719.510 193.360 719.830 193.420 ;
        RECT 718.590 193.220 719.830 193.360 ;
        RECT 718.590 193.160 718.910 193.220 ;
        RECT 719.510 193.160 719.830 193.220 ;
        RECT 718.590 137.940 718.910 138.000 ;
        RECT 719.970 137.940 720.290 138.000 ;
        RECT 718.590 137.800 720.290 137.940 ;
        RECT 718.590 137.740 718.910 137.800 ;
        RECT 719.970 137.740 720.290 137.800 ;
        RECT 710.310 19.280 710.630 19.340 ;
        RECT 719.510 19.280 719.830 19.340 ;
        RECT 710.310 19.140 719.830 19.280 ;
        RECT 710.310 19.080 710.630 19.140 ;
        RECT 719.510 19.080 719.830 19.140 ;
      LAYER via ;
        RECT 719.540 869.420 719.800 869.680 ;
        RECT 720.920 869.420 721.180 869.680 ;
        RECT 718.160 820.800 718.420 821.060 ;
        RECT 719.080 820.800 719.340 821.060 ;
        RECT 719.080 717.440 719.340 717.700 ;
        RECT 719.080 641.280 719.340 641.540 ;
        RECT 718.620 434.560 718.880 434.820 ;
        RECT 718.160 386.280 718.420 386.540 ;
        RECT 718.620 303.320 718.880 303.580 ;
        RECT 719.540 303.320 719.800 303.580 ;
        RECT 719.540 289.380 719.800 289.640 ;
        RECT 718.620 241.440 718.880 241.700 ;
        RECT 718.620 193.160 718.880 193.420 ;
        RECT 719.540 193.160 719.800 193.420 ;
        RECT 718.620 137.740 718.880 138.000 ;
        RECT 720.000 137.740 720.260 138.000 ;
        RECT 710.340 19.080 710.600 19.340 ;
        RECT 719.540 19.080 719.800 19.340 ;
      LAYER met2 ;
        RECT 723.570 960.570 723.850 964.000 ;
        RECT 720.060 960.430 723.850 960.570 ;
        RECT 720.060 917.845 720.200 960.430 ;
        RECT 723.570 960.000 723.850 960.430 ;
        RECT 719.990 917.475 720.270 917.845 ;
        RECT 720.910 917.475 721.190 917.845 ;
        RECT 720.980 869.710 721.120 917.475 ;
        RECT 719.540 869.390 719.800 869.710 ;
        RECT 720.920 869.390 721.180 869.710 ;
        RECT 719.600 834.770 719.740 869.390 ;
        RECT 719.140 834.630 719.740 834.770 ;
        RECT 719.140 821.090 719.280 834.630 ;
        RECT 718.160 820.770 718.420 821.090 ;
        RECT 719.080 820.770 719.340 821.090 ;
        RECT 718.220 773.005 718.360 820.770 ;
        RECT 718.150 772.635 718.430 773.005 ;
        RECT 719.530 772.635 719.810 773.005 ;
        RECT 719.600 738.210 719.740 772.635 ;
        RECT 719.140 738.070 719.740 738.210 ;
        RECT 719.140 717.730 719.280 738.070 ;
        RECT 719.080 717.410 719.340 717.730 ;
        RECT 719.080 641.250 719.340 641.570 ;
        RECT 719.140 603.570 719.280 641.250 ;
        RECT 718.220 603.430 719.280 603.570 ;
        RECT 718.220 579.885 718.360 603.430 ;
        RECT 718.150 579.515 718.430 579.885 ;
        RECT 719.530 579.515 719.810 579.885 ;
        RECT 719.600 545.090 719.740 579.515 ;
        RECT 719.140 544.950 719.740 545.090 ;
        RECT 719.140 507.010 719.280 544.950 ;
        RECT 718.220 506.870 719.280 507.010 ;
        RECT 718.220 483.325 718.360 506.870 ;
        RECT 718.150 482.955 718.430 483.325 ;
        RECT 719.530 482.955 719.810 483.325 ;
        RECT 719.600 448.530 719.740 482.955 ;
        RECT 718.680 448.390 719.740 448.530 ;
        RECT 718.680 434.850 718.820 448.390 ;
        RECT 718.620 434.530 718.880 434.850 ;
        RECT 718.160 386.250 718.420 386.570 ;
        RECT 718.220 351.290 718.360 386.250 ;
        RECT 718.220 351.150 718.820 351.290 ;
        RECT 718.680 303.610 718.820 351.150 ;
        RECT 718.620 303.290 718.880 303.610 ;
        RECT 719.540 303.290 719.800 303.610 ;
        RECT 719.600 289.670 719.740 303.290 ;
        RECT 719.540 289.350 719.800 289.670 ;
        RECT 718.620 241.410 718.880 241.730 ;
        RECT 718.680 193.450 718.820 241.410 ;
        RECT 718.620 193.130 718.880 193.450 ;
        RECT 719.540 193.130 719.800 193.450 ;
        RECT 719.600 145.250 719.740 193.130 ;
        RECT 718.680 145.110 719.740 145.250 ;
        RECT 718.680 138.030 718.820 145.110 ;
        RECT 718.620 137.710 718.880 138.030 ;
        RECT 720.000 137.710 720.260 138.030 ;
        RECT 720.060 62.290 720.200 137.710 ;
        RECT 719.600 62.150 720.200 62.290 ;
        RECT 719.600 19.370 719.740 62.150 ;
        RECT 710.340 19.050 710.600 19.370 ;
        RECT 719.540 19.050 719.800 19.370 ;
        RECT 710.400 2.400 710.540 19.050 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 719.990 917.520 720.270 917.800 ;
        RECT 720.910 917.520 721.190 917.800 ;
        RECT 718.150 772.680 718.430 772.960 ;
        RECT 719.530 772.680 719.810 772.960 ;
        RECT 718.150 579.560 718.430 579.840 ;
        RECT 719.530 579.560 719.810 579.840 ;
        RECT 718.150 483.000 718.430 483.280 ;
        RECT 719.530 483.000 719.810 483.280 ;
      LAYER met3 ;
        RECT 719.965 917.810 720.295 917.825 ;
        RECT 720.885 917.810 721.215 917.825 ;
        RECT 719.965 917.510 721.215 917.810 ;
        RECT 719.965 917.495 720.295 917.510 ;
        RECT 720.885 917.495 721.215 917.510 ;
        RECT 718.125 772.970 718.455 772.985 ;
        RECT 719.505 772.970 719.835 772.985 ;
        RECT 718.125 772.670 719.835 772.970 ;
        RECT 718.125 772.655 718.455 772.670 ;
        RECT 719.505 772.655 719.835 772.670 ;
        RECT 718.125 579.850 718.455 579.865 ;
        RECT 719.505 579.850 719.835 579.865 ;
        RECT 718.125 579.550 719.835 579.850 ;
        RECT 718.125 579.535 718.455 579.550 ;
        RECT 719.505 579.535 719.835 579.550 ;
        RECT 718.125 483.290 718.455 483.305 ;
        RECT 719.505 483.290 719.835 483.305 ;
        RECT 718.125 482.990 719.835 483.290 ;
        RECT 718.125 482.975 718.455 482.990 ;
        RECT 719.505 482.975 719.835 482.990 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1292.670 945.440 1292.990 945.500 ;
        RECT 1296.350 945.440 1296.670 945.500 ;
        RECT 1292.670 945.300 1296.670 945.440 ;
        RECT 1292.670 945.240 1292.990 945.300 ;
        RECT 1296.350 945.240 1296.670 945.300 ;
        RECT 1296.350 893.420 1296.670 893.480 ;
        RECT 1524.970 893.420 1525.290 893.480 ;
        RECT 1296.350 893.280 1525.290 893.420 ;
        RECT 1296.350 893.220 1296.670 893.280 ;
        RECT 1524.970 893.220 1525.290 893.280 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1530.950 17.580 1531.270 17.640 ;
        RECT 1524.970 17.440 1531.270 17.580 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
        RECT 1530.950 17.380 1531.270 17.440 ;
      LAYER via ;
        RECT 1292.700 945.240 1292.960 945.500 ;
        RECT 1296.380 945.240 1296.640 945.500 ;
        RECT 1296.380 893.220 1296.640 893.480 ;
        RECT 1525.000 893.220 1525.260 893.480 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
        RECT 1530.980 17.380 1531.240 17.640 ;
      LAYER met2 ;
        RECT 1292.590 960.500 1292.870 964.000 ;
        RECT 1292.590 960.000 1292.900 960.500 ;
        RECT 1292.760 945.530 1292.900 960.000 ;
        RECT 1292.700 945.210 1292.960 945.530 ;
        RECT 1296.380 945.210 1296.640 945.530 ;
        RECT 1296.440 893.510 1296.580 945.210 ;
        RECT 1296.380 893.190 1296.640 893.510 ;
        RECT 1525.000 893.190 1525.260 893.510 ;
        RECT 1525.060 17.670 1525.200 893.190 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1530.980 17.350 1531.240 17.670 ;
        RECT 1531.040 2.400 1531.180 17.350 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1305.090 946.800 1305.410 946.860 ;
        RECT 1310.610 946.800 1310.930 946.860 ;
        RECT 1305.090 946.660 1310.930 946.800 ;
        RECT 1305.090 946.600 1305.410 946.660 ;
        RECT 1310.610 946.600 1310.930 946.660 ;
        RECT 1310.610 197.100 1310.930 197.160 ;
        RECT 1545.670 197.100 1545.990 197.160 ;
        RECT 1310.610 196.960 1545.990 197.100 ;
        RECT 1310.610 196.900 1310.930 196.960 ;
        RECT 1545.670 196.900 1545.990 196.960 ;
      LAYER via ;
        RECT 1305.120 946.600 1305.380 946.860 ;
        RECT 1310.640 946.600 1310.900 946.860 ;
        RECT 1310.640 196.900 1310.900 197.160 ;
        RECT 1545.700 196.900 1545.960 197.160 ;
      LAYER met2 ;
        RECT 1305.010 960.500 1305.290 964.000 ;
        RECT 1305.010 960.000 1305.320 960.500 ;
        RECT 1305.180 946.890 1305.320 960.000 ;
        RECT 1305.120 946.570 1305.380 946.890 ;
        RECT 1310.640 946.570 1310.900 946.890 ;
        RECT 1310.700 197.190 1310.840 946.570 ;
        RECT 1310.640 196.870 1310.900 197.190 ;
        RECT 1545.700 196.870 1545.960 197.190 ;
        RECT 1545.760 16.730 1545.900 196.870 ;
        RECT 1545.760 16.590 1549.120 16.730 ;
        RECT 1548.980 2.400 1549.120 16.590 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 203.560 1317.370 203.620 ;
        RECT 1566.830 203.560 1567.150 203.620 ;
        RECT 1317.050 203.420 1567.150 203.560 ;
        RECT 1317.050 203.360 1317.370 203.420 ;
        RECT 1566.830 203.360 1567.150 203.420 ;
      LAYER via ;
        RECT 1317.080 203.360 1317.340 203.620 ;
        RECT 1566.860 203.360 1567.120 203.620 ;
      LAYER met2 ;
        RECT 1317.430 960.570 1317.710 964.000 ;
        RECT 1317.140 960.430 1317.710 960.570 ;
        RECT 1317.140 203.650 1317.280 960.430 ;
        RECT 1317.430 960.000 1317.710 960.430 ;
        RECT 1317.080 203.330 1317.340 203.650 ;
        RECT 1566.860 203.330 1567.120 203.650 ;
        RECT 1566.920 2.400 1567.060 203.330 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1330.850 210.700 1331.170 210.760 ;
        RECT 1580.170 210.700 1580.490 210.760 ;
        RECT 1330.850 210.560 1580.490 210.700 ;
        RECT 1330.850 210.500 1331.170 210.560 ;
        RECT 1580.170 210.500 1580.490 210.560 ;
      LAYER via ;
        RECT 1330.880 210.500 1331.140 210.760 ;
        RECT 1580.200 210.500 1580.460 210.760 ;
      LAYER met2 ;
        RECT 1329.850 960.570 1330.130 964.000 ;
        RECT 1329.850 960.430 1331.080 960.570 ;
        RECT 1329.850 960.000 1330.130 960.430 ;
        RECT 1330.940 210.790 1331.080 960.430 ;
        RECT 1330.880 210.470 1331.140 210.790 ;
        RECT 1580.200 210.470 1580.460 210.790 ;
        RECT 1580.260 17.410 1580.400 210.470 ;
        RECT 1580.260 17.270 1585.000 17.410 ;
        RECT 1584.860 2.400 1585.000 17.270 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 217.160 1345.430 217.220 ;
        RECT 1600.870 217.160 1601.190 217.220 ;
        RECT 1345.110 217.020 1601.190 217.160 ;
        RECT 1345.110 216.960 1345.430 217.020 ;
        RECT 1600.870 216.960 1601.190 217.020 ;
      LAYER via ;
        RECT 1345.140 216.960 1345.400 217.220 ;
        RECT 1600.900 216.960 1601.160 217.220 ;
      LAYER met2 ;
        RECT 1342.270 960.570 1342.550 964.000 ;
        RECT 1342.270 960.430 1345.340 960.570 ;
        RECT 1342.270 960.000 1342.550 960.430 ;
        RECT 1345.200 217.250 1345.340 960.430 ;
        RECT 1345.140 216.930 1345.400 217.250 ;
        RECT 1600.900 216.930 1601.160 217.250 ;
        RECT 1600.960 17.410 1601.100 216.930 ;
        RECT 1600.960 17.270 1602.480 17.410 ;
        RECT 1602.340 2.400 1602.480 17.270 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.310 946.460 1354.630 946.520 ;
        RECT 1359.830 946.460 1360.150 946.520 ;
        RECT 1354.310 946.320 1360.150 946.460 ;
        RECT 1354.310 946.260 1354.630 946.320 ;
        RECT 1359.830 946.260 1360.150 946.320 ;
        RECT 1359.830 934.900 1360.150 934.960 ;
        RECT 1614.670 934.900 1614.990 934.960 ;
        RECT 1359.830 934.760 1614.990 934.900 ;
        RECT 1359.830 934.700 1360.150 934.760 ;
        RECT 1614.670 934.700 1614.990 934.760 ;
      LAYER via ;
        RECT 1354.340 946.260 1354.600 946.520 ;
        RECT 1359.860 946.260 1360.120 946.520 ;
        RECT 1359.860 934.700 1360.120 934.960 ;
        RECT 1614.700 934.700 1614.960 934.960 ;
      LAYER met2 ;
        RECT 1354.230 960.500 1354.510 964.000 ;
        RECT 1354.230 960.000 1354.540 960.500 ;
        RECT 1354.400 946.550 1354.540 960.000 ;
        RECT 1354.340 946.230 1354.600 946.550 ;
        RECT 1359.860 946.230 1360.120 946.550 ;
        RECT 1359.920 934.990 1360.060 946.230 ;
        RECT 1359.860 934.670 1360.120 934.990 ;
        RECT 1614.700 934.670 1614.960 934.990 ;
        RECT 1614.760 17.410 1614.900 934.670 ;
        RECT 1614.760 17.270 1620.420 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1366.730 945.440 1367.050 945.500 ;
        RECT 1372.710 945.440 1373.030 945.500 ;
        RECT 1366.730 945.300 1373.030 945.440 ;
        RECT 1366.730 945.240 1367.050 945.300 ;
        RECT 1372.710 945.240 1373.030 945.300 ;
        RECT 1372.710 224.640 1373.030 224.700 ;
        RECT 1635.370 224.640 1635.690 224.700 ;
        RECT 1372.710 224.500 1635.690 224.640 ;
        RECT 1372.710 224.440 1373.030 224.500 ;
        RECT 1635.370 224.440 1635.690 224.500 ;
      LAYER via ;
        RECT 1366.760 945.240 1367.020 945.500 ;
        RECT 1372.740 945.240 1373.000 945.500 ;
        RECT 1372.740 224.440 1373.000 224.700 ;
        RECT 1635.400 224.440 1635.660 224.700 ;
      LAYER met2 ;
        RECT 1366.650 960.500 1366.930 964.000 ;
        RECT 1366.650 960.000 1366.960 960.500 ;
        RECT 1366.820 945.530 1366.960 960.000 ;
        RECT 1366.760 945.210 1367.020 945.530 ;
        RECT 1372.740 945.210 1373.000 945.530 ;
        RECT 1372.800 224.730 1372.940 945.210 ;
        RECT 1372.740 224.410 1373.000 224.730 ;
        RECT 1635.400 224.410 1635.660 224.730 ;
        RECT 1635.460 17.410 1635.600 224.410 ;
        RECT 1635.460 17.270 1638.360 17.410 ;
        RECT 1638.220 2.400 1638.360 17.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1379.610 237.900 1379.930 237.960 ;
        RECT 1656.530 237.900 1656.850 237.960 ;
        RECT 1379.610 237.760 1656.850 237.900 ;
        RECT 1379.610 237.700 1379.930 237.760 ;
        RECT 1656.530 237.700 1656.850 237.760 ;
      LAYER via ;
        RECT 1379.640 237.700 1379.900 237.960 ;
        RECT 1656.560 237.700 1656.820 237.960 ;
      LAYER met2 ;
        RECT 1379.070 960.570 1379.350 964.000 ;
        RECT 1379.070 960.430 1379.840 960.570 ;
        RECT 1379.070 960.000 1379.350 960.430 ;
        RECT 1379.700 237.990 1379.840 960.430 ;
        RECT 1379.640 237.670 1379.900 237.990 ;
        RECT 1656.560 237.670 1656.820 237.990 ;
        RECT 1656.620 17.410 1656.760 237.670 ;
        RECT 1656.160 17.270 1656.760 17.410 ;
        RECT 1656.160 2.400 1656.300 17.270 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1392.950 231.100 1393.270 231.160 ;
        RECT 1669.870 231.100 1670.190 231.160 ;
        RECT 1392.950 230.960 1670.190 231.100 ;
        RECT 1392.950 230.900 1393.270 230.960 ;
        RECT 1669.870 230.900 1670.190 230.960 ;
      LAYER via ;
        RECT 1392.980 230.900 1393.240 231.160 ;
        RECT 1669.900 230.900 1670.160 231.160 ;
      LAYER met2 ;
        RECT 1391.490 960.570 1391.770 964.000 ;
        RECT 1391.490 960.430 1393.180 960.570 ;
        RECT 1391.490 960.000 1391.770 960.430 ;
        RECT 1393.040 231.190 1393.180 960.430 ;
        RECT 1392.980 230.870 1393.240 231.190 ;
        RECT 1669.900 230.870 1670.160 231.190 ;
        RECT 1669.960 17.410 1670.100 230.870 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 155.280 1407.530 155.340 ;
        RECT 1690.570 155.280 1690.890 155.340 ;
        RECT 1407.210 155.140 1690.890 155.280 ;
        RECT 1407.210 155.080 1407.530 155.140 ;
        RECT 1690.570 155.080 1690.890 155.140 ;
      LAYER via ;
        RECT 1407.240 155.080 1407.500 155.340 ;
        RECT 1690.600 155.080 1690.860 155.340 ;
      LAYER met2 ;
        RECT 1403.910 960.570 1404.190 964.000 ;
        RECT 1403.910 960.430 1407.440 960.570 ;
        RECT 1403.910 960.000 1404.190 960.430 ;
        RECT 1407.300 155.370 1407.440 960.430 ;
        RECT 1407.240 155.050 1407.500 155.370 ;
        RECT 1690.600 155.050 1690.860 155.370 ;
        RECT 1690.660 17.410 1690.800 155.050 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 731.470 904.640 731.790 904.700 ;
        RECT 734.230 904.640 734.550 904.700 ;
        RECT 731.470 904.500 734.550 904.640 ;
        RECT 731.470 904.440 731.790 904.500 ;
        RECT 734.230 904.440 734.550 904.500 ;
        RECT 728.250 16.560 728.570 16.620 ;
        RECT 731.470 16.560 731.790 16.620 ;
        RECT 728.250 16.420 731.790 16.560 ;
        RECT 728.250 16.360 728.570 16.420 ;
        RECT 731.470 16.360 731.790 16.420 ;
      LAYER via ;
        RECT 731.500 904.440 731.760 904.700 ;
        RECT 734.260 904.440 734.520 904.700 ;
        RECT 728.280 16.360 728.540 16.620 ;
        RECT 731.500 16.360 731.760 16.620 ;
      LAYER met2 ;
        RECT 735.990 960.570 736.270 964.000 ;
        RECT 734.320 960.430 736.270 960.570 ;
        RECT 734.320 904.730 734.460 960.430 ;
        RECT 735.990 960.000 736.270 960.430 ;
        RECT 731.500 904.410 731.760 904.730 ;
        RECT 734.260 904.410 734.520 904.730 ;
        RECT 731.560 16.650 731.700 904.410 ;
        RECT 728.280 16.330 728.540 16.650 ;
        RECT 731.500 16.330 731.760 16.650 ;
        RECT 728.340 2.400 728.480 16.330 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1416.410 947.140 1416.730 947.200 ;
        RECT 1421.010 947.140 1421.330 947.200 ;
        RECT 1416.410 947.000 1421.330 947.140 ;
        RECT 1416.410 946.940 1416.730 947.000 ;
        RECT 1421.010 946.940 1421.330 947.000 ;
        RECT 1421.010 245.040 1421.330 245.100 ;
        RECT 1704.370 245.040 1704.690 245.100 ;
        RECT 1421.010 244.900 1704.690 245.040 ;
        RECT 1421.010 244.840 1421.330 244.900 ;
        RECT 1704.370 244.840 1704.690 244.900 ;
      LAYER via ;
        RECT 1416.440 946.940 1416.700 947.200 ;
        RECT 1421.040 946.940 1421.300 947.200 ;
        RECT 1421.040 244.840 1421.300 245.100 ;
        RECT 1704.400 244.840 1704.660 245.100 ;
      LAYER met2 ;
        RECT 1416.330 960.500 1416.610 964.000 ;
        RECT 1416.330 960.000 1416.640 960.500 ;
        RECT 1416.500 947.230 1416.640 960.000 ;
        RECT 1416.440 946.910 1416.700 947.230 ;
        RECT 1421.040 946.910 1421.300 947.230 ;
        RECT 1421.100 245.130 1421.240 946.910 ;
        RECT 1421.040 244.810 1421.300 245.130 ;
        RECT 1704.400 244.810 1704.660 245.130 ;
        RECT 1704.460 17.410 1704.600 244.810 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1428.830 947.480 1429.150 947.540 ;
        RECT 1434.810 947.480 1435.130 947.540 ;
        RECT 1428.830 947.340 1435.130 947.480 ;
        RECT 1428.830 947.280 1429.150 947.340 ;
        RECT 1434.810 947.280 1435.130 947.340 ;
        RECT 1434.810 168.880 1435.130 168.940 ;
        RECT 1725.070 168.880 1725.390 168.940 ;
        RECT 1434.810 168.740 1725.390 168.880 ;
        RECT 1434.810 168.680 1435.130 168.740 ;
        RECT 1725.070 168.680 1725.390 168.740 ;
      LAYER via ;
        RECT 1428.860 947.280 1429.120 947.540 ;
        RECT 1434.840 947.280 1435.100 947.540 ;
        RECT 1434.840 168.680 1435.100 168.940 ;
        RECT 1725.100 168.680 1725.360 168.940 ;
      LAYER met2 ;
        RECT 1428.750 960.500 1429.030 964.000 ;
        RECT 1428.750 960.000 1429.060 960.500 ;
        RECT 1428.920 947.570 1429.060 960.000 ;
        RECT 1428.860 947.250 1429.120 947.570 ;
        RECT 1434.840 947.250 1435.100 947.570 ;
        RECT 1434.900 168.970 1435.040 947.250 ;
        RECT 1434.840 168.650 1435.100 168.970 ;
        RECT 1725.100 168.650 1725.360 168.970 ;
        RECT 1725.160 17.410 1725.300 168.650 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.250 252.180 1441.570 252.240 ;
        RECT 1738.870 252.180 1739.190 252.240 ;
        RECT 1441.250 252.040 1739.190 252.180 ;
        RECT 1441.250 251.980 1441.570 252.040 ;
        RECT 1738.870 251.980 1739.190 252.040 ;
        RECT 1738.870 17.580 1739.190 17.640 ;
        RECT 1745.310 17.580 1745.630 17.640 ;
        RECT 1738.870 17.440 1745.630 17.580 ;
        RECT 1738.870 17.380 1739.190 17.440 ;
        RECT 1745.310 17.380 1745.630 17.440 ;
      LAYER via ;
        RECT 1441.280 251.980 1441.540 252.240 ;
        RECT 1738.900 251.980 1739.160 252.240 ;
        RECT 1738.900 17.380 1739.160 17.640 ;
        RECT 1745.340 17.380 1745.600 17.640 ;
      LAYER met2 ;
        RECT 1441.170 960.500 1441.450 964.000 ;
        RECT 1441.170 960.000 1441.480 960.500 ;
        RECT 1441.340 252.270 1441.480 960.000 ;
        RECT 1441.280 251.950 1441.540 252.270 ;
        RECT 1738.900 251.950 1739.160 252.270 ;
        RECT 1738.960 17.670 1739.100 251.950 ;
        RECT 1738.900 17.350 1739.160 17.670 ;
        RECT 1745.340 17.350 1745.600 17.670 ;
        RECT 1745.400 2.400 1745.540 17.350 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1455.050 258.980 1455.370 259.040 ;
        RECT 1759.570 258.980 1759.890 259.040 ;
        RECT 1455.050 258.840 1759.890 258.980 ;
        RECT 1455.050 258.780 1455.370 258.840 ;
        RECT 1759.570 258.780 1759.890 258.840 ;
      LAYER via ;
        RECT 1455.080 258.780 1455.340 259.040 ;
        RECT 1759.600 258.780 1759.860 259.040 ;
      LAYER met2 ;
        RECT 1453.590 960.570 1453.870 964.000 ;
        RECT 1453.590 960.430 1455.280 960.570 ;
        RECT 1453.590 960.000 1453.870 960.430 ;
        RECT 1455.140 259.070 1455.280 960.430 ;
        RECT 1455.080 258.750 1455.340 259.070 ;
        RECT 1759.600 258.750 1759.860 259.070 ;
        RECT 1759.660 18.090 1759.800 258.750 ;
        RECT 1759.660 17.950 1763.020 18.090 ;
        RECT 1762.880 2.400 1763.020 17.950 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1465.630 945.440 1465.950 945.500 ;
        RECT 1469.310 945.440 1469.630 945.500 ;
        RECT 1465.630 945.300 1469.630 945.440 ;
        RECT 1465.630 945.240 1465.950 945.300 ;
        RECT 1469.310 945.240 1469.630 945.300 ;
        RECT 1469.310 265.440 1469.630 265.500 ;
        RECT 1780.730 265.440 1781.050 265.500 ;
        RECT 1469.310 265.300 1781.050 265.440 ;
        RECT 1469.310 265.240 1469.630 265.300 ;
        RECT 1780.730 265.240 1781.050 265.300 ;
      LAYER via ;
        RECT 1465.660 945.240 1465.920 945.500 ;
        RECT 1469.340 945.240 1469.600 945.500 ;
        RECT 1469.340 265.240 1469.600 265.500 ;
        RECT 1780.760 265.240 1781.020 265.500 ;
      LAYER met2 ;
        RECT 1465.550 960.500 1465.830 964.000 ;
        RECT 1465.550 960.000 1465.860 960.500 ;
        RECT 1465.720 945.530 1465.860 960.000 ;
        RECT 1465.660 945.210 1465.920 945.530 ;
        RECT 1469.340 945.210 1469.600 945.530 ;
        RECT 1469.400 265.530 1469.540 945.210 ;
        RECT 1469.340 265.210 1469.600 265.530 ;
        RECT 1780.760 265.210 1781.020 265.530 ;
        RECT 1780.820 2.400 1780.960 265.210 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1478.050 945.440 1478.370 945.500 ;
        RECT 1483.110 945.440 1483.430 945.500 ;
        RECT 1478.050 945.300 1483.430 945.440 ;
        RECT 1478.050 945.240 1478.370 945.300 ;
        RECT 1483.110 945.240 1483.430 945.300 ;
        RECT 1483.110 183.160 1483.430 183.220 ;
        RECT 1794.070 183.160 1794.390 183.220 ;
        RECT 1483.110 183.020 1794.390 183.160 ;
        RECT 1483.110 182.960 1483.430 183.020 ;
        RECT 1794.070 182.960 1794.390 183.020 ;
      LAYER via ;
        RECT 1478.080 945.240 1478.340 945.500 ;
        RECT 1483.140 945.240 1483.400 945.500 ;
        RECT 1483.140 182.960 1483.400 183.220 ;
        RECT 1794.100 182.960 1794.360 183.220 ;
      LAYER met2 ;
        RECT 1477.970 960.500 1478.250 964.000 ;
        RECT 1477.970 960.000 1478.280 960.500 ;
        RECT 1478.140 945.530 1478.280 960.000 ;
        RECT 1478.080 945.210 1478.340 945.530 ;
        RECT 1483.140 945.210 1483.400 945.530 ;
        RECT 1483.200 183.250 1483.340 945.210 ;
        RECT 1483.140 182.930 1483.400 183.250 ;
        RECT 1794.100 182.930 1794.360 183.250 ;
        RECT 1794.160 16.730 1794.300 182.930 ;
        RECT 1794.160 16.590 1798.900 16.730 ;
        RECT 1798.760 2.400 1798.900 16.590 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1490.470 945.440 1490.790 945.500 ;
        RECT 1496.910 945.440 1497.230 945.500 ;
        RECT 1490.470 945.300 1497.230 945.440 ;
        RECT 1490.470 945.240 1490.790 945.300 ;
        RECT 1496.910 945.240 1497.230 945.300 ;
        RECT 1496.910 272.580 1497.230 272.640 ;
        RECT 1814.770 272.580 1815.090 272.640 ;
        RECT 1496.910 272.440 1815.090 272.580 ;
        RECT 1496.910 272.380 1497.230 272.440 ;
        RECT 1814.770 272.380 1815.090 272.440 ;
      LAYER via ;
        RECT 1490.500 945.240 1490.760 945.500 ;
        RECT 1496.940 945.240 1497.200 945.500 ;
        RECT 1496.940 272.380 1497.200 272.640 ;
        RECT 1814.800 272.380 1815.060 272.640 ;
      LAYER met2 ;
        RECT 1490.390 960.500 1490.670 964.000 ;
        RECT 1490.390 960.000 1490.700 960.500 ;
        RECT 1490.560 945.530 1490.700 960.000 ;
        RECT 1490.500 945.210 1490.760 945.530 ;
        RECT 1496.940 945.210 1497.200 945.530 ;
        RECT 1497.000 272.670 1497.140 945.210 ;
        RECT 1496.940 272.350 1497.200 272.670 ;
        RECT 1814.800 272.350 1815.060 272.670 ;
        RECT 1814.860 16.730 1815.000 272.350 ;
        RECT 1814.860 16.590 1816.840 16.730 ;
        RECT 1816.700 2.400 1816.840 16.590 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1503.350 279.380 1503.670 279.440 ;
        RECT 1828.570 279.380 1828.890 279.440 ;
        RECT 1503.350 279.240 1828.890 279.380 ;
        RECT 1503.350 279.180 1503.670 279.240 ;
        RECT 1828.570 279.180 1828.890 279.240 ;
        RECT 1828.570 17.920 1828.890 17.980 ;
        RECT 1834.550 17.920 1834.870 17.980 ;
        RECT 1828.570 17.780 1834.870 17.920 ;
        RECT 1828.570 17.720 1828.890 17.780 ;
        RECT 1834.550 17.720 1834.870 17.780 ;
      LAYER via ;
        RECT 1503.380 279.180 1503.640 279.440 ;
        RECT 1828.600 279.180 1828.860 279.440 ;
        RECT 1828.600 17.720 1828.860 17.980 ;
        RECT 1834.580 17.720 1834.840 17.980 ;
      LAYER met2 ;
        RECT 1502.810 960.570 1503.090 964.000 ;
        RECT 1502.810 960.430 1503.580 960.570 ;
        RECT 1502.810 960.000 1503.090 960.430 ;
        RECT 1503.440 279.470 1503.580 960.430 ;
        RECT 1503.380 279.150 1503.640 279.470 ;
        RECT 1828.600 279.150 1828.860 279.470 ;
        RECT 1828.660 18.010 1828.800 279.150 ;
        RECT 1828.600 17.690 1828.860 18.010 ;
        RECT 1834.580 17.690 1834.840 18.010 ;
        RECT 1834.640 2.400 1834.780 17.690 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1517.150 286.180 1517.470 286.240 ;
        RECT 1849.270 286.180 1849.590 286.240 ;
        RECT 1517.150 286.040 1849.590 286.180 ;
        RECT 1517.150 285.980 1517.470 286.040 ;
        RECT 1849.270 285.980 1849.590 286.040 ;
        RECT 1849.270 2.960 1849.590 3.020 ;
        RECT 1852.030 2.960 1852.350 3.020 ;
        RECT 1849.270 2.820 1852.350 2.960 ;
        RECT 1849.270 2.760 1849.590 2.820 ;
        RECT 1852.030 2.760 1852.350 2.820 ;
      LAYER via ;
        RECT 1517.180 285.980 1517.440 286.240 ;
        RECT 1849.300 285.980 1849.560 286.240 ;
        RECT 1849.300 2.760 1849.560 3.020 ;
        RECT 1852.060 2.760 1852.320 3.020 ;
      LAYER met2 ;
        RECT 1515.230 960.570 1515.510 964.000 ;
        RECT 1515.230 960.430 1517.380 960.570 ;
        RECT 1515.230 960.000 1515.510 960.430 ;
        RECT 1517.240 286.270 1517.380 960.430 ;
        RECT 1517.180 285.950 1517.440 286.270 ;
        RECT 1849.300 285.950 1849.560 286.270 ;
        RECT 1849.360 3.050 1849.500 285.950 ;
        RECT 1849.300 2.730 1849.560 3.050 ;
        RECT 1852.060 2.730 1852.320 3.050 ;
        RECT 1852.120 2.400 1852.260 2.730 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 293.320 1531.730 293.380 ;
        RECT 1870.430 293.320 1870.750 293.380 ;
        RECT 1531.410 293.180 1870.750 293.320 ;
        RECT 1531.410 293.120 1531.730 293.180 ;
        RECT 1870.430 293.120 1870.750 293.180 ;
      LAYER via ;
        RECT 1531.440 293.120 1531.700 293.380 ;
        RECT 1870.460 293.120 1870.720 293.380 ;
      LAYER met2 ;
        RECT 1527.650 960.570 1527.930 964.000 ;
        RECT 1527.650 960.430 1531.640 960.570 ;
        RECT 1527.650 960.000 1527.930 960.430 ;
        RECT 1531.500 293.410 1531.640 960.430 ;
        RECT 1531.440 293.090 1531.700 293.410 ;
        RECT 1870.460 293.090 1870.720 293.410 ;
        RECT 1870.520 17.410 1870.660 293.090 ;
        RECT 1870.060 17.270 1870.660 17.410 ;
        RECT 1870.060 2.400 1870.200 17.270 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.410 960.570 748.690 964.000 ;
        RECT 745.360 960.430 748.690 960.570 ;
        RECT 745.360 16.730 745.500 960.430 ;
        RECT 748.410 960.000 748.690 960.430 ;
        RECT 745.360 16.590 746.420 16.730 ;
        RECT 746.280 2.400 746.420 16.590 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1540.150 945.440 1540.470 945.500 ;
        RECT 1544.750 945.440 1545.070 945.500 ;
        RECT 1540.150 945.300 1545.070 945.440 ;
        RECT 1540.150 945.240 1540.470 945.300 ;
        RECT 1544.750 945.240 1545.070 945.300 ;
        RECT 1544.750 300.120 1545.070 300.180 ;
        RECT 1883.770 300.120 1884.090 300.180 ;
        RECT 1544.750 299.980 1884.090 300.120 ;
        RECT 1544.750 299.920 1545.070 299.980 ;
        RECT 1883.770 299.920 1884.090 299.980 ;
        RECT 1883.770 2.960 1884.090 3.020 ;
        RECT 1887.910 2.960 1888.230 3.020 ;
        RECT 1883.770 2.820 1888.230 2.960 ;
        RECT 1883.770 2.760 1884.090 2.820 ;
        RECT 1887.910 2.760 1888.230 2.820 ;
      LAYER via ;
        RECT 1540.180 945.240 1540.440 945.500 ;
        RECT 1544.780 945.240 1545.040 945.500 ;
        RECT 1544.780 299.920 1545.040 300.180 ;
        RECT 1883.800 299.920 1884.060 300.180 ;
        RECT 1883.800 2.760 1884.060 3.020 ;
        RECT 1887.940 2.760 1888.200 3.020 ;
      LAYER met2 ;
        RECT 1540.070 960.500 1540.350 964.000 ;
        RECT 1540.070 960.000 1540.380 960.500 ;
        RECT 1540.240 945.530 1540.380 960.000 ;
        RECT 1540.180 945.210 1540.440 945.530 ;
        RECT 1544.780 945.210 1545.040 945.530 ;
        RECT 1544.840 300.210 1544.980 945.210 ;
        RECT 1544.780 299.890 1545.040 300.210 ;
        RECT 1883.800 299.890 1884.060 300.210 ;
        RECT 1883.860 3.050 1884.000 299.890 ;
        RECT 1883.800 2.730 1884.060 3.050 ;
        RECT 1887.940 2.730 1888.200 3.050 ;
        RECT 1888.000 2.400 1888.140 2.730 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.570 949.520 1552.890 949.580 ;
        RECT 1576.490 949.520 1576.810 949.580 ;
        RECT 1552.570 949.380 1576.810 949.520 ;
        RECT 1552.570 949.320 1552.890 949.380 ;
        RECT 1576.490 949.320 1576.810 949.380 ;
        RECT 1576.490 306.920 1576.810 306.980 ;
        RECT 1904.470 306.920 1904.790 306.980 ;
        RECT 1576.490 306.780 1904.790 306.920 ;
        RECT 1576.490 306.720 1576.810 306.780 ;
        RECT 1904.470 306.720 1904.790 306.780 ;
      LAYER via ;
        RECT 1552.600 949.320 1552.860 949.580 ;
        RECT 1576.520 949.320 1576.780 949.580 ;
        RECT 1576.520 306.720 1576.780 306.980 ;
        RECT 1904.500 306.720 1904.760 306.980 ;
      LAYER met2 ;
        RECT 1552.490 960.500 1552.770 964.000 ;
        RECT 1552.490 960.000 1552.800 960.500 ;
        RECT 1552.660 949.610 1552.800 960.000 ;
        RECT 1552.600 949.290 1552.860 949.610 ;
        RECT 1576.520 949.290 1576.780 949.610 ;
        RECT 1576.580 307.010 1576.720 949.290 ;
        RECT 1576.520 306.690 1576.780 307.010 ;
        RECT 1904.500 306.690 1904.760 307.010 ;
        RECT 1904.560 3.130 1904.700 306.690 ;
        RECT 1904.560 2.990 1906.080 3.130 ;
        RECT 1905.940 2.400 1906.080 2.990 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1565.450 314.060 1565.770 314.120 ;
        RECT 1918.270 314.060 1918.590 314.120 ;
        RECT 1565.450 313.920 1918.590 314.060 ;
        RECT 1565.450 313.860 1565.770 313.920 ;
        RECT 1918.270 313.860 1918.590 313.920 ;
      LAYER via ;
        RECT 1565.480 313.860 1565.740 314.120 ;
        RECT 1918.300 313.860 1918.560 314.120 ;
      LAYER met2 ;
        RECT 1564.910 960.570 1565.190 964.000 ;
        RECT 1564.910 960.430 1565.680 960.570 ;
        RECT 1564.910 960.000 1565.190 960.430 ;
        RECT 1565.540 314.150 1565.680 960.430 ;
        RECT 1565.480 313.830 1565.740 314.150 ;
        RECT 1918.300 313.830 1918.560 314.150 ;
        RECT 1918.360 17.410 1918.500 313.830 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1579.710 210.360 1580.030 210.420 ;
        RECT 1938.970 210.360 1939.290 210.420 ;
        RECT 1579.710 210.220 1939.290 210.360 ;
        RECT 1579.710 210.160 1580.030 210.220 ;
        RECT 1938.970 210.160 1939.290 210.220 ;
      LAYER via ;
        RECT 1579.740 210.160 1580.000 210.420 ;
        RECT 1939.000 210.160 1939.260 210.420 ;
      LAYER met2 ;
        RECT 1576.870 960.570 1577.150 964.000 ;
        RECT 1576.870 960.430 1579.940 960.570 ;
        RECT 1576.870 960.000 1577.150 960.430 ;
        RECT 1579.800 210.450 1579.940 960.430 ;
        RECT 1579.740 210.130 1580.000 210.450 ;
        RECT 1939.000 210.130 1939.260 210.450 ;
        RECT 1939.060 17.410 1939.200 210.130 ;
        RECT 1939.060 17.270 1941.500 17.410 ;
        RECT 1941.360 2.400 1941.500 17.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1593.050 893.420 1593.370 893.480 ;
        RECT 1952.770 893.420 1953.090 893.480 ;
        RECT 1593.050 893.280 1953.090 893.420 ;
        RECT 1593.050 893.220 1593.370 893.280 ;
        RECT 1952.770 893.220 1953.090 893.280 ;
        RECT 1952.770 16.900 1953.090 16.960 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 1952.770 16.760 1959.530 16.900 ;
        RECT 1952.770 16.700 1953.090 16.760 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
      LAYER via ;
        RECT 1593.080 893.220 1593.340 893.480 ;
        RECT 1952.800 893.220 1953.060 893.480 ;
        RECT 1952.800 16.700 1953.060 16.960 ;
        RECT 1959.240 16.700 1959.500 16.960 ;
      LAYER met2 ;
        RECT 1589.290 960.570 1589.570 964.000 ;
        RECT 1589.290 960.430 1593.280 960.570 ;
        RECT 1589.290 960.000 1589.570 960.430 ;
        RECT 1593.140 893.510 1593.280 960.430 ;
        RECT 1593.080 893.190 1593.340 893.510 ;
        RECT 1952.800 893.190 1953.060 893.510 ;
        RECT 1952.860 16.990 1953.000 893.190 ;
        RECT 1952.800 16.670 1953.060 16.990 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 1959.300 2.400 1959.440 16.670 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1601.790 946.460 1602.110 946.520 ;
        RECT 1607.310 946.460 1607.630 946.520 ;
        RECT 1601.790 946.320 1607.630 946.460 ;
        RECT 1601.790 946.260 1602.110 946.320 ;
        RECT 1607.310 946.260 1607.630 946.320 ;
        RECT 1607.310 320.860 1607.630 320.920 ;
        RECT 1973.470 320.860 1973.790 320.920 ;
        RECT 1607.310 320.720 1973.790 320.860 ;
        RECT 1607.310 320.660 1607.630 320.720 ;
        RECT 1973.470 320.660 1973.790 320.720 ;
      LAYER via ;
        RECT 1601.820 946.260 1602.080 946.520 ;
        RECT 1607.340 946.260 1607.600 946.520 ;
        RECT 1607.340 320.660 1607.600 320.920 ;
        RECT 1973.500 320.660 1973.760 320.920 ;
      LAYER met2 ;
        RECT 1601.710 960.500 1601.990 964.000 ;
        RECT 1601.710 960.000 1602.020 960.500 ;
        RECT 1601.880 946.550 1602.020 960.000 ;
        RECT 1601.820 946.230 1602.080 946.550 ;
        RECT 1607.340 946.230 1607.600 946.550 ;
        RECT 1607.400 320.950 1607.540 946.230 ;
        RECT 1607.340 320.630 1607.600 320.950 ;
        RECT 1973.500 320.630 1973.760 320.950 ;
        RECT 1973.560 17.410 1973.700 320.630 ;
        RECT 1973.560 17.270 1977.380 17.410 ;
        RECT 1977.240 2.400 1977.380 17.270 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1613.750 327.660 1614.070 327.720 ;
        RECT 1994.170 327.660 1994.490 327.720 ;
        RECT 1613.750 327.520 1994.490 327.660 ;
        RECT 1613.750 327.460 1614.070 327.520 ;
        RECT 1994.170 327.460 1994.490 327.520 ;
      LAYER via ;
        RECT 1613.780 327.460 1614.040 327.720 ;
        RECT 1994.200 327.460 1994.460 327.720 ;
      LAYER met2 ;
        RECT 1614.130 960.570 1614.410 964.000 ;
        RECT 1613.840 960.430 1614.410 960.570 ;
        RECT 1613.840 327.750 1613.980 960.430 ;
        RECT 1614.130 960.000 1614.410 960.430 ;
        RECT 1613.780 327.430 1614.040 327.750 ;
        RECT 1994.200 327.430 1994.460 327.750 ;
        RECT 1994.260 17.410 1994.400 327.430 ;
        RECT 1994.260 17.270 1995.320 17.410 ;
        RECT 1995.180 2.400 1995.320 17.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.010 224.300 1628.330 224.360 ;
        RECT 2007.970 224.300 2008.290 224.360 ;
        RECT 1628.010 224.160 2008.290 224.300 ;
        RECT 1628.010 224.100 1628.330 224.160 ;
        RECT 2007.970 224.100 2008.290 224.160 ;
      LAYER via ;
        RECT 1628.040 224.100 1628.300 224.360 ;
        RECT 2008.000 224.100 2008.260 224.360 ;
      LAYER met2 ;
        RECT 1626.550 960.570 1626.830 964.000 ;
        RECT 1626.550 960.430 1628.240 960.570 ;
        RECT 1626.550 960.000 1626.830 960.430 ;
        RECT 1628.100 224.390 1628.240 960.430 ;
        RECT 1628.040 224.070 1628.300 224.390 ;
        RECT 2008.000 224.070 2008.260 224.390 ;
        RECT 2008.060 17.410 2008.200 224.070 ;
        RECT 2008.060 17.270 2012.800 17.410 ;
        RECT 2012.660 2.400 2012.800 17.270 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.810 451.760 1642.130 451.820 ;
        RECT 2028.670 451.760 2028.990 451.820 ;
        RECT 1641.810 451.620 2028.990 451.760 ;
        RECT 1641.810 451.560 1642.130 451.620 ;
        RECT 2028.670 451.560 2028.990 451.620 ;
      LAYER via ;
        RECT 1641.840 451.560 1642.100 451.820 ;
        RECT 2028.700 451.560 2028.960 451.820 ;
      LAYER met2 ;
        RECT 1638.970 960.570 1639.250 964.000 ;
        RECT 1638.970 960.430 1642.040 960.570 ;
        RECT 1638.970 960.000 1639.250 960.430 ;
        RECT 1641.900 451.850 1642.040 960.430 ;
        RECT 1641.840 451.530 1642.100 451.850 ;
        RECT 2028.700 451.530 2028.960 451.850 ;
        RECT 2028.760 17.410 2028.900 451.530 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1651.470 947.480 1651.790 947.540 ;
        RECT 1655.610 947.480 1655.930 947.540 ;
        RECT 1651.470 947.340 1655.930 947.480 ;
        RECT 1651.470 947.280 1651.790 947.340 ;
        RECT 1655.610 947.280 1655.930 947.340 ;
        RECT 1655.610 238.240 1655.930 238.300 ;
        RECT 2042.930 238.240 2043.250 238.300 ;
        RECT 1655.610 238.100 2043.250 238.240 ;
        RECT 1655.610 238.040 1655.930 238.100 ;
        RECT 2042.930 238.040 2043.250 238.100 ;
      LAYER via ;
        RECT 1651.500 947.280 1651.760 947.540 ;
        RECT 1655.640 947.280 1655.900 947.540 ;
        RECT 1655.640 238.040 1655.900 238.300 ;
        RECT 2042.960 238.040 2043.220 238.300 ;
      LAYER met2 ;
        RECT 1651.390 960.500 1651.670 964.000 ;
        RECT 1651.390 960.000 1651.700 960.500 ;
        RECT 1651.560 947.570 1651.700 960.000 ;
        RECT 1651.500 947.250 1651.760 947.570 ;
        RECT 1655.640 947.250 1655.900 947.570 ;
        RECT 1655.700 238.330 1655.840 947.250 ;
        RECT 1655.640 238.010 1655.900 238.330 ;
        RECT 2042.960 238.010 2043.220 238.330 ;
        RECT 2043.020 17.410 2043.160 238.010 ;
        RECT 2043.020 17.270 2048.680 17.410 ;
        RECT 2048.540 2.400 2048.680 17.270 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 759.070 17.580 759.390 17.640 ;
        RECT 763.670 17.580 763.990 17.640 ;
        RECT 759.070 17.440 763.990 17.580 ;
        RECT 759.070 17.380 759.390 17.440 ;
        RECT 763.670 17.380 763.990 17.440 ;
      LAYER via ;
        RECT 759.100 17.380 759.360 17.640 ;
        RECT 763.700 17.380 763.960 17.640 ;
      LAYER met2 ;
        RECT 760.830 960.570 761.110 964.000 ;
        RECT 759.160 960.430 761.110 960.570 ;
        RECT 759.160 17.670 759.300 960.430 ;
        RECT 760.830 960.000 761.110 960.430 ;
        RECT 759.100 17.350 759.360 17.670 ;
        RECT 763.700 17.350 763.960 17.670 ;
        RECT 763.760 2.400 763.900 17.350 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1663.890 951.220 1664.210 951.280 ;
        RECT 1669.410 951.220 1669.730 951.280 ;
        RECT 1663.890 951.080 1669.730 951.220 ;
        RECT 1663.890 951.020 1664.210 951.080 ;
        RECT 1669.410 951.020 1669.730 951.080 ;
        RECT 1669.410 334.460 1669.730 334.520 ;
        RECT 2063.170 334.460 2063.490 334.520 ;
        RECT 1669.410 334.320 2063.490 334.460 ;
        RECT 1669.410 334.260 1669.730 334.320 ;
        RECT 2063.170 334.260 2063.490 334.320 ;
      LAYER via ;
        RECT 1663.920 951.020 1664.180 951.280 ;
        RECT 1669.440 951.020 1669.700 951.280 ;
        RECT 1669.440 334.260 1669.700 334.520 ;
        RECT 2063.200 334.260 2063.460 334.520 ;
      LAYER met2 ;
        RECT 1663.810 960.500 1664.090 964.000 ;
        RECT 1663.810 960.000 1664.120 960.500 ;
        RECT 1663.980 951.310 1664.120 960.000 ;
        RECT 1663.920 950.990 1664.180 951.310 ;
        RECT 1669.440 950.990 1669.700 951.310 ;
        RECT 1669.500 334.550 1669.640 950.990 ;
        RECT 1669.440 334.230 1669.700 334.550 ;
        RECT 2063.200 334.230 2063.460 334.550 ;
        RECT 2063.260 17.410 2063.400 334.230 ;
        RECT 2063.260 17.270 2066.620 17.410 ;
        RECT 2066.480 2.400 2066.620 17.270 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 341.600 1676.630 341.660 ;
        RECT 2084.330 341.600 2084.650 341.660 ;
        RECT 1676.310 341.460 2084.650 341.600 ;
        RECT 1676.310 341.400 1676.630 341.460 ;
        RECT 2084.330 341.400 2084.650 341.460 ;
      LAYER via ;
        RECT 1676.340 341.400 1676.600 341.660 ;
        RECT 2084.360 341.400 2084.620 341.660 ;
      LAYER met2 ;
        RECT 1676.230 960.500 1676.510 964.000 ;
        RECT 1676.230 960.000 1676.540 960.500 ;
        RECT 1676.400 341.690 1676.540 960.000 ;
        RECT 1676.340 341.370 1676.600 341.690 ;
        RECT 2084.360 341.370 2084.620 341.690 ;
        RECT 2084.420 2.400 2084.560 341.370 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1689.650 348.400 1689.970 348.460 ;
        RECT 2097.670 348.400 2097.990 348.460 ;
        RECT 1689.650 348.260 2097.990 348.400 ;
        RECT 1689.650 348.200 1689.970 348.260 ;
        RECT 2097.670 348.200 2097.990 348.260 ;
      LAYER via ;
        RECT 1689.680 348.200 1689.940 348.460 ;
        RECT 2097.700 348.200 2097.960 348.460 ;
      LAYER met2 ;
        RECT 1688.190 960.570 1688.470 964.000 ;
        RECT 1688.190 960.430 1689.880 960.570 ;
        RECT 1688.190 960.000 1688.470 960.430 ;
        RECT 1689.740 348.490 1689.880 960.430 ;
        RECT 1689.680 348.170 1689.940 348.490 ;
        RECT 2097.700 348.170 2097.960 348.490 ;
        RECT 2097.760 17.410 2097.900 348.170 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.910 355.200 1704.230 355.260 ;
        RECT 2118.370 355.200 2118.690 355.260 ;
        RECT 1703.910 355.060 2118.690 355.200 ;
        RECT 1703.910 355.000 1704.230 355.060 ;
        RECT 2118.370 355.000 2118.690 355.060 ;
      LAYER via ;
        RECT 1703.940 355.000 1704.200 355.260 ;
        RECT 2118.400 355.000 2118.660 355.260 ;
      LAYER met2 ;
        RECT 1700.610 960.570 1700.890 964.000 ;
        RECT 1700.610 960.430 1704.140 960.570 ;
        RECT 1700.610 960.000 1700.890 960.430 ;
        RECT 1704.000 355.290 1704.140 960.430 ;
        RECT 1703.940 354.970 1704.200 355.290 ;
        RECT 2118.400 354.970 2118.660 355.290 ;
        RECT 2118.460 17.410 2118.600 354.970 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1713.110 945.440 1713.430 945.500 ;
        RECT 1721.390 945.440 1721.710 945.500 ;
        RECT 1713.110 945.300 1721.710 945.440 ;
        RECT 1713.110 945.240 1713.430 945.300 ;
        RECT 1721.390 945.240 1721.710 945.300 ;
        RECT 1721.390 362.340 1721.710 362.400 ;
        RECT 2132.170 362.340 2132.490 362.400 ;
        RECT 1721.390 362.200 2132.490 362.340 ;
        RECT 1721.390 362.140 1721.710 362.200 ;
        RECT 2132.170 362.140 2132.490 362.200 ;
      LAYER via ;
        RECT 1713.140 945.240 1713.400 945.500 ;
        RECT 1721.420 945.240 1721.680 945.500 ;
        RECT 1721.420 362.140 1721.680 362.400 ;
        RECT 2132.200 362.140 2132.460 362.400 ;
      LAYER met2 ;
        RECT 1713.030 960.500 1713.310 964.000 ;
        RECT 1713.030 960.000 1713.340 960.500 ;
        RECT 1713.200 945.530 1713.340 960.000 ;
        RECT 1713.140 945.210 1713.400 945.530 ;
        RECT 1721.420 945.210 1721.680 945.530 ;
        RECT 1721.480 362.430 1721.620 945.210 ;
        RECT 1721.420 362.110 1721.680 362.430 ;
        RECT 2132.200 362.110 2132.460 362.430 ;
        RECT 2132.260 17.410 2132.400 362.110 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1725.530 950.540 1725.850 950.600 ;
        RECT 1731.050 950.540 1731.370 950.600 ;
        RECT 1725.530 950.400 1731.370 950.540 ;
        RECT 1725.530 950.340 1725.850 950.400 ;
        RECT 1731.050 950.340 1731.370 950.400 ;
        RECT 1731.050 369.140 1731.370 369.200 ;
        RECT 2152.870 369.140 2153.190 369.200 ;
        RECT 1731.050 369.000 2153.190 369.140 ;
        RECT 1731.050 368.940 1731.370 369.000 ;
        RECT 2152.870 368.940 2153.190 369.000 ;
      LAYER via ;
        RECT 1725.560 950.340 1725.820 950.600 ;
        RECT 1731.080 950.340 1731.340 950.600 ;
        RECT 1731.080 368.940 1731.340 369.200 ;
        RECT 2152.900 368.940 2153.160 369.200 ;
      LAYER met2 ;
        RECT 1725.450 960.500 1725.730 964.000 ;
        RECT 1725.450 960.000 1725.760 960.500 ;
        RECT 1725.620 950.630 1725.760 960.000 ;
        RECT 1725.560 950.310 1725.820 950.630 ;
        RECT 1731.080 950.310 1731.340 950.630 ;
        RECT 1731.140 369.230 1731.280 950.310 ;
        RECT 1731.080 368.910 1731.340 369.230 ;
        RECT 2152.900 368.910 2153.160 369.230 ;
        RECT 2152.960 17.410 2153.100 368.910 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.410 375.940 1738.730 376.000 ;
        RECT 2166.670 375.940 2166.990 376.000 ;
        RECT 1738.410 375.800 2166.990 375.940 ;
        RECT 1738.410 375.740 1738.730 375.800 ;
        RECT 2166.670 375.740 2166.990 375.800 ;
        RECT 2166.670 16.900 2166.990 16.960 ;
        RECT 2173.110 16.900 2173.430 16.960 ;
        RECT 2166.670 16.760 2173.430 16.900 ;
        RECT 2166.670 16.700 2166.990 16.760 ;
        RECT 2173.110 16.700 2173.430 16.760 ;
      LAYER via ;
        RECT 1738.440 375.740 1738.700 376.000 ;
        RECT 2166.700 375.740 2166.960 376.000 ;
        RECT 2166.700 16.700 2166.960 16.960 ;
        RECT 2173.140 16.700 2173.400 16.960 ;
      LAYER met2 ;
        RECT 1737.870 960.570 1738.150 964.000 ;
        RECT 1737.870 960.430 1738.640 960.570 ;
        RECT 1737.870 960.000 1738.150 960.430 ;
        RECT 1738.500 376.030 1738.640 960.430 ;
        RECT 1738.440 375.710 1738.700 376.030 ;
        RECT 2166.700 375.710 2166.960 376.030 ;
        RECT 2166.760 16.990 2166.900 375.710 ;
        RECT 2166.700 16.670 2166.960 16.990 ;
        RECT 2173.140 16.670 2173.400 16.990 ;
        RECT 2173.200 2.400 2173.340 16.670 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1752.210 258.640 1752.530 258.700 ;
        RECT 2187.370 258.640 2187.690 258.700 ;
        RECT 1752.210 258.500 2187.690 258.640 ;
        RECT 1752.210 258.440 1752.530 258.500 ;
        RECT 2187.370 258.440 2187.690 258.500 ;
      LAYER via ;
        RECT 1752.240 258.440 1752.500 258.700 ;
        RECT 2187.400 258.440 2187.660 258.700 ;
      LAYER met2 ;
        RECT 1750.290 960.570 1750.570 964.000 ;
        RECT 1750.290 960.430 1752.440 960.570 ;
        RECT 1750.290 960.000 1750.570 960.430 ;
        RECT 1752.300 258.730 1752.440 960.430 ;
        RECT 1752.240 258.410 1752.500 258.730 ;
        RECT 2187.400 258.410 2187.660 258.730 ;
        RECT 2187.460 17.410 2187.600 258.410 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 382.740 1766.330 382.800 ;
        RECT 2208.070 382.740 2208.390 382.800 ;
        RECT 1766.010 382.600 2208.390 382.740 ;
        RECT 1766.010 382.540 1766.330 382.600 ;
        RECT 2208.070 382.540 2208.390 382.600 ;
      LAYER via ;
        RECT 1766.040 382.540 1766.300 382.800 ;
        RECT 2208.100 382.540 2208.360 382.800 ;
      LAYER met2 ;
        RECT 1762.710 960.570 1762.990 964.000 ;
        RECT 1762.710 960.430 1766.240 960.570 ;
        RECT 1762.710 960.000 1762.990 960.430 ;
        RECT 1766.100 382.830 1766.240 960.430 ;
        RECT 1766.040 382.510 1766.300 382.830 ;
        RECT 2208.100 382.510 2208.360 382.830 ;
        RECT 2208.160 16.730 2208.300 382.510 ;
        RECT 2208.160 16.590 2209.220 16.730 ;
        RECT 2209.080 2.400 2209.220 16.590 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1775.210 945.440 1775.530 945.500 ;
        RECT 1779.350 945.440 1779.670 945.500 ;
        RECT 1775.210 945.300 1779.670 945.440 ;
        RECT 1775.210 945.240 1775.530 945.300 ;
        RECT 1779.350 945.240 1779.670 945.300 ;
        RECT 1779.350 396.680 1779.670 396.740 ;
        RECT 2221.870 396.680 2222.190 396.740 ;
        RECT 1779.350 396.540 2222.190 396.680 ;
        RECT 1779.350 396.480 1779.670 396.540 ;
        RECT 2221.870 396.480 2222.190 396.540 ;
      LAYER via ;
        RECT 1775.240 945.240 1775.500 945.500 ;
        RECT 1779.380 945.240 1779.640 945.500 ;
        RECT 1779.380 396.480 1779.640 396.740 ;
        RECT 2221.900 396.480 2222.160 396.740 ;
      LAYER met2 ;
        RECT 1775.130 960.500 1775.410 964.000 ;
        RECT 1775.130 960.000 1775.440 960.500 ;
        RECT 1775.300 945.530 1775.440 960.000 ;
        RECT 1775.240 945.210 1775.500 945.530 ;
        RECT 1779.380 945.210 1779.640 945.530 ;
        RECT 1779.440 396.770 1779.580 945.210 ;
        RECT 1779.380 396.450 1779.640 396.770 ;
        RECT 2221.900 396.450 2222.160 396.770 ;
        RECT 2221.960 16.730 2222.100 396.450 ;
        RECT 2221.960 16.590 2227.160 16.730 ;
        RECT 2227.020 2.400 2227.160 16.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 773.330 950.540 773.650 950.600 ;
        RECT 778.850 950.540 779.170 950.600 ;
        RECT 773.330 950.400 779.170 950.540 ;
        RECT 773.330 950.340 773.650 950.400 ;
        RECT 778.850 950.340 779.170 950.400 ;
        RECT 778.850 17.580 779.170 17.640 ;
        RECT 781.610 17.580 781.930 17.640 ;
        RECT 778.850 17.440 781.930 17.580 ;
        RECT 778.850 17.380 779.170 17.440 ;
        RECT 781.610 17.380 781.930 17.440 ;
      LAYER via ;
        RECT 773.360 950.340 773.620 950.600 ;
        RECT 778.880 950.340 779.140 950.600 ;
        RECT 778.880 17.380 779.140 17.640 ;
        RECT 781.640 17.380 781.900 17.640 ;
      LAYER met2 ;
        RECT 773.250 960.500 773.530 964.000 ;
        RECT 773.250 960.000 773.560 960.500 ;
        RECT 773.420 950.630 773.560 960.000 ;
        RECT 773.360 950.310 773.620 950.630 ;
        RECT 778.880 950.310 779.140 950.630 ;
        RECT 778.940 17.670 779.080 950.310 ;
        RECT 778.880 17.350 779.140 17.670 ;
        RECT 781.640 17.350 781.900 17.670 ;
        RECT 781.700 2.400 781.840 17.350 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1787.630 949.860 1787.950 949.920 ;
        RECT 1793.150 949.860 1793.470 949.920 ;
        RECT 1787.630 949.720 1793.470 949.860 ;
        RECT 1787.630 949.660 1787.950 949.720 ;
        RECT 1793.150 949.660 1793.470 949.720 ;
        RECT 1793.150 265.440 1793.470 265.500 ;
        RECT 2242.570 265.440 2242.890 265.500 ;
        RECT 1793.150 265.300 2242.890 265.440 ;
        RECT 1793.150 265.240 1793.470 265.300 ;
        RECT 2242.570 265.240 2242.890 265.300 ;
      LAYER via ;
        RECT 1787.660 949.660 1787.920 949.920 ;
        RECT 1793.180 949.660 1793.440 949.920 ;
        RECT 1793.180 265.240 1793.440 265.500 ;
        RECT 2242.600 265.240 2242.860 265.500 ;
      LAYER met2 ;
        RECT 1787.550 960.500 1787.830 964.000 ;
        RECT 1787.550 960.000 1787.860 960.500 ;
        RECT 1787.720 949.950 1787.860 960.000 ;
        RECT 1787.660 949.630 1787.920 949.950 ;
        RECT 1793.180 949.630 1793.440 949.950 ;
        RECT 1793.240 265.530 1793.380 949.630 ;
        RECT 1793.180 265.210 1793.440 265.530 ;
        RECT 2242.600 265.210 2242.860 265.530 ;
        RECT 2242.660 16.730 2242.800 265.210 ;
        RECT 2242.660 16.590 2245.100 16.730 ;
        RECT 2244.960 2.400 2245.100 16.590 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.050 389.880 1800.370 389.940 ;
        RECT 2256.370 389.880 2256.690 389.940 ;
        RECT 1800.050 389.740 2256.690 389.880 ;
        RECT 1800.050 389.680 1800.370 389.740 ;
        RECT 2256.370 389.680 2256.690 389.740 ;
        RECT 2256.370 20.980 2256.690 21.040 ;
        RECT 2262.350 20.980 2262.670 21.040 ;
        RECT 2256.370 20.840 2262.670 20.980 ;
        RECT 2256.370 20.780 2256.690 20.840 ;
        RECT 2262.350 20.780 2262.670 20.840 ;
      LAYER via ;
        RECT 1800.080 389.680 1800.340 389.940 ;
        RECT 2256.400 389.680 2256.660 389.940 ;
        RECT 2256.400 20.780 2256.660 21.040 ;
        RECT 2262.380 20.780 2262.640 21.040 ;
      LAYER met2 ;
        RECT 1799.510 960.570 1799.790 964.000 ;
        RECT 1799.510 960.430 1800.280 960.570 ;
        RECT 1799.510 960.000 1799.790 960.430 ;
        RECT 1800.140 389.970 1800.280 960.430 ;
        RECT 1800.080 389.650 1800.340 389.970 ;
        RECT 2256.400 389.650 2256.660 389.970 ;
        RECT 2256.460 21.070 2256.600 389.650 ;
        RECT 2256.400 20.750 2256.660 21.070 ;
        RECT 2262.380 20.750 2262.640 21.070 ;
        RECT 2262.440 2.400 2262.580 20.750 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1813.850 403.480 1814.170 403.540 ;
        RECT 2277.070 403.480 2277.390 403.540 ;
        RECT 1813.850 403.340 2277.390 403.480 ;
        RECT 1813.850 403.280 1814.170 403.340 ;
        RECT 2277.070 403.280 2277.390 403.340 ;
      LAYER via ;
        RECT 1813.880 403.280 1814.140 403.540 ;
        RECT 2277.100 403.280 2277.360 403.540 ;
      LAYER met2 ;
        RECT 1811.930 960.570 1812.210 964.000 ;
        RECT 1811.930 960.430 1814.080 960.570 ;
        RECT 1811.930 960.000 1812.210 960.430 ;
        RECT 1813.940 403.570 1814.080 960.430 ;
        RECT 1813.880 403.250 1814.140 403.570 ;
        RECT 2277.100 403.250 2277.360 403.570 ;
        RECT 2277.160 17.410 2277.300 403.250 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1824.430 945.440 1824.750 945.500 ;
        RECT 1828.110 945.440 1828.430 945.500 ;
        RECT 1824.430 945.300 1828.430 945.440 ;
        RECT 1824.430 945.240 1824.750 945.300 ;
        RECT 1828.110 945.240 1828.430 945.300 ;
        RECT 1828.110 790.060 1828.430 790.120 ;
        RECT 2298.230 790.060 2298.550 790.120 ;
        RECT 1828.110 789.920 2298.550 790.060 ;
        RECT 1828.110 789.860 1828.430 789.920 ;
        RECT 2298.230 789.860 2298.550 789.920 ;
      LAYER via ;
        RECT 1824.460 945.240 1824.720 945.500 ;
        RECT 1828.140 945.240 1828.400 945.500 ;
        RECT 1828.140 789.860 1828.400 790.120 ;
        RECT 2298.260 789.860 2298.520 790.120 ;
      LAYER met2 ;
        RECT 1824.350 960.500 1824.630 964.000 ;
        RECT 1824.350 960.000 1824.660 960.500 ;
        RECT 1824.520 945.530 1824.660 960.000 ;
        RECT 1824.460 945.210 1824.720 945.530 ;
        RECT 1828.140 945.210 1828.400 945.530 ;
        RECT 1828.200 790.150 1828.340 945.210 ;
        RECT 1828.140 789.830 1828.400 790.150 ;
        RECT 2298.260 789.830 2298.520 790.150 ;
        RECT 2298.320 2.400 2298.460 789.830 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1836.850 907.360 1837.170 907.420 ;
        RECT 2311.570 907.360 2311.890 907.420 ;
        RECT 1836.850 907.220 2311.890 907.360 ;
        RECT 1836.850 907.160 1837.170 907.220 ;
        RECT 2311.570 907.160 2311.890 907.220 ;
      LAYER via ;
        RECT 1836.880 907.160 1837.140 907.420 ;
        RECT 2311.600 907.160 2311.860 907.420 ;
      LAYER met2 ;
        RECT 1836.770 960.500 1837.050 964.000 ;
        RECT 1836.770 960.000 1837.080 960.500 ;
        RECT 1836.940 907.450 1837.080 960.000 ;
        RECT 1836.880 907.130 1837.140 907.450 ;
        RECT 2311.600 907.130 2311.860 907.450 ;
        RECT 2311.660 17.410 2311.800 907.130 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1849.270 950.200 1849.590 950.260 ;
        RECT 1855.250 950.200 1855.570 950.260 ;
        RECT 1849.270 950.060 1855.570 950.200 ;
        RECT 1849.270 950.000 1849.590 950.060 ;
        RECT 1855.250 950.000 1855.570 950.060 ;
        RECT 1855.250 700.300 1855.570 700.360 ;
        RECT 2332.270 700.300 2332.590 700.360 ;
        RECT 1855.250 700.160 2332.590 700.300 ;
        RECT 1855.250 700.100 1855.570 700.160 ;
        RECT 2332.270 700.100 2332.590 700.160 ;
      LAYER via ;
        RECT 1849.300 950.000 1849.560 950.260 ;
        RECT 1855.280 950.000 1855.540 950.260 ;
        RECT 1855.280 700.100 1855.540 700.360 ;
        RECT 2332.300 700.100 2332.560 700.360 ;
      LAYER met2 ;
        RECT 1849.190 960.500 1849.470 964.000 ;
        RECT 1849.190 960.000 1849.500 960.500 ;
        RECT 1849.360 950.290 1849.500 960.000 ;
        RECT 1849.300 949.970 1849.560 950.290 ;
        RECT 1855.280 949.970 1855.540 950.290 ;
        RECT 1855.340 700.390 1855.480 949.970 ;
        RECT 1855.280 700.070 1855.540 700.390 ;
        RECT 2332.300 700.070 2332.560 700.390 ;
        RECT 2332.360 17.410 2332.500 700.070 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1862.150 555.460 1862.470 555.520 ;
        RECT 2346.070 555.460 2346.390 555.520 ;
        RECT 1862.150 555.320 2346.390 555.460 ;
        RECT 1862.150 555.260 1862.470 555.320 ;
        RECT 2346.070 555.260 2346.390 555.320 ;
      LAYER via ;
        RECT 1862.180 555.260 1862.440 555.520 ;
        RECT 2346.100 555.260 2346.360 555.520 ;
      LAYER met2 ;
        RECT 1861.610 960.570 1861.890 964.000 ;
        RECT 1861.610 960.430 1862.380 960.570 ;
        RECT 1861.610 960.000 1861.890 960.430 ;
        RECT 1862.240 555.550 1862.380 960.430 ;
        RECT 1862.180 555.230 1862.440 555.550 ;
        RECT 2346.100 555.230 2346.360 555.550 ;
        RECT 2346.160 17.410 2346.300 555.230 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1875.950 438.160 1876.270 438.220 ;
        RECT 2366.770 438.160 2367.090 438.220 ;
        RECT 1875.950 438.020 2367.090 438.160 ;
        RECT 1875.950 437.960 1876.270 438.020 ;
        RECT 2366.770 437.960 2367.090 438.020 ;
      LAYER via ;
        RECT 1875.980 437.960 1876.240 438.220 ;
        RECT 2366.800 437.960 2367.060 438.220 ;
      LAYER met2 ;
        RECT 1874.030 960.570 1874.310 964.000 ;
        RECT 1874.030 960.430 1876.180 960.570 ;
        RECT 1874.030 960.000 1874.310 960.430 ;
        RECT 1876.040 438.250 1876.180 960.430 ;
        RECT 1875.980 437.930 1876.240 438.250 ;
        RECT 2366.800 437.930 2367.060 438.250 ;
        RECT 2366.860 17.410 2367.000 437.930 ;
        RECT 2366.860 17.270 2369.760 17.410 ;
        RECT 2369.620 2.400 2369.760 17.270 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 272.580 1890.530 272.640 ;
        RECT 2387.930 272.580 2388.250 272.640 ;
        RECT 1890.210 272.440 2388.250 272.580 ;
        RECT 1890.210 272.380 1890.530 272.440 ;
        RECT 2387.930 272.380 2388.250 272.440 ;
      LAYER via ;
        RECT 1890.240 272.380 1890.500 272.640 ;
        RECT 2387.960 272.380 2388.220 272.640 ;
      LAYER met2 ;
        RECT 1886.450 960.570 1886.730 964.000 ;
        RECT 1886.450 960.430 1890.440 960.570 ;
        RECT 1886.450 960.000 1886.730 960.430 ;
        RECT 1890.300 272.670 1890.440 960.430 ;
        RECT 1890.240 272.350 1890.500 272.670 ;
        RECT 2387.960 272.350 2388.220 272.670 ;
        RECT 2388.020 17.410 2388.160 272.350 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1898.950 945.440 1899.270 945.500 ;
        RECT 1903.550 945.440 1903.870 945.500 ;
        RECT 1898.950 945.300 1903.870 945.440 ;
        RECT 1898.950 945.240 1899.270 945.300 ;
        RECT 1903.550 945.240 1903.870 945.300 ;
        RECT 1903.550 693.500 1903.870 693.560 ;
        RECT 2401.270 693.500 2401.590 693.560 ;
        RECT 1903.550 693.360 2401.590 693.500 ;
        RECT 1903.550 693.300 1903.870 693.360 ;
        RECT 2401.270 693.300 2401.590 693.360 ;
      LAYER via ;
        RECT 1898.980 945.240 1899.240 945.500 ;
        RECT 1903.580 945.240 1903.840 945.500 ;
        RECT 1903.580 693.300 1903.840 693.560 ;
        RECT 2401.300 693.300 2401.560 693.560 ;
      LAYER met2 ;
        RECT 1898.870 960.500 1899.150 964.000 ;
        RECT 1898.870 960.000 1899.180 960.500 ;
        RECT 1899.040 945.530 1899.180 960.000 ;
        RECT 1898.980 945.210 1899.240 945.530 ;
        RECT 1903.580 945.210 1903.840 945.530 ;
        RECT 1903.640 693.590 1903.780 945.210 ;
        RECT 1903.580 693.270 1903.840 693.590 ;
        RECT 2401.300 693.270 2401.560 693.590 ;
        RECT 2401.360 17.410 2401.500 693.270 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 785.750 15.200 786.070 15.260 ;
        RECT 799.550 15.200 799.870 15.260 ;
        RECT 785.750 15.060 799.870 15.200 ;
        RECT 785.750 15.000 786.070 15.060 ;
        RECT 799.550 15.000 799.870 15.060 ;
      LAYER via ;
        RECT 785.780 15.000 786.040 15.260 ;
        RECT 799.580 15.000 799.840 15.260 ;
      LAYER met2 ;
        RECT 785.210 960.570 785.490 964.000 ;
        RECT 785.210 960.430 785.980 960.570 ;
        RECT 785.210 960.000 785.490 960.430 ;
        RECT 785.840 15.290 785.980 960.430 ;
        RECT 785.780 14.970 786.040 15.290 ;
        RECT 799.580 14.970 799.840 15.290 ;
        RECT 799.640 2.400 799.780 14.970 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 19.960 645.310 20.020 ;
        RECT 676.270 19.960 676.590 20.020 ;
        RECT 644.990 19.820 676.590 19.960 ;
        RECT 644.990 19.760 645.310 19.820 ;
        RECT 676.270 19.760 676.590 19.820 ;
      LAYER via ;
        RECT 645.020 19.760 645.280 20.020 ;
        RECT 676.300 19.760 676.560 20.020 ;
      LAYER met2 ;
        RECT 678.030 960.570 678.310 964.000 ;
        RECT 676.360 960.430 678.310 960.570 ;
        RECT 676.360 20.050 676.500 960.430 ;
        RECT 678.030 960.000 678.310 960.430 ;
        RECT 645.020 19.730 645.280 20.050 ;
        RECT 676.300 19.730 676.560 20.050 ;
        RECT 645.080 2.400 645.220 19.730 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 286.180 1918.130 286.240 ;
        RECT 2429.330 286.180 2429.650 286.240 ;
        RECT 1917.810 286.040 2429.650 286.180 ;
        RECT 1917.810 285.980 1918.130 286.040 ;
        RECT 2429.330 285.980 2429.650 286.040 ;
      LAYER via ;
        RECT 1917.840 285.980 1918.100 286.240 ;
        RECT 2429.360 285.980 2429.620 286.240 ;
      LAYER met2 ;
        RECT 1914.970 960.570 1915.250 964.000 ;
        RECT 1914.970 960.430 1918.040 960.570 ;
        RECT 1914.970 960.000 1915.250 960.430 ;
        RECT 1917.900 286.270 1918.040 960.430 ;
        RECT 1917.840 285.950 1918.100 286.270 ;
        RECT 2429.360 285.950 2429.620 286.270 ;
        RECT 2429.420 17.410 2429.560 285.950 ;
        RECT 2428.960 17.270 2429.560 17.410 ;
        RECT 2428.960 2.400 2429.100 17.270 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1927.470 945.440 1927.790 945.500 ;
        RECT 1931.150 945.440 1931.470 945.500 ;
        RECT 1927.470 945.300 1931.470 945.440 ;
        RECT 1927.470 945.240 1927.790 945.300 ;
        RECT 1931.150 945.240 1931.470 945.300 ;
        RECT 1931.150 686.360 1931.470 686.420 ;
        RECT 2442.670 686.360 2442.990 686.420 ;
        RECT 1931.150 686.220 2442.990 686.360 ;
        RECT 1931.150 686.160 1931.470 686.220 ;
        RECT 2442.670 686.160 2442.990 686.220 ;
      LAYER via ;
        RECT 1927.500 945.240 1927.760 945.500 ;
        RECT 1931.180 945.240 1931.440 945.500 ;
        RECT 1931.180 686.160 1931.440 686.420 ;
        RECT 2442.700 686.160 2442.960 686.420 ;
      LAYER met2 ;
        RECT 1927.390 960.500 1927.670 964.000 ;
        RECT 1927.390 960.000 1927.700 960.500 ;
        RECT 1927.560 945.530 1927.700 960.000 ;
        RECT 1927.500 945.210 1927.760 945.530 ;
        RECT 1931.180 945.210 1931.440 945.530 ;
        RECT 1931.240 686.450 1931.380 945.210 ;
        RECT 1931.180 686.130 1931.440 686.450 ;
        RECT 2442.700 686.130 2442.960 686.450 ;
        RECT 2442.760 17.410 2442.900 686.130 ;
        RECT 2442.760 17.270 2447.040 17.410 ;
        RECT 2446.900 2.400 2447.040 17.270 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1939.890 945.440 1940.210 945.500 ;
        RECT 1944.950 945.440 1945.270 945.500 ;
        RECT 1939.890 945.300 1945.270 945.440 ;
        RECT 1939.890 945.240 1940.210 945.300 ;
        RECT 1944.950 945.240 1945.270 945.300 ;
        RECT 1944.950 279.380 1945.270 279.440 ;
        RECT 2463.370 279.380 2463.690 279.440 ;
        RECT 1944.950 279.240 2463.690 279.380 ;
        RECT 1944.950 279.180 1945.270 279.240 ;
        RECT 2463.370 279.180 2463.690 279.240 ;
      LAYER via ;
        RECT 1939.920 945.240 1940.180 945.500 ;
        RECT 1944.980 945.240 1945.240 945.500 ;
        RECT 1944.980 279.180 1945.240 279.440 ;
        RECT 2463.400 279.180 2463.660 279.440 ;
      LAYER met2 ;
        RECT 1939.810 960.500 1940.090 964.000 ;
        RECT 1939.810 960.000 1940.120 960.500 ;
        RECT 1939.980 945.530 1940.120 960.000 ;
        RECT 1939.920 945.210 1940.180 945.530 ;
        RECT 1944.980 945.210 1945.240 945.530 ;
        RECT 1945.040 279.470 1945.180 945.210 ;
        RECT 1944.980 279.150 1945.240 279.470 ;
        RECT 2463.400 279.150 2463.660 279.470 ;
        RECT 2463.460 17.410 2463.600 279.150 ;
        RECT 2463.460 17.270 2464.980 17.410 ;
        RECT 2464.840 2.400 2464.980 17.270 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1951.850 679.560 1952.170 679.620 ;
        RECT 2477.170 679.560 2477.490 679.620 ;
        RECT 1951.850 679.420 2477.490 679.560 ;
        RECT 1951.850 679.360 1952.170 679.420 ;
        RECT 2477.170 679.360 2477.490 679.420 ;
      LAYER via ;
        RECT 1951.880 679.360 1952.140 679.620 ;
        RECT 2477.200 679.360 2477.460 679.620 ;
      LAYER met2 ;
        RECT 1952.230 960.570 1952.510 964.000 ;
        RECT 1951.940 960.430 1952.510 960.570 ;
        RECT 1951.940 679.650 1952.080 960.430 ;
        RECT 1952.230 960.000 1952.510 960.430 ;
        RECT 1951.880 679.330 1952.140 679.650 ;
        RECT 2477.200 679.330 2477.460 679.650 ;
        RECT 2477.260 17.410 2477.400 679.330 ;
        RECT 2477.260 17.270 2482.920 17.410 ;
        RECT 2482.780 2.400 2482.920 17.270 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 293.320 1966.430 293.380 ;
        RECT 2497.870 293.320 2498.190 293.380 ;
        RECT 1966.110 293.180 2498.190 293.320 ;
        RECT 1966.110 293.120 1966.430 293.180 ;
        RECT 2497.870 293.120 2498.190 293.180 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 1966.140 293.120 1966.400 293.380 ;
        RECT 2497.900 293.120 2498.160 293.380 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 1964.650 960.570 1964.930 964.000 ;
        RECT 1964.650 960.430 1966.340 960.570 ;
        RECT 1964.650 960.000 1964.930 960.430 ;
        RECT 1966.200 293.410 1966.340 960.430 ;
        RECT 1966.140 293.090 1966.400 293.410 ;
        RECT 2497.900 293.090 2498.160 293.410 ;
        RECT 2497.960 3.050 2498.100 293.090 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 410.620 1980.230 410.680 ;
        RECT 2511.670 410.620 2511.990 410.680 ;
        RECT 1979.910 410.480 2511.990 410.620 ;
        RECT 1979.910 410.420 1980.230 410.480 ;
        RECT 2511.670 410.420 2511.990 410.480 ;
        RECT 2511.670 13.840 2511.990 13.900 ;
        RECT 2518.110 13.840 2518.430 13.900 ;
        RECT 2511.670 13.700 2518.430 13.840 ;
        RECT 2511.670 13.640 2511.990 13.700 ;
        RECT 2518.110 13.640 2518.430 13.700 ;
      LAYER via ;
        RECT 1979.940 410.420 1980.200 410.680 ;
        RECT 2511.700 410.420 2511.960 410.680 ;
        RECT 2511.700 13.640 2511.960 13.900 ;
        RECT 2518.140 13.640 2518.400 13.900 ;
      LAYER met2 ;
        RECT 1977.070 960.570 1977.350 964.000 ;
        RECT 1977.070 960.430 1980.140 960.570 ;
        RECT 1977.070 960.000 1977.350 960.430 ;
        RECT 1980.000 410.710 1980.140 960.430 ;
        RECT 1979.940 410.390 1980.200 410.710 ;
        RECT 2511.700 410.390 2511.960 410.710 ;
        RECT 2511.760 13.930 2511.900 410.390 ;
        RECT 2511.700 13.610 2511.960 13.930 ;
        RECT 2518.140 13.610 2518.400 13.930 ;
        RECT 2518.200 2.400 2518.340 13.610 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.250 665.960 1993.570 666.020 ;
        RECT 2532.370 665.960 2532.690 666.020 ;
        RECT 1993.250 665.820 2532.690 665.960 ;
        RECT 1993.250 665.760 1993.570 665.820 ;
        RECT 2532.370 665.760 2532.690 665.820 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 1993.280 665.760 1993.540 666.020 ;
        RECT 2532.400 665.760 2532.660 666.020 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 1989.490 960.570 1989.770 964.000 ;
        RECT 1989.490 960.430 1993.480 960.570 ;
        RECT 1989.490 960.000 1989.770 960.430 ;
        RECT 1993.340 666.050 1993.480 960.430 ;
        RECT 1993.280 665.730 1993.540 666.050 ;
        RECT 2532.400 665.730 2532.660 666.050 ;
        RECT 2532.460 3.050 2532.600 665.730 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2001.990 945.440 2002.310 945.500 ;
        RECT 2007.510 945.440 2007.830 945.500 ;
        RECT 2001.990 945.300 2007.830 945.440 ;
        RECT 2001.990 945.240 2002.310 945.300 ;
        RECT 2007.510 945.240 2007.830 945.300 ;
        RECT 2007.510 658.820 2007.830 658.880 ;
        RECT 2553.070 658.820 2553.390 658.880 ;
        RECT 2007.510 658.680 2553.390 658.820 ;
        RECT 2007.510 658.620 2007.830 658.680 ;
        RECT 2553.070 658.620 2553.390 658.680 ;
      LAYER via ;
        RECT 2002.020 945.240 2002.280 945.500 ;
        RECT 2007.540 945.240 2007.800 945.500 ;
        RECT 2007.540 658.620 2007.800 658.880 ;
        RECT 2553.100 658.620 2553.360 658.880 ;
      LAYER met2 ;
        RECT 2001.910 960.500 2002.190 964.000 ;
        RECT 2001.910 960.000 2002.220 960.500 ;
        RECT 2002.080 945.530 2002.220 960.000 ;
        RECT 2002.020 945.210 2002.280 945.530 ;
        RECT 2007.540 945.210 2007.800 945.530 ;
        RECT 2007.600 658.910 2007.740 945.210 ;
        RECT 2007.540 658.590 2007.800 658.910 ;
        RECT 2553.100 658.590 2553.360 658.910 ;
        RECT 2553.160 17.410 2553.300 658.590 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2013.950 652.020 2014.270 652.080 ;
        RECT 2566.870 652.020 2567.190 652.080 ;
        RECT 2013.950 651.880 2567.190 652.020 ;
        RECT 2013.950 651.820 2014.270 651.880 ;
        RECT 2566.870 651.820 2567.190 651.880 ;
      LAYER via ;
        RECT 2013.980 651.820 2014.240 652.080 ;
        RECT 2566.900 651.820 2567.160 652.080 ;
      LAYER met2 ;
        RECT 2014.330 960.570 2014.610 964.000 ;
        RECT 2014.040 960.430 2014.610 960.570 ;
        RECT 2014.040 652.110 2014.180 960.430 ;
        RECT 2014.330 960.000 2014.610 960.430 ;
        RECT 2013.980 651.790 2014.240 652.110 ;
        RECT 2566.900 651.790 2567.160 652.110 ;
        RECT 2566.960 17.410 2567.100 651.790 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.400 2572.160 17.270 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.210 314.060 2028.530 314.120 ;
        RECT 2587.570 314.060 2587.890 314.120 ;
        RECT 2028.210 313.920 2587.890 314.060 ;
        RECT 2028.210 313.860 2028.530 313.920 ;
        RECT 2587.570 313.860 2587.890 313.920 ;
      LAYER via ;
        RECT 2028.240 313.860 2028.500 314.120 ;
        RECT 2587.600 313.860 2587.860 314.120 ;
      LAYER met2 ;
        RECT 2026.290 960.570 2026.570 964.000 ;
        RECT 2026.290 960.430 2028.440 960.570 ;
        RECT 2026.290 960.000 2026.570 960.430 ;
        RECT 2028.300 314.150 2028.440 960.430 ;
        RECT 2028.240 313.830 2028.500 314.150 ;
        RECT 2587.600 313.830 2587.860 314.150 ;
        RECT 2587.660 17.410 2587.800 313.830 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 801.850 945.780 802.170 945.840 ;
        RECT 806.910 945.780 807.230 945.840 ;
        RECT 801.850 945.640 807.230 945.780 ;
        RECT 801.850 945.580 802.170 945.640 ;
        RECT 806.910 945.580 807.230 945.640 ;
        RECT 806.910 17.920 807.230 17.980 ;
        RECT 823.470 17.920 823.790 17.980 ;
        RECT 806.910 17.780 823.790 17.920 ;
        RECT 806.910 17.720 807.230 17.780 ;
        RECT 823.470 17.720 823.790 17.780 ;
      LAYER via ;
        RECT 801.880 945.580 802.140 945.840 ;
        RECT 806.940 945.580 807.200 945.840 ;
        RECT 806.940 17.720 807.200 17.980 ;
        RECT 823.500 17.720 823.760 17.980 ;
      LAYER met2 ;
        RECT 801.770 960.500 802.050 964.000 ;
        RECT 801.770 960.000 802.080 960.500 ;
        RECT 801.940 945.870 802.080 960.000 ;
        RECT 801.880 945.550 802.140 945.870 ;
        RECT 806.940 945.550 807.200 945.870 ;
        RECT 807.000 18.010 807.140 945.550 ;
        RECT 806.940 17.690 807.200 18.010 ;
        RECT 823.500 17.690 823.760 18.010 ;
        RECT 823.560 2.400 823.700 17.690 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 431.360 2042.330 431.420 ;
        RECT 2601.370 431.360 2601.690 431.420 ;
        RECT 2042.010 431.220 2601.690 431.360 ;
        RECT 2042.010 431.160 2042.330 431.220 ;
        RECT 2601.370 431.160 2601.690 431.220 ;
        RECT 2601.370 17.920 2601.690 17.980 ;
        RECT 2607.350 17.920 2607.670 17.980 ;
        RECT 2601.370 17.780 2607.670 17.920 ;
        RECT 2601.370 17.720 2601.690 17.780 ;
        RECT 2607.350 17.720 2607.670 17.780 ;
      LAYER via ;
        RECT 2042.040 431.160 2042.300 431.420 ;
        RECT 2601.400 431.160 2601.660 431.420 ;
        RECT 2601.400 17.720 2601.660 17.980 ;
        RECT 2607.380 17.720 2607.640 17.980 ;
      LAYER met2 ;
        RECT 2038.710 960.570 2038.990 964.000 ;
        RECT 2038.710 960.430 2042.240 960.570 ;
        RECT 2038.710 960.000 2038.990 960.430 ;
        RECT 2042.100 431.450 2042.240 960.430 ;
        RECT 2042.040 431.130 2042.300 431.450 ;
        RECT 2601.400 431.130 2601.660 431.450 ;
        RECT 2601.460 18.010 2601.600 431.130 ;
        RECT 2601.400 17.690 2601.660 18.010 ;
        RECT 2607.380 17.690 2607.640 18.010 ;
        RECT 2607.440 2.400 2607.580 17.690 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2051.210 945.440 2051.530 945.500 ;
        RECT 2055.810 945.440 2056.130 945.500 ;
        RECT 2051.210 945.300 2056.130 945.440 ;
        RECT 2051.210 945.240 2051.530 945.300 ;
        RECT 2055.810 945.240 2056.130 945.300 ;
        RECT 2055.810 300.120 2056.130 300.180 ;
        RECT 2622.070 300.120 2622.390 300.180 ;
        RECT 2055.810 299.980 2622.390 300.120 ;
        RECT 2055.810 299.920 2056.130 299.980 ;
        RECT 2622.070 299.920 2622.390 299.980 ;
      LAYER via ;
        RECT 2051.240 945.240 2051.500 945.500 ;
        RECT 2055.840 945.240 2056.100 945.500 ;
        RECT 2055.840 299.920 2056.100 300.180 ;
        RECT 2622.100 299.920 2622.360 300.180 ;
      LAYER met2 ;
        RECT 2051.130 960.500 2051.410 964.000 ;
        RECT 2051.130 960.000 2051.440 960.500 ;
        RECT 2051.300 945.530 2051.440 960.000 ;
        RECT 2051.240 945.210 2051.500 945.530 ;
        RECT 2055.840 945.210 2056.100 945.530 ;
        RECT 2055.900 300.210 2056.040 945.210 ;
        RECT 2055.840 299.890 2056.100 300.210 ;
        RECT 2622.100 299.890 2622.360 300.210 ;
        RECT 2622.160 17.410 2622.300 299.890 ;
        RECT 2622.160 17.270 2625.520 17.410 ;
        RECT 2625.380 2.400 2625.520 17.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2063.630 946.800 2063.950 946.860 ;
        RECT 2069.610 946.800 2069.930 946.860 ;
        RECT 2063.630 946.660 2069.930 946.800 ;
        RECT 2063.630 946.600 2063.950 946.660 ;
        RECT 2069.610 946.600 2069.930 946.660 ;
        RECT 2069.610 306.920 2069.930 306.980 ;
        RECT 2643.230 306.920 2643.550 306.980 ;
        RECT 2069.610 306.780 2643.550 306.920 ;
        RECT 2069.610 306.720 2069.930 306.780 ;
        RECT 2643.230 306.720 2643.550 306.780 ;
      LAYER via ;
        RECT 2063.660 946.600 2063.920 946.860 ;
        RECT 2069.640 946.600 2069.900 946.860 ;
        RECT 2069.640 306.720 2069.900 306.980 ;
        RECT 2643.260 306.720 2643.520 306.980 ;
      LAYER met2 ;
        RECT 2063.550 960.500 2063.830 964.000 ;
        RECT 2063.550 960.000 2063.860 960.500 ;
        RECT 2063.720 946.890 2063.860 960.000 ;
        RECT 2063.660 946.570 2063.920 946.890 ;
        RECT 2069.640 946.570 2069.900 946.890 ;
        RECT 2069.700 307.010 2069.840 946.570 ;
        RECT 2069.640 306.690 2069.900 307.010 ;
        RECT 2643.260 306.690 2643.520 307.010 ;
        RECT 2643.320 2.400 2643.460 306.690 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.510 645.220 2076.830 645.280 ;
        RECT 2656.570 645.220 2656.890 645.280 ;
        RECT 2076.510 645.080 2656.890 645.220 ;
        RECT 2076.510 645.020 2076.830 645.080 ;
        RECT 2656.570 645.020 2656.890 645.080 ;
      LAYER via ;
        RECT 2076.540 645.020 2076.800 645.280 ;
        RECT 2656.600 645.020 2656.860 645.280 ;
      LAYER met2 ;
        RECT 2075.970 960.570 2076.250 964.000 ;
        RECT 2075.970 960.430 2076.740 960.570 ;
        RECT 2075.970 960.000 2076.250 960.430 ;
        RECT 2076.600 645.310 2076.740 960.430 ;
        RECT 2076.540 644.990 2076.800 645.310 ;
        RECT 2656.600 644.990 2656.860 645.310 ;
        RECT 2656.660 17.410 2656.800 644.990 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 341.600 2090.630 341.660 ;
        RECT 2677.270 341.600 2677.590 341.660 ;
        RECT 2090.310 341.460 2677.590 341.600 ;
        RECT 2090.310 341.400 2090.630 341.460 ;
        RECT 2677.270 341.400 2677.590 341.460 ;
      LAYER via ;
        RECT 2090.340 341.400 2090.600 341.660 ;
        RECT 2677.300 341.400 2677.560 341.660 ;
      LAYER met2 ;
        RECT 2088.390 960.570 2088.670 964.000 ;
        RECT 2088.390 960.430 2090.540 960.570 ;
        RECT 2088.390 960.000 2088.670 960.430 ;
        RECT 2090.400 341.690 2090.540 960.430 ;
        RECT 2090.340 341.370 2090.600 341.690 ;
        RECT 2677.300 341.370 2677.560 341.690 ;
        RECT 2677.360 17.410 2677.500 341.370 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 417.420 2104.430 417.480 ;
        RECT 2691.070 417.420 2691.390 417.480 ;
        RECT 2104.110 417.280 2691.390 417.420 ;
        RECT 2104.110 417.220 2104.430 417.280 ;
        RECT 2691.070 417.220 2691.390 417.280 ;
      LAYER via ;
        RECT 2104.140 417.220 2104.400 417.480 ;
        RECT 2691.100 417.220 2691.360 417.480 ;
      LAYER met2 ;
        RECT 2100.810 960.570 2101.090 964.000 ;
        RECT 2100.810 960.430 2104.340 960.570 ;
        RECT 2100.810 960.000 2101.090 960.430 ;
        RECT 2104.200 417.510 2104.340 960.430 ;
        RECT 2104.140 417.190 2104.400 417.510 ;
        RECT 2691.100 417.190 2691.360 417.510 ;
        RECT 2691.160 17.410 2691.300 417.190 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2113.310 945.440 2113.630 945.500 ;
        RECT 2117.450 945.440 2117.770 945.500 ;
        RECT 2113.310 945.300 2117.770 945.440 ;
        RECT 2113.310 945.240 2113.630 945.300 ;
        RECT 2117.450 945.240 2117.770 945.300 ;
        RECT 2117.450 638.080 2117.770 638.140 ;
        RECT 2711.770 638.080 2712.090 638.140 ;
        RECT 2117.450 637.940 2712.090 638.080 ;
        RECT 2117.450 637.880 2117.770 637.940 ;
        RECT 2711.770 637.880 2712.090 637.940 ;
      LAYER via ;
        RECT 2113.340 945.240 2113.600 945.500 ;
        RECT 2117.480 945.240 2117.740 945.500 ;
        RECT 2117.480 637.880 2117.740 638.140 ;
        RECT 2711.800 637.880 2712.060 638.140 ;
      LAYER met2 ;
        RECT 2113.230 960.500 2113.510 964.000 ;
        RECT 2113.230 960.000 2113.540 960.500 ;
        RECT 2113.400 945.530 2113.540 960.000 ;
        RECT 2113.340 945.210 2113.600 945.530 ;
        RECT 2117.480 945.210 2117.740 945.530 ;
        RECT 2117.540 638.170 2117.680 945.210 ;
        RECT 2117.480 637.850 2117.740 638.170 ;
        RECT 2711.800 637.850 2712.060 638.170 ;
        RECT 2711.860 17.410 2712.000 637.850 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2125.730 946.460 2126.050 946.520 ;
        RECT 2131.710 946.460 2132.030 946.520 ;
        RECT 2125.730 946.320 2132.030 946.460 ;
        RECT 2125.730 946.260 2126.050 946.320 ;
        RECT 2131.710 946.260 2132.030 946.320 ;
        RECT 2131.710 327.660 2132.030 327.720 ;
        RECT 2732.930 327.660 2733.250 327.720 ;
        RECT 2131.710 327.520 2733.250 327.660 ;
        RECT 2131.710 327.460 2132.030 327.520 ;
        RECT 2732.930 327.460 2733.250 327.520 ;
      LAYER via ;
        RECT 2125.760 946.260 2126.020 946.520 ;
        RECT 2131.740 946.260 2132.000 946.520 ;
        RECT 2131.740 327.460 2132.000 327.720 ;
        RECT 2732.960 327.460 2733.220 327.720 ;
      LAYER met2 ;
        RECT 2125.650 960.500 2125.930 964.000 ;
        RECT 2125.650 960.000 2125.960 960.500 ;
        RECT 2125.820 946.550 2125.960 960.000 ;
        RECT 2125.760 946.230 2126.020 946.550 ;
        RECT 2131.740 946.230 2132.000 946.550 ;
        RECT 2131.800 327.750 2131.940 946.230 ;
        RECT 2131.740 327.430 2132.000 327.750 ;
        RECT 2732.960 327.430 2733.220 327.750 ;
        RECT 2733.020 17.410 2733.160 327.430 ;
        RECT 2732.560 17.270 2733.160 17.410 ;
        RECT 2732.560 2.400 2732.700 17.270 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2138.610 424.220 2138.930 424.280 ;
        RECT 2746.270 424.220 2746.590 424.280 ;
        RECT 2138.610 424.080 2746.590 424.220 ;
        RECT 2138.610 424.020 2138.930 424.080 ;
        RECT 2746.270 424.020 2746.590 424.080 ;
      LAYER via ;
        RECT 2138.640 424.020 2138.900 424.280 ;
        RECT 2746.300 424.020 2746.560 424.280 ;
      LAYER met2 ;
        RECT 2138.070 960.570 2138.350 964.000 ;
        RECT 2138.070 960.430 2138.840 960.570 ;
        RECT 2138.070 960.000 2138.350 960.430 ;
        RECT 2138.700 424.310 2138.840 960.430 ;
        RECT 2138.640 423.990 2138.900 424.310 ;
        RECT 2746.300 423.990 2746.560 424.310 ;
        RECT 2746.360 17.410 2746.500 423.990 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.410 334.460 2152.730 334.520 ;
        RECT 2766.970 334.460 2767.290 334.520 ;
        RECT 2152.410 334.320 2767.290 334.460 ;
        RECT 2152.410 334.260 2152.730 334.320 ;
        RECT 2766.970 334.260 2767.290 334.320 ;
      LAYER via ;
        RECT 2152.440 334.260 2152.700 334.520 ;
        RECT 2767.000 334.260 2767.260 334.520 ;
      LAYER met2 ;
        RECT 2150.030 960.570 2150.310 964.000 ;
        RECT 2150.030 960.430 2152.640 960.570 ;
        RECT 2150.030 960.000 2150.310 960.430 ;
        RECT 2152.500 334.550 2152.640 960.430 ;
        RECT 2152.440 334.230 2152.700 334.550 ;
        RECT 2767.000 334.230 2767.260 334.550 ;
        RECT 2767.060 17.410 2767.200 334.230 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 814.270 949.860 814.590 949.920 ;
        RECT 820.250 949.860 820.570 949.920 ;
        RECT 814.270 949.720 820.570 949.860 ;
        RECT 814.270 949.660 814.590 949.720 ;
        RECT 820.250 949.660 820.570 949.720 ;
        RECT 820.250 16.560 820.570 16.620 ;
        RECT 840.950 16.560 841.270 16.620 ;
        RECT 820.250 16.420 841.270 16.560 ;
        RECT 820.250 16.360 820.570 16.420 ;
        RECT 840.950 16.360 841.270 16.420 ;
      LAYER via ;
        RECT 814.300 949.660 814.560 949.920 ;
        RECT 820.280 949.660 820.540 949.920 ;
        RECT 820.280 16.360 820.540 16.620 ;
        RECT 840.980 16.360 841.240 16.620 ;
      LAYER met2 ;
        RECT 814.190 960.500 814.470 964.000 ;
        RECT 814.190 960.000 814.500 960.500 ;
        RECT 814.360 949.950 814.500 960.000 ;
        RECT 814.300 949.630 814.560 949.950 ;
        RECT 820.280 949.630 820.540 949.950 ;
        RECT 820.340 16.650 820.480 949.630 ;
        RECT 820.280 16.330 820.540 16.650 ;
        RECT 840.980 16.330 841.240 16.650 ;
        RECT 841.040 2.400 841.180 16.330 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 631.280 2166.530 631.340 ;
        RECT 2780.770 631.280 2781.090 631.340 ;
        RECT 2166.210 631.140 2781.090 631.280 ;
        RECT 2166.210 631.080 2166.530 631.140 ;
        RECT 2780.770 631.080 2781.090 631.140 ;
      LAYER via ;
        RECT 2166.240 631.080 2166.500 631.340 ;
        RECT 2780.800 631.080 2781.060 631.340 ;
      LAYER met2 ;
        RECT 2162.450 960.570 2162.730 964.000 ;
        RECT 2162.450 960.430 2166.440 960.570 ;
        RECT 2162.450 960.000 2162.730 960.430 ;
        RECT 2166.300 631.370 2166.440 960.430 ;
        RECT 2166.240 631.050 2166.500 631.370 ;
        RECT 2780.800 631.050 2781.060 631.370 ;
        RECT 2780.860 17.410 2781.000 631.050 ;
        RECT 2780.860 17.270 2786.060 17.410 ;
        RECT 2785.920 2.400 2786.060 17.270 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2174.950 951.220 2175.270 951.280 ;
        RECT 2179.550 951.220 2179.870 951.280 ;
        RECT 2174.950 951.080 2179.870 951.220 ;
        RECT 2174.950 951.020 2175.270 951.080 ;
        RECT 2179.550 951.020 2179.870 951.080 ;
        RECT 2179.550 624.480 2179.870 624.540 ;
        RECT 2801.470 624.480 2801.790 624.540 ;
        RECT 2179.550 624.340 2801.790 624.480 ;
        RECT 2179.550 624.280 2179.870 624.340 ;
        RECT 2801.470 624.280 2801.790 624.340 ;
      LAYER via ;
        RECT 2174.980 951.020 2175.240 951.280 ;
        RECT 2179.580 951.020 2179.840 951.280 ;
        RECT 2179.580 624.280 2179.840 624.540 ;
        RECT 2801.500 624.280 2801.760 624.540 ;
      LAYER met2 ;
        RECT 2174.870 960.500 2175.150 964.000 ;
        RECT 2174.870 960.000 2175.180 960.500 ;
        RECT 2175.040 951.310 2175.180 960.000 ;
        RECT 2174.980 950.990 2175.240 951.310 ;
        RECT 2179.580 950.990 2179.840 951.310 ;
        RECT 2179.640 624.570 2179.780 950.990 ;
        RECT 2179.580 624.250 2179.840 624.570 ;
        RECT 2801.500 624.250 2801.760 624.570 ;
        RECT 2801.560 17.410 2801.700 624.250 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2187.370 946.460 2187.690 946.520 ;
        RECT 2193.810 946.460 2194.130 946.520 ;
        RECT 2187.370 946.320 2194.130 946.460 ;
        RECT 2187.370 946.260 2187.690 946.320 ;
        RECT 2193.810 946.260 2194.130 946.320 ;
        RECT 2193.810 348.400 2194.130 348.460 ;
        RECT 2815.730 348.400 2816.050 348.460 ;
        RECT 2193.810 348.260 2816.050 348.400 ;
        RECT 2193.810 348.200 2194.130 348.260 ;
        RECT 2815.730 348.200 2816.050 348.260 ;
        RECT 2815.730 17.920 2816.050 17.980 ;
        RECT 2821.710 17.920 2822.030 17.980 ;
        RECT 2815.730 17.780 2822.030 17.920 ;
        RECT 2815.730 17.720 2816.050 17.780 ;
        RECT 2821.710 17.720 2822.030 17.780 ;
      LAYER via ;
        RECT 2187.400 946.260 2187.660 946.520 ;
        RECT 2193.840 946.260 2194.100 946.520 ;
        RECT 2193.840 348.200 2194.100 348.460 ;
        RECT 2815.760 348.200 2816.020 348.460 ;
        RECT 2815.760 17.720 2816.020 17.980 ;
        RECT 2821.740 17.720 2822.000 17.980 ;
      LAYER met2 ;
        RECT 2187.290 960.500 2187.570 964.000 ;
        RECT 2187.290 960.000 2187.600 960.500 ;
        RECT 2187.460 946.550 2187.600 960.000 ;
        RECT 2187.400 946.230 2187.660 946.550 ;
        RECT 2193.840 946.230 2194.100 946.550 ;
        RECT 2193.900 348.490 2194.040 946.230 ;
        RECT 2193.840 348.170 2194.100 348.490 ;
        RECT 2815.760 348.170 2816.020 348.490 ;
        RECT 2815.820 18.010 2815.960 348.170 ;
        RECT 2815.760 17.690 2816.020 18.010 ;
        RECT 2821.740 17.690 2822.000 18.010 ;
        RECT 2821.800 2.400 2821.940 17.690 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2200.710 355.200 2201.030 355.260 ;
        RECT 2835.970 355.200 2836.290 355.260 ;
        RECT 2200.710 355.060 2836.290 355.200 ;
        RECT 2200.710 355.000 2201.030 355.060 ;
        RECT 2835.970 355.000 2836.290 355.060 ;
      LAYER via ;
        RECT 2200.740 355.000 2201.000 355.260 ;
        RECT 2836.000 355.000 2836.260 355.260 ;
      LAYER met2 ;
        RECT 2199.710 960.570 2199.990 964.000 ;
        RECT 2199.710 960.430 2200.940 960.570 ;
        RECT 2199.710 960.000 2199.990 960.430 ;
        RECT 2200.800 355.290 2200.940 960.430 ;
        RECT 2200.740 354.970 2201.000 355.290 ;
        RECT 2836.000 354.970 2836.260 355.290 ;
        RECT 2836.060 17.410 2836.200 354.970 ;
        RECT 2836.060 17.270 2839.420 17.410 ;
        RECT 2839.280 2.400 2839.420 17.270 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 362.340 2214.830 362.400 ;
        RECT 2857.130 362.340 2857.450 362.400 ;
        RECT 2214.510 362.200 2857.450 362.340 ;
        RECT 2214.510 362.140 2214.830 362.200 ;
        RECT 2857.130 362.140 2857.450 362.200 ;
      LAYER via ;
        RECT 2214.540 362.140 2214.800 362.400 ;
        RECT 2857.160 362.140 2857.420 362.400 ;
      LAYER met2 ;
        RECT 2212.130 960.570 2212.410 964.000 ;
        RECT 2212.130 960.430 2214.740 960.570 ;
        RECT 2212.130 960.000 2212.410 960.430 ;
        RECT 2214.600 362.430 2214.740 960.430 ;
        RECT 2214.540 362.110 2214.800 362.430 ;
        RECT 2857.160 362.110 2857.420 362.430 ;
        RECT 2857.220 2.400 2857.360 362.110 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2224.630 945.440 2224.950 945.500 ;
        RECT 2228.310 945.440 2228.630 945.500 ;
        RECT 2224.630 945.300 2228.630 945.440 ;
        RECT 2224.630 945.240 2224.950 945.300 ;
        RECT 2228.310 945.240 2228.630 945.300 ;
        RECT 2228.310 396.680 2228.630 396.740 ;
        RECT 2870.470 396.680 2870.790 396.740 ;
        RECT 2228.310 396.540 2870.790 396.680 ;
        RECT 2228.310 396.480 2228.630 396.540 ;
        RECT 2870.470 396.480 2870.790 396.540 ;
      LAYER via ;
        RECT 2224.660 945.240 2224.920 945.500 ;
        RECT 2228.340 945.240 2228.600 945.500 ;
        RECT 2228.340 396.480 2228.600 396.740 ;
        RECT 2870.500 396.480 2870.760 396.740 ;
      LAYER met2 ;
        RECT 2224.550 960.500 2224.830 964.000 ;
        RECT 2224.550 960.000 2224.860 960.500 ;
        RECT 2224.720 945.530 2224.860 960.000 ;
        RECT 2224.660 945.210 2224.920 945.530 ;
        RECT 2228.340 945.210 2228.600 945.530 ;
        RECT 2228.400 396.770 2228.540 945.210 ;
        RECT 2228.340 396.450 2228.600 396.770 ;
        RECT 2870.500 396.450 2870.760 396.770 ;
        RECT 2870.560 17.410 2870.700 396.450 ;
        RECT 2870.560 17.270 2875.300 17.410 ;
        RECT 2875.160 2.400 2875.300 17.270 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2237.050 945.440 2237.370 945.500 ;
        RECT 2242.110 945.440 2242.430 945.500 ;
        RECT 2237.050 945.300 2242.430 945.440 ;
        RECT 2237.050 945.240 2237.370 945.300 ;
        RECT 2242.110 945.240 2242.430 945.300 ;
        RECT 2242.110 17.580 2242.430 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2242.110 17.440 2893.330 17.580 ;
        RECT 2242.110 17.380 2242.430 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 2237.080 945.240 2237.340 945.500 ;
        RECT 2242.140 945.240 2242.400 945.500 ;
        RECT 2242.140 17.380 2242.400 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 2236.970 960.500 2237.250 964.000 ;
        RECT 2236.970 960.000 2237.280 960.500 ;
        RECT 2237.140 945.530 2237.280 960.000 ;
        RECT 2237.080 945.210 2237.340 945.530 ;
        RECT 2242.140 945.210 2242.400 945.530 ;
        RECT 2242.200 17.670 2242.340 945.210 ;
        RECT 2242.140 17.350 2242.400 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2249.470 945.440 2249.790 945.500 ;
        RECT 2255.910 945.440 2256.230 945.500 ;
        RECT 2249.470 945.300 2256.230 945.440 ;
        RECT 2249.470 945.240 2249.790 945.300 ;
        RECT 2255.910 945.240 2256.230 945.300 ;
        RECT 2255.910 17.240 2256.230 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2255.910 17.100 2911.270 17.240 ;
        RECT 2255.910 17.040 2256.230 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 2249.500 945.240 2249.760 945.500 ;
        RECT 2255.940 945.240 2256.200 945.500 ;
        RECT 2255.940 17.040 2256.200 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 2249.390 960.500 2249.670 964.000 ;
        RECT 2249.390 960.000 2249.700 960.500 ;
        RECT 2249.560 945.530 2249.700 960.000 ;
        RECT 2249.500 945.210 2249.760 945.530 ;
        RECT 2255.940 945.210 2256.200 945.530 ;
        RECT 2256.000 17.330 2256.140 945.210 ;
        RECT 2255.940 17.010 2256.200 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 15.200 827.930 15.260 ;
        RECT 858.890 15.200 859.210 15.260 ;
        RECT 827.610 15.060 859.210 15.200 ;
        RECT 827.610 15.000 827.930 15.060 ;
        RECT 858.890 15.000 859.210 15.060 ;
      LAYER via ;
        RECT 827.640 15.000 827.900 15.260 ;
        RECT 858.920 15.000 859.180 15.260 ;
      LAYER met2 ;
        RECT 826.610 960.570 826.890 964.000 ;
        RECT 826.610 960.430 827.840 960.570 ;
        RECT 826.610 960.000 826.890 960.430 ;
        RECT 827.700 15.290 827.840 960.430 ;
        RECT 827.640 14.970 827.900 15.290 ;
        RECT 858.920 14.970 859.180 15.290 ;
        RECT 858.980 2.400 859.120 14.970 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 17.580 841.730 17.640 ;
        RECT 876.830 17.580 877.150 17.640 ;
        RECT 841.410 17.440 877.150 17.580 ;
        RECT 841.410 17.380 841.730 17.440 ;
        RECT 876.830 17.380 877.150 17.440 ;
      LAYER via ;
        RECT 841.440 17.380 841.700 17.640 ;
        RECT 876.860 17.380 877.120 17.640 ;
      LAYER met2 ;
        RECT 839.030 960.570 839.310 964.000 ;
        RECT 839.030 960.430 841.640 960.570 ;
        RECT 839.030 960.000 839.310 960.430 ;
        RECT 841.500 17.670 841.640 960.430 ;
        RECT 841.440 17.350 841.700 17.670 ;
        RECT 876.860 17.350 877.120 17.670 ;
        RECT 876.920 2.400 877.060 17.350 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.210 17.240 855.530 17.300 ;
        RECT 894.770 17.240 895.090 17.300 ;
        RECT 855.210 17.100 895.090 17.240 ;
        RECT 855.210 17.040 855.530 17.100 ;
        RECT 894.770 17.040 895.090 17.100 ;
      LAYER via ;
        RECT 855.240 17.040 855.500 17.300 ;
        RECT 894.800 17.040 895.060 17.300 ;
      LAYER met2 ;
        RECT 851.450 960.570 851.730 964.000 ;
        RECT 851.450 960.430 855.440 960.570 ;
        RECT 851.450 960.000 851.730 960.430 ;
        RECT 855.300 17.330 855.440 960.430 ;
        RECT 855.240 17.010 855.500 17.330 ;
        RECT 894.800 17.010 895.060 17.330 ;
        RECT 894.860 2.400 895.000 17.010 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 863.950 946.800 864.270 946.860 ;
        RECT 869.010 946.800 869.330 946.860 ;
        RECT 863.950 946.660 869.330 946.800 ;
        RECT 863.950 946.600 864.270 946.660 ;
        RECT 869.010 946.600 869.330 946.660 ;
        RECT 912.710 18.940 913.030 19.000 ;
        RECT 889.340 18.800 913.030 18.940 ;
        RECT 869.010 18.600 869.330 18.660 ;
        RECT 889.340 18.600 889.480 18.800 ;
        RECT 912.710 18.740 913.030 18.800 ;
        RECT 869.010 18.460 889.480 18.600 ;
        RECT 869.010 18.400 869.330 18.460 ;
      LAYER via ;
        RECT 863.980 946.600 864.240 946.860 ;
        RECT 869.040 946.600 869.300 946.860 ;
        RECT 869.040 18.400 869.300 18.660 ;
        RECT 912.740 18.740 913.000 19.000 ;
      LAYER met2 ;
        RECT 863.870 960.500 864.150 964.000 ;
        RECT 863.870 960.000 864.180 960.500 ;
        RECT 864.040 946.890 864.180 960.000 ;
        RECT 863.980 946.570 864.240 946.890 ;
        RECT 869.040 946.570 869.300 946.890 ;
        RECT 869.100 18.690 869.240 946.570 ;
        RECT 912.740 18.710 913.000 19.030 ;
        RECT 869.040 18.370 869.300 18.690 ;
        RECT 912.800 2.400 912.940 18.710 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.370 946.460 876.690 946.520 ;
        RECT 882.810 946.460 883.130 946.520 ;
        RECT 876.370 946.320 883.130 946.460 ;
        RECT 876.370 946.260 876.690 946.320 ;
        RECT 882.810 946.260 883.130 946.320 ;
        RECT 882.810 19.960 883.130 20.020 ;
        RECT 930.190 19.960 930.510 20.020 ;
        RECT 882.810 19.820 930.510 19.960 ;
        RECT 882.810 19.760 883.130 19.820 ;
        RECT 930.190 19.760 930.510 19.820 ;
      LAYER via ;
        RECT 876.400 946.260 876.660 946.520 ;
        RECT 882.840 946.260 883.100 946.520 ;
        RECT 882.840 19.760 883.100 20.020 ;
        RECT 930.220 19.760 930.480 20.020 ;
      LAYER met2 ;
        RECT 876.290 960.500 876.570 964.000 ;
        RECT 876.290 960.000 876.600 960.500 ;
        RECT 876.460 946.550 876.600 960.000 ;
        RECT 876.400 946.230 876.660 946.550 ;
        RECT 882.840 946.230 883.100 946.550 ;
        RECT 882.900 20.050 883.040 946.230 ;
        RECT 882.840 19.730 883.100 20.050 ;
        RECT 930.220 19.730 930.480 20.050 ;
        RECT 930.280 2.400 930.420 19.730 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 889.710 17.580 890.030 17.640 ;
        RECT 948.130 17.580 948.450 17.640 ;
        RECT 889.710 17.440 948.450 17.580 ;
        RECT 889.710 17.380 890.030 17.440 ;
        RECT 948.130 17.380 948.450 17.440 ;
      LAYER via ;
        RECT 889.740 17.380 890.000 17.640 ;
        RECT 948.160 17.380 948.420 17.640 ;
      LAYER met2 ;
        RECT 888.710 960.570 888.990 964.000 ;
        RECT 888.710 960.430 889.940 960.570 ;
        RECT 888.710 960.000 888.990 960.430 ;
        RECT 889.800 17.670 889.940 960.430 ;
        RECT 889.740 17.350 890.000 17.670 ;
        RECT 948.160 17.350 948.420 17.670 ;
        RECT 948.220 2.400 948.360 17.350 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.510 18.600 903.830 18.660 ;
        RECT 966.070 18.600 966.390 18.660 ;
        RECT 903.510 18.460 966.390 18.600 ;
        RECT 903.510 18.400 903.830 18.460 ;
        RECT 966.070 18.400 966.390 18.460 ;
      LAYER via ;
        RECT 903.540 18.400 903.800 18.660 ;
        RECT 966.100 18.400 966.360 18.660 ;
      LAYER met2 ;
        RECT 900.670 960.570 900.950 964.000 ;
        RECT 900.670 960.430 903.740 960.570 ;
        RECT 900.670 960.000 900.950 960.430 ;
        RECT 903.600 18.690 903.740 960.430 ;
        RECT 903.540 18.370 903.800 18.690 ;
        RECT 966.100 18.370 966.360 18.690 ;
        RECT 966.160 2.400 966.300 18.370 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 913.170 947.140 913.490 947.200 ;
        RECT 917.310 947.140 917.630 947.200 ;
        RECT 913.170 947.000 917.630 947.140 ;
        RECT 913.170 946.940 913.490 947.000 ;
        RECT 917.310 946.940 917.630 947.000 ;
        RECT 917.310 18.940 917.630 19.000 ;
        RECT 984.010 18.940 984.330 19.000 ;
        RECT 917.310 18.800 984.330 18.940 ;
        RECT 917.310 18.740 917.630 18.800 ;
        RECT 984.010 18.740 984.330 18.800 ;
      LAYER via ;
        RECT 913.200 946.940 913.460 947.200 ;
        RECT 917.340 946.940 917.600 947.200 ;
        RECT 917.340 18.740 917.600 19.000 ;
        RECT 984.040 18.740 984.300 19.000 ;
      LAYER met2 ;
        RECT 913.090 960.500 913.370 964.000 ;
        RECT 913.090 960.000 913.400 960.500 ;
        RECT 913.260 947.230 913.400 960.000 ;
        RECT 913.200 946.910 913.460 947.230 ;
        RECT 917.340 946.910 917.600 947.230 ;
        RECT 917.400 19.030 917.540 946.910 ;
        RECT 917.340 18.710 917.600 19.030 ;
        RECT 984.040 18.710 984.300 19.030 ;
        RECT 984.100 2.400 984.240 18.710 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 17.920 663.250 17.980 ;
        RECT 690.070 17.920 690.390 17.980 ;
        RECT 662.930 17.780 690.390 17.920 ;
        RECT 662.930 17.720 663.250 17.780 ;
        RECT 690.070 17.720 690.390 17.780 ;
      LAYER via ;
        RECT 662.960 17.720 663.220 17.980 ;
        RECT 690.100 17.720 690.360 17.980 ;
      LAYER met2 ;
        RECT 690.450 960.570 690.730 964.000 ;
        RECT 690.160 960.430 690.730 960.570 ;
        RECT 690.160 18.010 690.300 960.430 ;
        RECT 690.450 960.000 690.730 960.430 ;
        RECT 662.960 17.690 663.220 18.010 ;
        RECT 690.100 17.690 690.360 18.010 ;
        RECT 663.020 2.400 663.160 17.690 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 925.590 946.460 925.910 946.520 ;
        RECT 931.110 946.460 931.430 946.520 ;
        RECT 925.590 946.320 931.430 946.460 ;
        RECT 925.590 946.260 925.910 946.320 ;
        RECT 931.110 946.260 931.430 946.320 ;
        RECT 931.110 18.260 931.430 18.320 ;
        RECT 1001.950 18.260 1002.270 18.320 ;
        RECT 931.110 18.120 1002.270 18.260 ;
        RECT 931.110 18.060 931.430 18.120 ;
        RECT 1001.950 18.060 1002.270 18.120 ;
      LAYER via ;
        RECT 925.620 946.260 925.880 946.520 ;
        RECT 931.140 946.260 931.400 946.520 ;
        RECT 931.140 18.060 931.400 18.320 ;
        RECT 1001.980 18.060 1002.240 18.320 ;
      LAYER met2 ;
        RECT 925.510 960.500 925.790 964.000 ;
        RECT 925.510 960.000 925.820 960.500 ;
        RECT 925.680 946.550 925.820 960.000 ;
        RECT 925.620 946.230 925.880 946.550 ;
        RECT 931.140 946.230 931.400 946.550 ;
        RECT 931.200 18.350 931.340 946.230 ;
        RECT 931.140 18.030 931.400 18.350 ;
        RECT 1001.980 18.030 1002.240 18.350 ;
        RECT 1002.040 2.400 1002.180 18.030 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.010 17.920 938.330 17.980 ;
        RECT 1019.430 17.920 1019.750 17.980 ;
        RECT 938.010 17.780 1019.750 17.920 ;
        RECT 938.010 17.720 938.330 17.780 ;
        RECT 1019.430 17.720 1019.750 17.780 ;
      LAYER via ;
        RECT 938.040 17.720 938.300 17.980 ;
        RECT 1019.460 17.720 1019.720 17.980 ;
      LAYER met2 ;
        RECT 937.930 960.500 938.210 964.000 ;
        RECT 937.930 960.000 938.240 960.500 ;
        RECT 938.100 18.010 938.240 960.000 ;
        RECT 938.040 17.690 938.300 18.010 ;
        RECT 1019.460 17.690 1019.720 18.010 ;
        RECT 1019.520 2.400 1019.660 17.690 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1007.085 16.745 1007.255 17.595 ;
      LAYER mcon ;
        RECT 1007.085 17.425 1007.255 17.595 ;
      LAYER met1 ;
        RECT 951.810 17.580 952.130 17.640 ;
        RECT 1007.025 17.580 1007.315 17.625 ;
        RECT 951.810 17.440 1007.315 17.580 ;
        RECT 951.810 17.380 952.130 17.440 ;
        RECT 1007.025 17.395 1007.315 17.440 ;
        RECT 1007.025 16.900 1007.315 16.945 ;
        RECT 1037.370 16.900 1037.690 16.960 ;
        RECT 1007.025 16.760 1037.690 16.900 ;
        RECT 1007.025 16.715 1007.315 16.760 ;
        RECT 1037.370 16.700 1037.690 16.760 ;
      LAYER via ;
        RECT 951.840 17.380 952.100 17.640 ;
        RECT 1037.400 16.700 1037.660 16.960 ;
      LAYER met2 ;
        RECT 950.350 960.570 950.630 964.000 ;
        RECT 950.350 960.430 952.040 960.570 ;
        RECT 950.350 960.000 950.630 960.430 ;
        RECT 951.900 17.670 952.040 960.430 ;
        RECT 951.840 17.350 952.100 17.670 ;
        RECT 1037.400 16.670 1037.660 16.990 ;
        RECT 1037.460 2.400 1037.600 16.670 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 965.610 17.240 965.930 17.300 ;
        RECT 1055.310 17.240 1055.630 17.300 ;
        RECT 965.610 17.100 1055.630 17.240 ;
        RECT 965.610 17.040 965.930 17.100 ;
        RECT 1055.310 17.040 1055.630 17.100 ;
      LAYER via ;
        RECT 965.640 17.040 965.900 17.300 ;
        RECT 1055.340 17.040 1055.600 17.300 ;
      LAYER met2 ;
        RECT 962.770 960.570 963.050 964.000 ;
        RECT 962.770 960.430 965.840 960.570 ;
        RECT 962.770 960.000 963.050 960.430 ;
        RECT 965.700 17.330 965.840 960.430 ;
        RECT 965.640 17.010 965.900 17.330 ;
        RECT 1055.340 17.010 1055.600 17.330 ;
        RECT 1055.400 2.400 1055.540 17.010 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 975.270 945.440 975.590 945.500 ;
        RECT 979.410 945.440 979.730 945.500 ;
        RECT 975.270 945.300 979.730 945.440 ;
        RECT 975.270 945.240 975.590 945.300 ;
        RECT 979.410 945.240 979.730 945.300 ;
        RECT 979.410 19.620 979.730 19.680 ;
        RECT 1073.250 19.620 1073.570 19.680 ;
        RECT 979.410 19.480 1073.570 19.620 ;
        RECT 979.410 19.420 979.730 19.480 ;
        RECT 1073.250 19.420 1073.570 19.480 ;
      LAYER via ;
        RECT 975.300 945.240 975.560 945.500 ;
        RECT 979.440 945.240 979.700 945.500 ;
        RECT 979.440 19.420 979.700 19.680 ;
        RECT 1073.280 19.420 1073.540 19.680 ;
      LAYER met2 ;
        RECT 975.190 960.500 975.470 964.000 ;
        RECT 975.190 960.000 975.500 960.500 ;
        RECT 975.360 945.530 975.500 960.000 ;
        RECT 975.300 945.210 975.560 945.530 ;
        RECT 979.440 945.210 979.700 945.530 ;
        RECT 979.500 19.710 979.640 945.210 ;
        RECT 979.440 19.390 979.700 19.710 ;
        RECT 1073.280 19.390 1073.540 19.710 ;
        RECT 1073.340 2.400 1073.480 19.390 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 987.690 946.800 988.010 946.860 ;
        RECT 993.210 946.800 993.530 946.860 ;
        RECT 987.690 946.660 993.530 946.800 ;
        RECT 987.690 946.600 988.010 946.660 ;
        RECT 993.210 946.600 993.530 946.660 ;
        RECT 993.210 19.280 993.530 19.340 ;
        RECT 1090.730 19.280 1091.050 19.340 ;
        RECT 993.210 19.140 1091.050 19.280 ;
        RECT 993.210 19.080 993.530 19.140 ;
        RECT 1090.730 19.080 1091.050 19.140 ;
      LAYER via ;
        RECT 987.720 946.600 987.980 946.860 ;
        RECT 993.240 946.600 993.500 946.860 ;
        RECT 993.240 19.080 993.500 19.340 ;
        RECT 1090.760 19.080 1091.020 19.340 ;
      LAYER met2 ;
        RECT 987.610 960.500 987.890 964.000 ;
        RECT 987.610 960.000 987.920 960.500 ;
        RECT 987.780 946.890 987.920 960.000 ;
        RECT 987.720 946.570 987.980 946.890 ;
        RECT 993.240 946.570 993.500 946.890 ;
        RECT 993.300 19.370 993.440 946.570 ;
        RECT 993.240 19.050 993.500 19.370 ;
        RECT 1090.760 19.050 1091.020 19.370 ;
        RECT 1090.820 2.400 1090.960 19.050 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.110 18.940 1000.430 19.000 ;
        RECT 1108.670 18.940 1108.990 19.000 ;
        RECT 1000.110 18.800 1108.990 18.940 ;
        RECT 1000.110 18.740 1000.430 18.800 ;
        RECT 1108.670 18.740 1108.990 18.800 ;
      LAYER via ;
        RECT 1000.140 18.740 1000.400 19.000 ;
        RECT 1108.700 18.740 1108.960 19.000 ;
      LAYER met2 ;
        RECT 1000.030 960.500 1000.310 964.000 ;
        RECT 1000.030 960.000 1000.340 960.500 ;
        RECT 1000.200 19.030 1000.340 960.000 ;
        RECT 1000.140 18.710 1000.400 19.030 ;
        RECT 1108.700 18.710 1108.960 19.030 ;
        RECT 1108.760 2.400 1108.900 18.710 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1013.910 18.260 1014.230 18.320 ;
        RECT 1126.610 18.260 1126.930 18.320 ;
        RECT 1013.910 18.120 1126.930 18.260 ;
        RECT 1013.910 18.060 1014.230 18.120 ;
        RECT 1126.610 18.060 1126.930 18.120 ;
      LAYER via ;
        RECT 1013.940 18.060 1014.200 18.320 ;
        RECT 1126.640 18.060 1126.900 18.320 ;
      LAYER met2 ;
        RECT 1011.990 960.570 1012.270 964.000 ;
        RECT 1011.990 960.430 1014.140 960.570 ;
        RECT 1011.990 960.000 1012.270 960.430 ;
        RECT 1014.000 18.350 1014.140 960.430 ;
        RECT 1013.940 18.030 1014.200 18.350 ;
        RECT 1126.640 18.030 1126.900 18.350 ;
        RECT 1126.700 2.400 1126.840 18.030 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 18.600 1028.030 18.660 ;
        RECT 1144.550 18.600 1144.870 18.660 ;
        RECT 1027.710 18.460 1144.870 18.600 ;
        RECT 1027.710 18.400 1028.030 18.460 ;
        RECT 1144.550 18.400 1144.870 18.460 ;
      LAYER via ;
        RECT 1027.740 18.400 1028.000 18.660 ;
        RECT 1144.580 18.400 1144.840 18.660 ;
      LAYER met2 ;
        RECT 1024.410 960.570 1024.690 964.000 ;
        RECT 1024.410 960.430 1027.940 960.570 ;
        RECT 1024.410 960.000 1024.690 960.430 ;
        RECT 1027.800 18.690 1027.940 960.430 ;
        RECT 1027.740 18.370 1028.000 18.690 ;
        RECT 1144.580 18.370 1144.840 18.690 ;
        RECT 1144.640 2.400 1144.780 18.370 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1036.910 945.440 1037.230 945.500 ;
        RECT 1041.510 945.440 1041.830 945.500 ;
        RECT 1036.910 945.300 1041.830 945.440 ;
        RECT 1036.910 945.240 1037.230 945.300 ;
        RECT 1041.510 945.240 1041.830 945.300 ;
        RECT 1041.510 17.920 1041.830 17.980 ;
        RECT 1162.490 17.920 1162.810 17.980 ;
        RECT 1041.510 17.780 1162.810 17.920 ;
        RECT 1041.510 17.720 1041.830 17.780 ;
        RECT 1162.490 17.720 1162.810 17.780 ;
      LAYER via ;
        RECT 1036.940 945.240 1037.200 945.500 ;
        RECT 1041.540 945.240 1041.800 945.500 ;
        RECT 1041.540 17.720 1041.800 17.980 ;
        RECT 1162.520 17.720 1162.780 17.980 ;
      LAYER met2 ;
        RECT 1036.830 960.500 1037.110 964.000 ;
        RECT 1036.830 960.000 1037.140 960.500 ;
        RECT 1037.000 945.530 1037.140 960.000 ;
        RECT 1036.940 945.210 1037.200 945.530 ;
        RECT 1041.540 945.210 1041.800 945.530 ;
        RECT 1041.600 18.010 1041.740 945.210 ;
        RECT 1041.540 17.690 1041.800 18.010 ;
        RECT 1162.520 17.690 1162.780 18.010 ;
        RECT 1162.580 2.400 1162.720 17.690 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 680.410 16.900 680.730 16.960 ;
        RECT 697.430 16.900 697.750 16.960 ;
        RECT 680.410 16.760 697.750 16.900 ;
        RECT 680.410 16.700 680.730 16.760 ;
        RECT 697.430 16.700 697.750 16.760 ;
      LAYER via ;
        RECT 680.440 16.700 680.700 16.960 ;
        RECT 697.460 16.700 697.720 16.960 ;
      LAYER met2 ;
        RECT 702.870 961.250 703.150 964.000 ;
        RECT 699.360 961.110 703.150 961.250 ;
        RECT 699.360 946.290 699.500 961.110 ;
        RECT 702.870 960.000 703.150 961.110 ;
        RECT 698.900 946.150 699.500 946.290 ;
        RECT 698.900 883.730 699.040 946.150 ;
        RECT 698.440 883.590 699.040 883.730 ;
        RECT 698.440 883.050 698.580 883.590 ;
        RECT 697.980 882.910 698.580 883.050 ;
        RECT 697.980 835.450 698.120 882.910 ;
        RECT 697.520 835.310 698.120 835.450 ;
        RECT 697.520 16.990 697.660 835.310 ;
        RECT 680.440 16.670 680.700 16.990 ;
        RECT 697.460 16.670 697.720 16.990 ;
        RECT 680.500 2.400 680.640 16.670 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1049.330 946.460 1049.650 946.520 ;
        RECT 1055.310 946.460 1055.630 946.520 ;
        RECT 1049.330 946.320 1055.630 946.460 ;
        RECT 1049.330 946.260 1049.650 946.320 ;
        RECT 1055.310 946.260 1055.630 946.320 ;
        RECT 1055.770 17.580 1056.090 17.640 ;
        RECT 1179.970 17.580 1180.290 17.640 ;
        RECT 1055.770 17.440 1180.290 17.580 ;
        RECT 1055.770 17.380 1056.090 17.440 ;
        RECT 1179.970 17.380 1180.290 17.440 ;
      LAYER via ;
        RECT 1049.360 946.260 1049.620 946.520 ;
        RECT 1055.340 946.260 1055.600 946.520 ;
        RECT 1055.800 17.380 1056.060 17.640 ;
        RECT 1180.000 17.380 1180.260 17.640 ;
      LAYER met2 ;
        RECT 1049.250 960.500 1049.530 964.000 ;
        RECT 1049.250 960.000 1049.560 960.500 ;
        RECT 1049.420 946.550 1049.560 960.000 ;
        RECT 1049.360 946.230 1049.620 946.550 ;
        RECT 1055.340 946.230 1055.600 946.550 ;
        RECT 1055.400 18.090 1055.540 946.230 ;
        RECT 1055.400 17.950 1056.000 18.090 ;
        RECT 1055.860 17.670 1056.000 17.950 ;
        RECT 1055.800 17.350 1056.060 17.670 ;
        RECT 1180.000 17.350 1180.260 17.670 ;
        RECT 1180.060 2.400 1180.200 17.350 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1062.210 17.240 1062.530 17.300 ;
        RECT 1197.910 17.240 1198.230 17.300 ;
        RECT 1062.210 17.100 1198.230 17.240 ;
        RECT 1062.210 17.040 1062.530 17.100 ;
        RECT 1197.910 17.040 1198.230 17.100 ;
      LAYER via ;
        RECT 1062.240 17.040 1062.500 17.300 ;
        RECT 1197.940 17.040 1198.200 17.300 ;
      LAYER met2 ;
        RECT 1061.670 960.570 1061.950 964.000 ;
        RECT 1061.670 960.430 1062.440 960.570 ;
        RECT 1061.670 960.000 1061.950 960.430 ;
        RECT 1062.300 17.330 1062.440 960.430 ;
        RECT 1062.240 17.010 1062.500 17.330 ;
        RECT 1197.940 17.010 1198.200 17.330 ;
        RECT 1198.000 2.400 1198.140 17.010 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1075.550 162.080 1075.870 162.140 ;
        RECT 1214.470 162.080 1214.790 162.140 ;
        RECT 1075.550 161.940 1214.790 162.080 ;
        RECT 1075.550 161.880 1075.870 161.940 ;
        RECT 1214.470 161.880 1214.790 161.940 ;
      LAYER via ;
        RECT 1075.580 161.880 1075.840 162.140 ;
        RECT 1214.500 161.880 1214.760 162.140 ;
      LAYER met2 ;
        RECT 1074.090 960.570 1074.370 964.000 ;
        RECT 1074.090 960.430 1075.780 960.570 ;
        RECT 1074.090 960.000 1074.370 960.430 ;
        RECT 1075.640 162.170 1075.780 960.430 ;
        RECT 1075.580 161.850 1075.840 162.170 ;
        RECT 1214.500 161.850 1214.760 162.170 ;
        RECT 1214.560 17.410 1214.700 161.850 ;
        RECT 1214.560 17.270 1216.080 17.410 ;
        RECT 1215.940 2.400 1216.080 17.270 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1089.810 168.880 1090.130 168.940 ;
        RECT 1228.270 168.880 1228.590 168.940 ;
        RECT 1089.810 168.740 1228.590 168.880 ;
        RECT 1089.810 168.680 1090.130 168.740 ;
        RECT 1228.270 168.680 1228.590 168.740 ;
      LAYER via ;
        RECT 1089.840 168.680 1090.100 168.940 ;
        RECT 1228.300 168.680 1228.560 168.940 ;
      LAYER met2 ;
        RECT 1086.510 960.570 1086.790 964.000 ;
        RECT 1086.510 960.430 1090.040 960.570 ;
        RECT 1086.510 960.000 1086.790 960.430 ;
        RECT 1089.900 168.970 1090.040 960.430 ;
        RECT 1089.840 168.650 1090.100 168.970 ;
        RECT 1228.300 168.650 1228.560 168.970 ;
        RECT 1228.360 17.410 1228.500 168.650 ;
        RECT 1228.360 17.270 1234.020 17.410 ;
        RECT 1233.880 2.400 1234.020 17.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1099.010 947.140 1099.330 947.200 ;
        RECT 1103.150 947.140 1103.470 947.200 ;
        RECT 1099.010 947.000 1103.470 947.140 ;
        RECT 1099.010 946.940 1099.330 947.000 ;
        RECT 1103.150 946.940 1103.470 947.000 ;
        RECT 1103.150 182.820 1103.470 182.880 ;
        RECT 1248.970 182.820 1249.290 182.880 ;
        RECT 1103.150 182.680 1249.290 182.820 ;
        RECT 1103.150 182.620 1103.470 182.680 ;
        RECT 1248.970 182.620 1249.290 182.680 ;
      LAYER via ;
        RECT 1099.040 946.940 1099.300 947.200 ;
        RECT 1103.180 946.940 1103.440 947.200 ;
        RECT 1103.180 182.620 1103.440 182.880 ;
        RECT 1249.000 182.620 1249.260 182.880 ;
      LAYER met2 ;
        RECT 1098.930 960.500 1099.210 964.000 ;
        RECT 1098.930 960.000 1099.240 960.500 ;
        RECT 1099.100 947.230 1099.240 960.000 ;
        RECT 1099.040 946.910 1099.300 947.230 ;
        RECT 1103.180 946.910 1103.440 947.230 ;
        RECT 1103.240 182.910 1103.380 946.910 ;
        RECT 1103.180 182.590 1103.440 182.910 ;
        RECT 1249.000 182.590 1249.260 182.910 ;
        RECT 1249.060 17.410 1249.200 182.590 ;
        RECT 1249.060 17.270 1251.960 17.410 ;
        RECT 1251.820 2.400 1251.960 17.270 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.430 947.480 1111.750 947.540 ;
        RECT 1117.410 947.480 1117.730 947.540 ;
        RECT 1111.430 947.340 1117.730 947.480 ;
        RECT 1111.430 947.280 1111.750 947.340 ;
        RECT 1117.410 947.280 1117.730 947.340 ;
        RECT 1117.410 893.420 1117.730 893.480 ;
        RECT 1262.770 893.420 1263.090 893.480 ;
        RECT 1117.410 893.280 1263.090 893.420 ;
        RECT 1117.410 893.220 1117.730 893.280 ;
        RECT 1262.770 893.220 1263.090 893.280 ;
        RECT 1262.770 17.580 1263.090 17.640 ;
        RECT 1269.210 17.580 1269.530 17.640 ;
        RECT 1262.770 17.440 1269.530 17.580 ;
        RECT 1262.770 17.380 1263.090 17.440 ;
        RECT 1269.210 17.380 1269.530 17.440 ;
      LAYER via ;
        RECT 1111.460 947.280 1111.720 947.540 ;
        RECT 1117.440 947.280 1117.700 947.540 ;
        RECT 1117.440 893.220 1117.700 893.480 ;
        RECT 1262.800 893.220 1263.060 893.480 ;
        RECT 1262.800 17.380 1263.060 17.640 ;
        RECT 1269.240 17.380 1269.500 17.640 ;
      LAYER met2 ;
        RECT 1111.350 960.500 1111.630 964.000 ;
        RECT 1111.350 960.000 1111.660 960.500 ;
        RECT 1111.520 947.570 1111.660 960.000 ;
        RECT 1111.460 947.250 1111.720 947.570 ;
        RECT 1117.440 947.250 1117.700 947.570 ;
        RECT 1117.500 893.510 1117.640 947.250 ;
        RECT 1117.440 893.190 1117.700 893.510 ;
        RECT 1262.800 893.190 1263.060 893.510 ;
        RECT 1262.860 17.670 1263.000 893.190 ;
        RECT 1262.800 17.350 1263.060 17.670 ;
        RECT 1269.240 17.350 1269.500 17.670 ;
        RECT 1269.300 2.400 1269.440 17.350 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1123.850 196.760 1124.170 196.820 ;
        RECT 1283.470 196.760 1283.790 196.820 ;
        RECT 1123.850 196.620 1283.790 196.760 ;
        RECT 1123.850 196.560 1124.170 196.620 ;
        RECT 1283.470 196.560 1283.790 196.620 ;
      LAYER via ;
        RECT 1123.880 196.560 1124.140 196.820 ;
        RECT 1283.500 196.560 1283.760 196.820 ;
      LAYER met2 ;
        RECT 1123.310 960.570 1123.590 964.000 ;
        RECT 1123.310 960.430 1124.080 960.570 ;
        RECT 1123.310 960.000 1123.590 960.430 ;
        RECT 1123.940 196.850 1124.080 960.430 ;
        RECT 1123.880 196.530 1124.140 196.850 ;
        RECT 1283.500 196.530 1283.760 196.850 ;
        RECT 1283.560 17.410 1283.700 196.530 ;
        RECT 1283.560 17.270 1287.380 17.410 ;
        RECT 1287.240 2.400 1287.380 17.270 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 203.560 1138.430 203.620 ;
        RECT 1304.170 203.560 1304.490 203.620 ;
        RECT 1138.110 203.420 1304.490 203.560 ;
        RECT 1138.110 203.360 1138.430 203.420 ;
        RECT 1304.170 203.360 1304.490 203.420 ;
      LAYER via ;
        RECT 1138.140 203.360 1138.400 203.620 ;
        RECT 1304.200 203.360 1304.460 203.620 ;
      LAYER met2 ;
        RECT 1135.730 960.570 1136.010 964.000 ;
        RECT 1135.730 960.430 1138.340 960.570 ;
        RECT 1135.730 960.000 1136.010 960.430 ;
        RECT 1138.200 203.650 1138.340 960.430 ;
        RECT 1138.140 203.330 1138.400 203.650 ;
        RECT 1304.200 203.330 1304.460 203.650 ;
        RECT 1304.260 17.410 1304.400 203.330 ;
        RECT 1304.260 17.270 1305.320 17.410 ;
        RECT 1305.180 2.400 1305.320 17.270 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1148.230 948.500 1148.550 948.560 ;
        RECT 1151.910 948.500 1152.230 948.560 ;
        RECT 1148.230 948.360 1152.230 948.500 ;
        RECT 1148.230 948.300 1148.550 948.360 ;
        RECT 1151.910 948.300 1152.230 948.360 ;
        RECT 1151.910 210.360 1152.230 210.420 ;
        RECT 1317.970 210.360 1318.290 210.420 ;
        RECT 1151.910 210.220 1318.290 210.360 ;
        RECT 1151.910 210.160 1152.230 210.220 ;
        RECT 1317.970 210.160 1318.290 210.220 ;
      LAYER via ;
        RECT 1148.260 948.300 1148.520 948.560 ;
        RECT 1151.940 948.300 1152.200 948.560 ;
        RECT 1151.940 210.160 1152.200 210.420 ;
        RECT 1318.000 210.160 1318.260 210.420 ;
      LAYER met2 ;
        RECT 1148.150 960.500 1148.430 964.000 ;
        RECT 1148.150 960.000 1148.460 960.500 ;
        RECT 1148.320 948.590 1148.460 960.000 ;
        RECT 1148.260 948.270 1148.520 948.590 ;
        RECT 1151.940 948.270 1152.200 948.590 ;
        RECT 1152.000 210.450 1152.140 948.270 ;
        RECT 1151.940 210.130 1152.200 210.450 ;
        RECT 1318.000 210.130 1318.260 210.450 ;
        RECT 1318.060 17.410 1318.200 210.130 ;
        RECT 1318.060 17.270 1323.260 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1160.650 945.440 1160.970 945.500 ;
        RECT 1165.250 945.440 1165.570 945.500 ;
        RECT 1160.650 945.300 1165.570 945.440 ;
        RECT 1160.650 945.240 1160.970 945.300 ;
        RECT 1165.250 945.240 1165.570 945.300 ;
        RECT 1165.250 224.300 1165.570 224.360 ;
        RECT 1338.670 224.300 1338.990 224.360 ;
        RECT 1165.250 224.160 1338.990 224.300 ;
        RECT 1165.250 224.100 1165.570 224.160 ;
        RECT 1338.670 224.100 1338.990 224.160 ;
      LAYER via ;
        RECT 1160.680 945.240 1160.940 945.500 ;
        RECT 1165.280 945.240 1165.540 945.500 ;
        RECT 1165.280 224.100 1165.540 224.360 ;
        RECT 1338.700 224.100 1338.960 224.360 ;
      LAYER met2 ;
        RECT 1160.570 960.500 1160.850 964.000 ;
        RECT 1160.570 960.000 1160.880 960.500 ;
        RECT 1160.740 945.530 1160.880 960.000 ;
        RECT 1160.680 945.210 1160.940 945.530 ;
        RECT 1165.280 945.210 1165.540 945.530 ;
        RECT 1165.340 224.390 1165.480 945.210 ;
        RECT 1165.280 224.070 1165.540 224.390 ;
        RECT 1338.700 224.070 1338.960 224.390 ;
        RECT 1338.760 17.410 1338.900 224.070 ;
        RECT 1338.760 17.270 1340.740 17.410 ;
        RECT 1340.600 2.400 1340.740 17.270 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.770 907.360 711.090 907.420 ;
        RECT 713.990 907.360 714.310 907.420 ;
        RECT 710.770 907.220 714.310 907.360 ;
        RECT 710.770 907.160 711.090 907.220 ;
        RECT 713.990 907.160 714.310 907.220 ;
        RECT 698.350 19.620 698.670 19.680 ;
        RECT 710.770 19.620 711.090 19.680 ;
        RECT 698.350 19.480 711.090 19.620 ;
        RECT 698.350 19.420 698.670 19.480 ;
        RECT 710.770 19.420 711.090 19.480 ;
      LAYER via ;
        RECT 710.800 907.160 711.060 907.420 ;
        RECT 714.020 907.160 714.280 907.420 ;
        RECT 698.380 19.420 698.640 19.680 ;
        RECT 710.800 19.420 711.060 19.680 ;
      LAYER met2 ;
        RECT 715.290 960.570 715.570 964.000 ;
        RECT 714.080 960.430 715.570 960.570 ;
        RECT 714.080 907.450 714.220 960.430 ;
        RECT 715.290 960.000 715.570 960.430 ;
        RECT 710.800 907.130 711.060 907.450 ;
        RECT 714.020 907.130 714.280 907.450 ;
        RECT 710.860 19.710 711.000 907.130 ;
        RECT 698.380 19.390 698.640 19.710 ;
        RECT 710.800 19.390 711.060 19.710 ;
        RECT 698.440 2.400 698.580 19.390 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.070 946.460 1173.390 946.520 ;
        RECT 1179.510 946.460 1179.830 946.520 ;
        RECT 1173.070 946.320 1179.830 946.460 ;
        RECT 1173.070 946.260 1173.390 946.320 ;
        RECT 1179.510 946.260 1179.830 946.320 ;
        RECT 1179.510 231.100 1179.830 231.160 ;
        RECT 1352.470 231.100 1352.790 231.160 ;
        RECT 1179.510 230.960 1352.790 231.100 ;
        RECT 1179.510 230.900 1179.830 230.960 ;
        RECT 1352.470 230.900 1352.790 230.960 ;
        RECT 1352.470 17.920 1352.790 17.980 ;
        RECT 1358.450 17.920 1358.770 17.980 ;
        RECT 1352.470 17.780 1358.770 17.920 ;
        RECT 1352.470 17.720 1352.790 17.780 ;
        RECT 1358.450 17.720 1358.770 17.780 ;
      LAYER via ;
        RECT 1173.100 946.260 1173.360 946.520 ;
        RECT 1179.540 946.260 1179.800 946.520 ;
        RECT 1179.540 230.900 1179.800 231.160 ;
        RECT 1352.500 230.900 1352.760 231.160 ;
        RECT 1352.500 17.720 1352.760 17.980 ;
        RECT 1358.480 17.720 1358.740 17.980 ;
      LAYER met2 ;
        RECT 1172.990 960.500 1173.270 964.000 ;
        RECT 1172.990 960.000 1173.300 960.500 ;
        RECT 1173.160 946.550 1173.300 960.000 ;
        RECT 1173.100 946.230 1173.360 946.550 ;
        RECT 1179.540 946.230 1179.800 946.550 ;
        RECT 1179.600 231.190 1179.740 946.230 ;
        RECT 1179.540 230.870 1179.800 231.190 ;
        RECT 1352.500 230.870 1352.760 231.190 ;
        RECT 1352.560 18.010 1352.700 230.870 ;
        RECT 1352.500 17.690 1352.760 18.010 ;
        RECT 1358.480 17.690 1358.740 18.010 ;
        RECT 1358.540 2.400 1358.680 17.690 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 237.900 1186.270 237.960 ;
        RECT 1373.170 237.900 1373.490 237.960 ;
        RECT 1185.950 237.760 1373.490 237.900 ;
        RECT 1185.950 237.700 1186.270 237.760 ;
        RECT 1373.170 237.700 1373.490 237.760 ;
      LAYER via ;
        RECT 1185.980 237.700 1186.240 237.960 ;
        RECT 1373.200 237.700 1373.460 237.960 ;
      LAYER met2 ;
        RECT 1185.410 960.570 1185.690 964.000 ;
        RECT 1185.410 960.430 1186.180 960.570 ;
        RECT 1185.410 960.000 1185.690 960.430 ;
        RECT 1186.040 237.990 1186.180 960.430 ;
        RECT 1185.980 237.670 1186.240 237.990 ;
        RECT 1373.200 237.670 1373.460 237.990 ;
        RECT 1373.260 17.410 1373.400 237.670 ;
        RECT 1373.260 17.270 1376.620 17.410 ;
        RECT 1376.480 2.400 1376.620 17.270 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1199.750 245.040 1200.070 245.100 ;
        RECT 1393.870 245.040 1394.190 245.100 ;
        RECT 1199.750 244.900 1394.190 245.040 ;
        RECT 1199.750 244.840 1200.070 244.900 ;
        RECT 1393.870 244.840 1394.190 244.900 ;
      LAYER via ;
        RECT 1199.780 244.840 1200.040 245.100 ;
        RECT 1393.900 244.840 1394.160 245.100 ;
      LAYER met2 ;
        RECT 1197.830 960.570 1198.110 964.000 ;
        RECT 1197.830 960.430 1199.980 960.570 ;
        RECT 1197.830 960.000 1198.110 960.430 ;
        RECT 1199.840 245.130 1199.980 960.430 ;
        RECT 1199.780 244.810 1200.040 245.130 ;
        RECT 1393.900 244.810 1394.160 245.130 ;
        RECT 1393.960 17.410 1394.100 244.810 ;
        RECT 1393.960 17.270 1394.560 17.410 ;
        RECT 1394.420 2.400 1394.560 17.270 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.010 251.840 1214.330 251.900 ;
        RECT 1407.670 251.840 1407.990 251.900 ;
        RECT 1214.010 251.700 1407.990 251.840 ;
        RECT 1214.010 251.640 1214.330 251.700 ;
        RECT 1407.670 251.640 1407.990 251.700 ;
      LAYER via ;
        RECT 1214.040 251.640 1214.300 251.900 ;
        RECT 1407.700 251.640 1407.960 251.900 ;
      LAYER met2 ;
        RECT 1210.250 960.570 1210.530 964.000 ;
        RECT 1210.250 960.430 1214.240 960.570 ;
        RECT 1210.250 960.000 1210.530 960.430 ;
        RECT 1214.100 251.930 1214.240 960.430 ;
        RECT 1214.040 251.610 1214.300 251.930 ;
        RECT 1407.700 251.610 1407.960 251.930 ;
        RECT 1407.760 16.730 1407.900 251.610 ;
        RECT 1407.760 16.590 1412.500 16.730 ;
        RECT 1412.360 2.400 1412.500 16.590 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1222.750 950.540 1223.070 950.600 ;
        RECT 1227.350 950.540 1227.670 950.600 ;
        RECT 1222.750 950.400 1227.670 950.540 ;
        RECT 1222.750 950.340 1223.070 950.400 ;
        RECT 1227.350 950.340 1227.670 950.400 ;
        RECT 1227.350 258.640 1227.670 258.700 ;
        RECT 1428.370 258.640 1428.690 258.700 ;
        RECT 1227.350 258.500 1428.690 258.640 ;
        RECT 1227.350 258.440 1227.670 258.500 ;
        RECT 1428.370 258.440 1428.690 258.500 ;
      LAYER via ;
        RECT 1222.780 950.340 1223.040 950.600 ;
        RECT 1227.380 950.340 1227.640 950.600 ;
        RECT 1227.380 258.440 1227.640 258.700 ;
        RECT 1428.400 258.440 1428.660 258.700 ;
      LAYER met2 ;
        RECT 1222.670 960.500 1222.950 964.000 ;
        RECT 1222.670 960.000 1222.980 960.500 ;
        RECT 1222.840 950.630 1222.980 960.000 ;
        RECT 1222.780 950.310 1223.040 950.630 ;
        RECT 1227.380 950.310 1227.640 950.630 ;
        RECT 1227.440 258.730 1227.580 950.310 ;
        RECT 1227.380 258.410 1227.640 258.730 ;
        RECT 1428.400 258.410 1428.660 258.730 ;
        RECT 1428.460 16.730 1428.600 258.410 ;
        RECT 1428.460 16.590 1429.980 16.730 ;
        RECT 1429.840 2.400 1429.980 16.590 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.250 265.440 1234.570 265.500 ;
        RECT 1442.170 265.440 1442.490 265.500 ;
        RECT 1234.250 265.300 1442.490 265.440 ;
        RECT 1234.250 265.240 1234.570 265.300 ;
        RECT 1442.170 265.240 1442.490 265.300 ;
      LAYER via ;
        RECT 1234.280 265.240 1234.540 265.500 ;
        RECT 1442.200 265.240 1442.460 265.500 ;
      LAYER met2 ;
        RECT 1234.630 960.570 1234.910 964.000 ;
        RECT 1234.340 960.430 1234.910 960.570 ;
        RECT 1234.340 265.530 1234.480 960.430 ;
        RECT 1234.630 960.000 1234.910 960.430 ;
        RECT 1234.280 265.210 1234.540 265.530 ;
        RECT 1442.200 265.210 1442.460 265.530 ;
        RECT 1442.260 17.410 1442.400 265.210 ;
        RECT 1442.260 17.270 1447.920 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.050 272.580 1248.370 272.640 ;
        RECT 1462.870 272.580 1463.190 272.640 ;
        RECT 1248.050 272.440 1463.190 272.580 ;
        RECT 1248.050 272.380 1248.370 272.440 ;
        RECT 1462.870 272.380 1463.190 272.440 ;
      LAYER via ;
        RECT 1248.080 272.380 1248.340 272.640 ;
        RECT 1462.900 272.380 1463.160 272.640 ;
      LAYER met2 ;
        RECT 1247.050 960.570 1247.330 964.000 ;
        RECT 1247.050 960.430 1248.280 960.570 ;
        RECT 1247.050 960.000 1247.330 960.430 ;
        RECT 1248.140 272.670 1248.280 960.430 ;
        RECT 1248.080 272.350 1248.340 272.670 ;
        RECT 1462.900 272.350 1463.160 272.670 ;
        RECT 1462.960 17.410 1463.100 272.350 ;
        RECT 1462.960 17.270 1465.860 17.410 ;
        RECT 1465.720 2.400 1465.860 17.270 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 279.380 1262.630 279.440 ;
        RECT 1484.030 279.380 1484.350 279.440 ;
        RECT 1262.310 279.240 1484.350 279.380 ;
        RECT 1262.310 279.180 1262.630 279.240 ;
        RECT 1484.030 279.180 1484.350 279.240 ;
      LAYER via ;
        RECT 1262.340 279.180 1262.600 279.440 ;
        RECT 1484.060 279.180 1484.320 279.440 ;
      LAYER met2 ;
        RECT 1259.470 960.570 1259.750 964.000 ;
        RECT 1259.470 960.430 1262.540 960.570 ;
        RECT 1259.470 960.000 1259.750 960.430 ;
        RECT 1262.400 279.470 1262.540 960.430 ;
        RECT 1262.340 279.150 1262.600 279.470 ;
        RECT 1484.060 279.150 1484.320 279.470 ;
        RECT 1484.120 7.210 1484.260 279.150 ;
        RECT 1483.660 7.070 1484.260 7.210 ;
        RECT 1483.660 2.400 1483.800 7.070 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1275.650 286.180 1275.970 286.240 ;
        RECT 1497.370 286.180 1497.690 286.240 ;
        RECT 1275.650 286.040 1497.690 286.180 ;
        RECT 1275.650 285.980 1275.970 286.040 ;
        RECT 1497.370 285.980 1497.690 286.040 ;
      LAYER via ;
        RECT 1275.680 285.980 1275.940 286.240 ;
        RECT 1497.400 285.980 1497.660 286.240 ;
      LAYER met2 ;
        RECT 1271.890 960.570 1272.170 964.000 ;
        RECT 1271.890 960.430 1275.880 960.570 ;
        RECT 1271.890 960.000 1272.170 960.430 ;
        RECT 1275.740 286.270 1275.880 960.430 ;
        RECT 1275.680 285.950 1275.940 286.270 ;
        RECT 1497.400 285.950 1497.660 286.270 ;
        RECT 1497.460 17.410 1497.600 285.950 ;
        RECT 1497.460 17.270 1501.740 17.410 ;
        RECT 1501.600 2.400 1501.740 17.270 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1284.390 945.440 1284.710 945.500 ;
        RECT 1289.910 945.440 1290.230 945.500 ;
        RECT 1284.390 945.300 1290.230 945.440 ;
        RECT 1284.390 945.240 1284.710 945.300 ;
        RECT 1289.910 945.240 1290.230 945.300 ;
        RECT 1289.910 293.320 1290.230 293.380 ;
        RECT 1518.070 293.320 1518.390 293.380 ;
        RECT 1289.910 293.180 1518.390 293.320 ;
        RECT 1289.910 293.120 1290.230 293.180 ;
        RECT 1518.070 293.120 1518.390 293.180 ;
      LAYER via ;
        RECT 1284.420 945.240 1284.680 945.500 ;
        RECT 1289.940 945.240 1290.200 945.500 ;
        RECT 1289.940 293.120 1290.200 293.380 ;
        RECT 1518.100 293.120 1518.360 293.380 ;
      LAYER met2 ;
        RECT 1284.310 960.500 1284.590 964.000 ;
        RECT 1284.310 960.000 1284.620 960.500 ;
        RECT 1284.480 945.530 1284.620 960.000 ;
        RECT 1284.420 945.210 1284.680 945.530 ;
        RECT 1289.940 945.210 1290.200 945.530 ;
        RECT 1290.000 293.410 1290.140 945.210 ;
        RECT 1289.940 293.090 1290.200 293.410 ;
        RECT 1518.100 293.090 1518.360 293.410 ;
        RECT 1518.160 17.410 1518.300 293.090 ;
        RECT 1518.160 17.270 1519.220 17.410 ;
        RECT 1519.080 2.400 1519.220 17.270 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 716.290 18.940 716.610 19.000 ;
        RECT 724.570 18.940 724.890 19.000 ;
        RECT 716.290 18.800 724.890 18.940 ;
        RECT 716.290 18.740 716.610 18.800 ;
        RECT 724.570 18.740 724.890 18.800 ;
      LAYER via ;
        RECT 716.320 18.740 716.580 19.000 ;
        RECT 724.600 18.740 724.860 19.000 ;
      LAYER met2 ;
        RECT 727.710 960.570 727.990 964.000 ;
        RECT 724.660 960.430 727.990 960.570 ;
        RECT 724.660 19.030 724.800 960.430 ;
        RECT 727.710 960.000 727.990 960.430 ;
        RECT 716.320 18.710 716.580 19.030 ;
        RECT 724.600 18.710 724.860 19.030 ;
        RECT 716.380 2.400 716.520 18.710 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 141.680 1297.130 141.740 ;
        RECT 1531.870 141.680 1532.190 141.740 ;
        RECT 1296.810 141.540 1532.190 141.680 ;
        RECT 1296.810 141.480 1297.130 141.540 ;
        RECT 1531.870 141.480 1532.190 141.540 ;
      LAYER via ;
        RECT 1296.840 141.480 1297.100 141.740 ;
        RECT 1531.900 141.480 1532.160 141.740 ;
      LAYER met2 ;
        RECT 1296.730 960.500 1297.010 964.000 ;
        RECT 1296.730 960.000 1297.040 960.500 ;
        RECT 1296.900 141.770 1297.040 960.000 ;
        RECT 1296.840 141.450 1297.100 141.770 ;
        RECT 1531.900 141.450 1532.160 141.770 ;
        RECT 1531.960 16.730 1532.100 141.450 ;
        RECT 1531.960 16.590 1537.160 16.730 ;
        RECT 1537.020 2.400 1537.160 16.590 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.150 306.920 1310.470 306.980 ;
        RECT 1552.570 306.920 1552.890 306.980 ;
        RECT 1310.150 306.780 1552.890 306.920 ;
        RECT 1310.150 306.720 1310.470 306.780 ;
        RECT 1552.570 306.720 1552.890 306.780 ;
      LAYER via ;
        RECT 1310.180 306.720 1310.440 306.980 ;
        RECT 1552.600 306.720 1552.860 306.980 ;
      LAYER met2 ;
        RECT 1309.150 960.570 1309.430 964.000 ;
        RECT 1309.150 960.430 1310.380 960.570 ;
        RECT 1309.150 960.000 1309.430 960.430 ;
        RECT 1310.240 307.010 1310.380 960.430 ;
        RECT 1310.180 306.690 1310.440 307.010 ;
        RECT 1552.600 306.690 1552.860 307.010 ;
        RECT 1552.660 16.730 1552.800 306.690 ;
        RECT 1552.660 16.590 1555.100 16.730 ;
        RECT 1554.960 2.400 1555.100 16.590 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 320.860 1324.730 320.920 ;
        RECT 1566.370 320.860 1566.690 320.920 ;
        RECT 1324.410 320.720 1566.690 320.860 ;
        RECT 1324.410 320.660 1324.730 320.720 ;
        RECT 1566.370 320.660 1566.690 320.720 ;
        RECT 1566.370 17.580 1566.690 17.640 ;
        RECT 1572.810 17.580 1573.130 17.640 ;
        RECT 1566.370 17.440 1573.130 17.580 ;
        RECT 1566.370 17.380 1566.690 17.440 ;
        RECT 1572.810 17.380 1573.130 17.440 ;
      LAYER via ;
        RECT 1324.440 320.660 1324.700 320.920 ;
        RECT 1566.400 320.660 1566.660 320.920 ;
        RECT 1566.400 17.380 1566.660 17.640 ;
        RECT 1572.840 17.380 1573.100 17.640 ;
      LAYER met2 ;
        RECT 1321.570 960.570 1321.850 964.000 ;
        RECT 1321.570 960.430 1324.640 960.570 ;
        RECT 1321.570 960.000 1321.850 960.430 ;
        RECT 1324.500 320.950 1324.640 960.430 ;
        RECT 1324.440 320.630 1324.700 320.950 ;
        RECT 1566.400 320.630 1566.660 320.950 ;
        RECT 1566.460 17.670 1566.600 320.630 ;
        RECT 1566.400 17.350 1566.660 17.670 ;
        RECT 1572.840 17.350 1573.100 17.670 ;
        RECT 1572.900 2.400 1573.040 17.350 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1334.070 945.440 1334.390 945.500 ;
        RECT 1337.750 945.440 1338.070 945.500 ;
        RECT 1334.070 945.300 1338.070 945.440 ;
        RECT 1334.070 945.240 1334.390 945.300 ;
        RECT 1337.750 945.240 1338.070 945.300 ;
        RECT 1337.750 327.660 1338.070 327.720 ;
        RECT 1587.070 327.660 1587.390 327.720 ;
        RECT 1337.750 327.520 1587.390 327.660 ;
        RECT 1337.750 327.460 1338.070 327.520 ;
        RECT 1587.070 327.460 1587.390 327.520 ;
      LAYER via ;
        RECT 1334.100 945.240 1334.360 945.500 ;
        RECT 1337.780 945.240 1338.040 945.500 ;
        RECT 1337.780 327.460 1338.040 327.720 ;
        RECT 1587.100 327.460 1587.360 327.720 ;
      LAYER met2 ;
        RECT 1333.990 960.500 1334.270 964.000 ;
        RECT 1333.990 960.000 1334.300 960.500 ;
        RECT 1334.160 945.530 1334.300 960.000 ;
        RECT 1334.100 945.210 1334.360 945.530 ;
        RECT 1337.780 945.210 1338.040 945.530 ;
        RECT 1337.840 327.750 1337.980 945.210 ;
        RECT 1337.780 327.430 1338.040 327.750 ;
        RECT 1587.100 327.430 1587.360 327.750 ;
        RECT 1587.160 17.410 1587.300 327.430 ;
        RECT 1587.160 17.270 1590.520 17.410 ;
        RECT 1590.380 2.400 1590.520 17.270 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 949.860 1346.350 949.920 ;
        RECT 1351.550 949.860 1351.870 949.920 ;
        RECT 1346.030 949.720 1351.870 949.860 ;
        RECT 1346.030 949.660 1346.350 949.720 ;
        RECT 1351.550 949.660 1351.870 949.720 ;
        RECT 1351.550 334.460 1351.870 334.520 ;
        RECT 1607.770 334.460 1608.090 334.520 ;
        RECT 1351.550 334.320 1608.090 334.460 ;
        RECT 1351.550 334.260 1351.870 334.320 ;
        RECT 1607.770 334.260 1608.090 334.320 ;
      LAYER via ;
        RECT 1346.060 949.660 1346.320 949.920 ;
        RECT 1351.580 949.660 1351.840 949.920 ;
        RECT 1351.580 334.260 1351.840 334.520 ;
        RECT 1607.800 334.260 1608.060 334.520 ;
      LAYER met2 ;
        RECT 1345.950 960.500 1346.230 964.000 ;
        RECT 1345.950 960.000 1346.260 960.500 ;
        RECT 1346.120 949.950 1346.260 960.000 ;
        RECT 1346.060 949.630 1346.320 949.950 ;
        RECT 1351.580 949.630 1351.840 949.950 ;
        RECT 1351.640 334.550 1351.780 949.630 ;
        RECT 1351.580 334.230 1351.840 334.550 ;
        RECT 1607.800 334.230 1608.060 334.550 ;
        RECT 1607.860 17.410 1608.000 334.230 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.910 341.600 1359.230 341.660 ;
        RECT 1621.570 341.600 1621.890 341.660 ;
        RECT 1358.910 341.460 1621.890 341.600 ;
        RECT 1358.910 341.400 1359.230 341.460 ;
        RECT 1621.570 341.400 1621.890 341.460 ;
      LAYER via ;
        RECT 1358.940 341.400 1359.200 341.660 ;
        RECT 1621.600 341.400 1621.860 341.660 ;
      LAYER met2 ;
        RECT 1358.370 960.570 1358.650 964.000 ;
        RECT 1358.370 960.430 1359.140 960.570 ;
        RECT 1358.370 960.000 1358.650 960.430 ;
        RECT 1359.000 341.690 1359.140 960.430 ;
        RECT 1358.940 341.370 1359.200 341.690 ;
        RECT 1621.600 341.370 1621.860 341.690 ;
        RECT 1621.660 17.410 1621.800 341.370 ;
        RECT 1621.660 17.270 1626.400 17.410 ;
        RECT 1626.260 2.400 1626.400 17.270 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.250 348.400 1372.570 348.460 ;
        RECT 1642.270 348.400 1642.590 348.460 ;
        RECT 1372.250 348.260 1642.590 348.400 ;
        RECT 1372.250 348.200 1372.570 348.260 ;
        RECT 1642.270 348.200 1642.590 348.260 ;
      LAYER via ;
        RECT 1372.280 348.200 1372.540 348.460 ;
        RECT 1642.300 348.200 1642.560 348.460 ;
      LAYER met2 ;
        RECT 1370.790 960.570 1371.070 964.000 ;
        RECT 1370.790 960.430 1372.480 960.570 ;
        RECT 1370.790 960.000 1371.070 960.430 ;
        RECT 1372.340 348.490 1372.480 960.430 ;
        RECT 1372.280 348.170 1372.540 348.490 ;
        RECT 1642.300 348.170 1642.560 348.490 ;
        RECT 1642.360 17.410 1642.500 348.170 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 355.200 1386.830 355.260 ;
        RECT 1656.070 355.200 1656.390 355.260 ;
        RECT 1386.510 355.060 1656.390 355.200 ;
        RECT 1386.510 355.000 1386.830 355.060 ;
        RECT 1656.070 355.000 1656.390 355.060 ;
        RECT 1656.070 17.920 1656.390 17.980 ;
        RECT 1662.050 17.920 1662.370 17.980 ;
        RECT 1656.070 17.780 1662.370 17.920 ;
        RECT 1656.070 17.720 1656.390 17.780 ;
        RECT 1662.050 17.720 1662.370 17.780 ;
      LAYER via ;
        RECT 1386.540 355.000 1386.800 355.260 ;
        RECT 1656.100 355.000 1656.360 355.260 ;
        RECT 1656.100 17.720 1656.360 17.980 ;
        RECT 1662.080 17.720 1662.340 17.980 ;
      LAYER met2 ;
        RECT 1383.210 960.570 1383.490 964.000 ;
        RECT 1383.210 960.430 1386.740 960.570 ;
        RECT 1383.210 960.000 1383.490 960.430 ;
        RECT 1386.600 355.290 1386.740 960.430 ;
        RECT 1386.540 354.970 1386.800 355.290 ;
        RECT 1656.100 354.970 1656.360 355.290 ;
        RECT 1656.160 18.010 1656.300 354.970 ;
        RECT 1656.100 17.690 1656.360 18.010 ;
        RECT 1662.080 17.690 1662.340 18.010 ;
        RECT 1662.140 2.400 1662.280 17.690 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 945.440 1396.030 945.500 ;
        RECT 1399.850 945.440 1400.170 945.500 ;
        RECT 1395.710 945.300 1400.170 945.440 ;
        RECT 1395.710 945.240 1396.030 945.300 ;
        RECT 1399.850 945.240 1400.170 945.300 ;
        RECT 1399.850 369.140 1400.170 369.200 ;
        RECT 1676.770 369.140 1677.090 369.200 ;
        RECT 1399.850 369.000 1677.090 369.140 ;
        RECT 1399.850 368.940 1400.170 369.000 ;
        RECT 1676.770 368.940 1677.090 369.000 ;
      LAYER via ;
        RECT 1395.740 945.240 1396.000 945.500 ;
        RECT 1399.880 945.240 1400.140 945.500 ;
        RECT 1399.880 368.940 1400.140 369.200 ;
        RECT 1676.800 368.940 1677.060 369.200 ;
      LAYER met2 ;
        RECT 1395.630 960.500 1395.910 964.000 ;
        RECT 1395.630 960.000 1395.940 960.500 ;
        RECT 1395.800 945.530 1395.940 960.000 ;
        RECT 1395.740 945.210 1396.000 945.530 ;
        RECT 1399.880 945.210 1400.140 945.530 ;
        RECT 1399.940 369.230 1400.080 945.210 ;
        RECT 1399.880 368.910 1400.140 369.230 ;
        RECT 1676.800 368.910 1677.060 369.230 ;
        RECT 1676.860 17.410 1677.000 368.910 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1408.130 950.880 1408.450 950.940 ;
        RECT 1413.650 950.880 1413.970 950.940 ;
        RECT 1408.130 950.740 1413.970 950.880 ;
        RECT 1408.130 950.680 1408.450 950.740 ;
        RECT 1413.650 950.680 1413.970 950.740 ;
        RECT 1413.650 362.340 1413.970 362.400 ;
        RECT 1697.470 362.340 1697.790 362.400 ;
        RECT 1413.650 362.200 1697.790 362.340 ;
        RECT 1413.650 362.140 1413.970 362.200 ;
        RECT 1697.470 362.140 1697.790 362.200 ;
      LAYER via ;
        RECT 1408.160 950.680 1408.420 950.940 ;
        RECT 1413.680 950.680 1413.940 950.940 ;
        RECT 1413.680 362.140 1413.940 362.400 ;
        RECT 1697.500 362.140 1697.760 362.400 ;
      LAYER met2 ;
        RECT 1408.050 960.500 1408.330 964.000 ;
        RECT 1408.050 960.000 1408.360 960.500 ;
        RECT 1408.220 950.970 1408.360 960.000 ;
        RECT 1408.160 950.650 1408.420 950.970 ;
        RECT 1413.680 950.650 1413.940 950.970 ;
        RECT 1413.740 362.430 1413.880 950.650 ;
        RECT 1413.680 362.110 1413.940 362.430 ;
        RECT 1697.500 362.110 1697.760 362.430 ;
        RECT 1697.560 2.400 1697.700 362.110 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.230 17.920 734.550 17.980 ;
        RECT 738.830 17.920 739.150 17.980 ;
        RECT 734.230 17.780 739.150 17.920 ;
        RECT 734.230 17.720 734.550 17.780 ;
        RECT 738.830 17.720 739.150 17.780 ;
      LAYER via ;
        RECT 734.260 17.720 734.520 17.980 ;
        RECT 738.860 17.720 739.120 17.980 ;
      LAYER met2 ;
        RECT 740.130 960.570 740.410 964.000 ;
        RECT 738.920 960.430 740.410 960.570 ;
        RECT 738.920 18.010 739.060 960.430 ;
        RECT 740.130 960.000 740.410 960.430 ;
        RECT 734.260 17.690 734.520 18.010 ;
        RECT 738.860 17.690 739.120 18.010 ;
        RECT 734.320 2.400 734.460 17.690 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1420.550 375.940 1420.870 376.000 ;
        RECT 1711.270 375.940 1711.590 376.000 ;
        RECT 1420.550 375.800 1711.590 375.940 ;
        RECT 1420.550 375.740 1420.870 375.800 ;
        RECT 1711.270 375.740 1711.590 375.800 ;
      LAYER via ;
        RECT 1420.580 375.740 1420.840 376.000 ;
        RECT 1711.300 375.740 1711.560 376.000 ;
      LAYER met2 ;
        RECT 1420.470 960.500 1420.750 964.000 ;
        RECT 1420.470 960.000 1420.780 960.500 ;
        RECT 1420.640 376.030 1420.780 960.000 ;
        RECT 1420.580 375.710 1420.840 376.030 ;
        RECT 1711.300 375.710 1711.560 376.030 ;
        RECT 1711.360 17.410 1711.500 375.710 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.350 382.740 1434.670 382.800 ;
        RECT 1731.970 382.740 1732.290 382.800 ;
        RECT 1434.350 382.600 1732.290 382.740 ;
        RECT 1434.350 382.540 1434.670 382.600 ;
        RECT 1731.970 382.540 1732.290 382.600 ;
      LAYER via ;
        RECT 1434.380 382.540 1434.640 382.800 ;
        RECT 1732.000 382.540 1732.260 382.800 ;
      LAYER met2 ;
        RECT 1432.890 960.570 1433.170 964.000 ;
        RECT 1432.890 960.430 1434.580 960.570 ;
        RECT 1432.890 960.000 1433.170 960.430 ;
        RECT 1434.440 382.830 1434.580 960.430 ;
        RECT 1434.380 382.510 1434.640 382.830 ;
        RECT 1732.000 382.510 1732.260 382.830 ;
        RECT 1732.060 17.410 1732.200 382.510 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 389.880 1448.930 389.940 ;
        RECT 1745.770 389.880 1746.090 389.940 ;
        RECT 1448.610 389.740 1746.090 389.880 ;
        RECT 1448.610 389.680 1448.930 389.740 ;
        RECT 1745.770 389.680 1746.090 389.740 ;
      LAYER via ;
        RECT 1448.640 389.680 1448.900 389.940 ;
        RECT 1745.800 389.680 1746.060 389.940 ;
      LAYER met2 ;
        RECT 1445.310 960.570 1445.590 964.000 ;
        RECT 1445.310 960.430 1448.840 960.570 ;
        RECT 1445.310 960.000 1445.590 960.430 ;
        RECT 1448.700 389.970 1448.840 960.430 ;
        RECT 1448.640 389.650 1448.900 389.970 ;
        RECT 1745.800 389.650 1746.060 389.970 ;
        RECT 1745.860 17.410 1746.000 389.650 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1457.810 945.440 1458.130 945.500 ;
        RECT 1461.950 945.440 1462.270 945.500 ;
        RECT 1457.810 945.300 1462.270 945.440 ;
        RECT 1457.810 945.240 1458.130 945.300 ;
        RECT 1461.950 945.240 1462.270 945.300 ;
        RECT 1461.950 396.680 1462.270 396.740 ;
        RECT 1766.470 396.680 1766.790 396.740 ;
        RECT 1461.950 396.540 1766.790 396.680 ;
        RECT 1461.950 396.480 1462.270 396.540 ;
        RECT 1766.470 396.480 1766.790 396.540 ;
      LAYER via ;
        RECT 1457.840 945.240 1458.100 945.500 ;
        RECT 1461.980 945.240 1462.240 945.500 ;
        RECT 1461.980 396.480 1462.240 396.740 ;
        RECT 1766.500 396.480 1766.760 396.740 ;
      LAYER met2 ;
        RECT 1457.730 960.500 1458.010 964.000 ;
        RECT 1457.730 960.000 1458.040 960.500 ;
        RECT 1457.900 945.530 1458.040 960.000 ;
        RECT 1457.840 945.210 1458.100 945.530 ;
        RECT 1461.980 945.210 1462.240 945.530 ;
        RECT 1462.040 396.770 1462.180 945.210 ;
        RECT 1461.980 396.450 1462.240 396.770 ;
        RECT 1766.500 396.450 1766.760 396.770 ;
        RECT 1766.560 17.410 1766.700 396.450 ;
        RECT 1766.560 17.270 1769.000 17.410 ;
        RECT 1768.860 2.400 1769.000 17.270 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.770 947.140 1470.090 947.200 ;
        RECT 1476.210 947.140 1476.530 947.200 ;
        RECT 1469.770 947.000 1476.530 947.140 ;
        RECT 1469.770 946.940 1470.090 947.000 ;
        RECT 1476.210 946.940 1476.530 947.000 ;
        RECT 1476.210 403.480 1476.530 403.540 ;
        RECT 1780.270 403.480 1780.590 403.540 ;
        RECT 1476.210 403.340 1780.590 403.480 ;
        RECT 1476.210 403.280 1476.530 403.340 ;
        RECT 1780.270 403.280 1780.590 403.340 ;
        RECT 1780.270 17.580 1780.590 17.640 ;
        RECT 1786.710 17.580 1787.030 17.640 ;
        RECT 1780.270 17.440 1787.030 17.580 ;
        RECT 1780.270 17.380 1780.590 17.440 ;
        RECT 1786.710 17.380 1787.030 17.440 ;
      LAYER via ;
        RECT 1469.800 946.940 1470.060 947.200 ;
        RECT 1476.240 946.940 1476.500 947.200 ;
        RECT 1476.240 403.280 1476.500 403.540 ;
        RECT 1780.300 403.280 1780.560 403.540 ;
        RECT 1780.300 17.380 1780.560 17.640 ;
        RECT 1786.740 17.380 1787.000 17.640 ;
      LAYER met2 ;
        RECT 1469.690 960.500 1469.970 964.000 ;
        RECT 1469.690 960.000 1470.000 960.500 ;
        RECT 1469.860 947.230 1470.000 960.000 ;
        RECT 1469.800 946.910 1470.060 947.230 ;
        RECT 1476.240 946.910 1476.500 947.230 ;
        RECT 1476.300 403.570 1476.440 946.910 ;
        RECT 1476.240 403.250 1476.500 403.570 ;
        RECT 1780.300 403.250 1780.560 403.570 ;
        RECT 1780.360 17.670 1780.500 403.250 ;
        RECT 1780.300 17.350 1780.560 17.670 ;
        RECT 1786.740 17.350 1787.000 17.670 ;
        RECT 1786.800 2.400 1786.940 17.350 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1482.650 196.760 1482.970 196.820 ;
        RECT 1800.970 196.760 1801.290 196.820 ;
        RECT 1482.650 196.620 1801.290 196.760 ;
        RECT 1482.650 196.560 1482.970 196.620 ;
        RECT 1800.970 196.560 1801.290 196.620 ;
      LAYER via ;
        RECT 1482.680 196.560 1482.940 196.820 ;
        RECT 1801.000 196.560 1801.260 196.820 ;
      LAYER met2 ;
        RECT 1482.110 960.570 1482.390 964.000 ;
        RECT 1482.110 960.430 1482.880 960.570 ;
        RECT 1482.110 960.000 1482.390 960.430 ;
        RECT 1482.740 196.850 1482.880 960.430 ;
        RECT 1482.680 196.530 1482.940 196.850 ;
        RECT 1801.000 196.530 1801.260 196.850 ;
        RECT 1801.060 16.730 1801.200 196.530 ;
        RECT 1801.060 16.590 1804.880 16.730 ;
        RECT 1804.740 2.400 1804.880 16.590 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.450 410.620 1496.770 410.680 ;
        RECT 1821.670 410.620 1821.990 410.680 ;
        RECT 1496.450 410.480 1821.990 410.620 ;
        RECT 1496.450 410.420 1496.770 410.480 ;
        RECT 1821.670 410.420 1821.990 410.480 ;
        RECT 1821.670 2.960 1821.990 3.020 ;
        RECT 1822.590 2.960 1822.910 3.020 ;
        RECT 1821.670 2.820 1822.910 2.960 ;
        RECT 1821.670 2.760 1821.990 2.820 ;
        RECT 1822.590 2.760 1822.910 2.820 ;
      LAYER via ;
        RECT 1496.480 410.420 1496.740 410.680 ;
        RECT 1821.700 410.420 1821.960 410.680 ;
        RECT 1821.700 2.760 1821.960 3.020 ;
        RECT 1822.620 2.760 1822.880 3.020 ;
      LAYER met2 ;
        RECT 1494.530 960.570 1494.810 964.000 ;
        RECT 1494.530 960.430 1496.680 960.570 ;
        RECT 1494.530 960.000 1494.810 960.430 ;
        RECT 1496.540 410.710 1496.680 960.430 ;
        RECT 1496.480 410.390 1496.740 410.710 ;
        RECT 1821.700 410.390 1821.960 410.710 ;
        RECT 1821.760 3.050 1821.900 410.390 ;
        RECT 1821.700 2.730 1821.960 3.050 ;
        RECT 1822.620 2.730 1822.880 3.050 ;
        RECT 1822.680 2.400 1822.820 2.730 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.030 945.440 1507.350 945.500 ;
        RECT 1510.710 945.440 1511.030 945.500 ;
        RECT 1507.030 945.300 1511.030 945.440 ;
        RECT 1507.030 945.240 1507.350 945.300 ;
        RECT 1510.710 945.240 1511.030 945.300 ;
        RECT 1510.710 417.420 1511.030 417.480 ;
        RECT 1835.470 417.420 1835.790 417.480 ;
        RECT 1510.710 417.280 1835.790 417.420 ;
        RECT 1510.710 417.220 1511.030 417.280 ;
        RECT 1835.470 417.220 1835.790 417.280 ;
        RECT 1835.470 2.960 1835.790 3.020 ;
        RECT 1840.070 2.960 1840.390 3.020 ;
        RECT 1835.470 2.820 1840.390 2.960 ;
        RECT 1835.470 2.760 1835.790 2.820 ;
        RECT 1840.070 2.760 1840.390 2.820 ;
      LAYER via ;
        RECT 1507.060 945.240 1507.320 945.500 ;
        RECT 1510.740 945.240 1511.000 945.500 ;
        RECT 1510.740 417.220 1511.000 417.480 ;
        RECT 1835.500 417.220 1835.760 417.480 ;
        RECT 1835.500 2.760 1835.760 3.020 ;
        RECT 1840.100 2.760 1840.360 3.020 ;
      LAYER met2 ;
        RECT 1506.950 960.500 1507.230 964.000 ;
        RECT 1506.950 960.000 1507.260 960.500 ;
        RECT 1507.120 945.530 1507.260 960.000 ;
        RECT 1507.060 945.210 1507.320 945.530 ;
        RECT 1510.740 945.210 1511.000 945.530 ;
        RECT 1510.800 417.510 1510.940 945.210 ;
        RECT 1510.740 417.190 1511.000 417.510 ;
        RECT 1835.500 417.190 1835.760 417.510 ;
        RECT 1835.560 3.050 1835.700 417.190 ;
        RECT 1835.500 2.730 1835.760 3.050 ;
        RECT 1840.100 2.730 1840.360 3.050 ;
        RECT 1840.160 2.400 1840.300 2.730 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1519.450 951.900 1519.770 951.960 ;
        RECT 1524.050 951.900 1524.370 951.960 ;
        RECT 1519.450 951.760 1524.370 951.900 ;
        RECT 1519.450 951.700 1519.770 951.760 ;
        RECT 1524.050 951.700 1524.370 951.760 ;
        RECT 1524.050 431.360 1524.370 431.420 ;
        RECT 1856.170 431.360 1856.490 431.420 ;
        RECT 1524.050 431.220 1856.490 431.360 ;
        RECT 1524.050 431.160 1524.370 431.220 ;
        RECT 1856.170 431.160 1856.490 431.220 ;
      LAYER via ;
        RECT 1519.480 951.700 1519.740 951.960 ;
        RECT 1524.080 951.700 1524.340 951.960 ;
        RECT 1524.080 431.160 1524.340 431.420 ;
        RECT 1856.200 431.160 1856.460 431.420 ;
      LAYER met2 ;
        RECT 1519.370 960.500 1519.650 964.000 ;
        RECT 1519.370 960.000 1519.680 960.500 ;
        RECT 1519.540 951.990 1519.680 960.000 ;
        RECT 1519.480 951.670 1519.740 951.990 ;
        RECT 1524.080 951.670 1524.340 951.990 ;
        RECT 1524.140 431.450 1524.280 951.670 ;
        RECT 1524.080 431.130 1524.340 431.450 ;
        RECT 1856.200 431.130 1856.460 431.450 ;
        RECT 1856.260 3.130 1856.400 431.130 ;
        RECT 1856.260 2.990 1858.240 3.130 ;
        RECT 1858.100 2.400 1858.240 2.990 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.870 946.460 1532.190 946.520 ;
        RECT 1538.310 946.460 1538.630 946.520 ;
        RECT 1531.870 946.320 1538.630 946.460 ;
        RECT 1531.870 946.260 1532.190 946.320 ;
        RECT 1538.310 946.260 1538.630 946.320 ;
        RECT 1538.310 424.220 1538.630 424.280 ;
        RECT 1869.970 424.220 1870.290 424.280 ;
        RECT 1538.310 424.080 1870.290 424.220 ;
        RECT 1538.310 424.020 1538.630 424.080 ;
        RECT 1869.970 424.020 1870.290 424.080 ;
        RECT 1869.970 17.920 1870.290 17.980 ;
        RECT 1875.950 17.920 1876.270 17.980 ;
        RECT 1869.970 17.780 1876.270 17.920 ;
        RECT 1869.970 17.720 1870.290 17.780 ;
        RECT 1875.950 17.720 1876.270 17.780 ;
      LAYER via ;
        RECT 1531.900 946.260 1532.160 946.520 ;
        RECT 1538.340 946.260 1538.600 946.520 ;
        RECT 1538.340 424.020 1538.600 424.280 ;
        RECT 1870.000 424.020 1870.260 424.280 ;
        RECT 1870.000 17.720 1870.260 17.980 ;
        RECT 1875.980 17.720 1876.240 17.980 ;
      LAYER met2 ;
        RECT 1531.790 960.500 1532.070 964.000 ;
        RECT 1531.790 960.000 1532.100 960.500 ;
        RECT 1531.960 946.550 1532.100 960.000 ;
        RECT 1531.900 946.230 1532.160 946.550 ;
        RECT 1538.340 946.230 1538.600 946.550 ;
        RECT 1538.400 424.310 1538.540 946.230 ;
        RECT 1538.340 423.990 1538.600 424.310 ;
        RECT 1870.000 423.990 1870.260 424.310 ;
        RECT 1870.060 18.010 1870.200 423.990 ;
        RECT 1870.000 17.690 1870.260 18.010 ;
        RECT 1875.980 17.690 1876.240 18.010 ;
        RECT 1876.040 2.400 1876.180 17.690 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.550 960.500 752.830 964.000 ;
        RECT 752.550 960.000 752.860 960.500 ;
        RECT 752.720 17.410 752.860 960.000 ;
        RECT 752.260 17.270 752.860 17.410 ;
        RECT 752.260 2.400 752.400 17.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 24.040 1545.530 24.100 ;
        RECT 1893.890 24.040 1894.210 24.100 ;
        RECT 1545.210 23.900 1894.210 24.040 ;
        RECT 1545.210 23.840 1545.530 23.900 ;
        RECT 1893.890 23.840 1894.210 23.900 ;
      LAYER via ;
        RECT 1545.240 23.840 1545.500 24.100 ;
        RECT 1893.920 23.840 1894.180 24.100 ;
      LAYER met2 ;
        RECT 1544.210 960.570 1544.490 964.000 ;
        RECT 1544.210 960.430 1545.440 960.570 ;
        RECT 1544.210 960.000 1544.490 960.430 ;
        RECT 1545.300 24.130 1545.440 960.430 ;
        RECT 1545.240 23.810 1545.500 24.130 ;
        RECT 1893.920 23.810 1894.180 24.130 ;
        RECT 1893.980 2.400 1894.120 23.810 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 444.960 1559.330 445.020 ;
        RECT 1911.370 444.960 1911.690 445.020 ;
        RECT 1559.010 444.820 1911.690 444.960 ;
        RECT 1559.010 444.760 1559.330 444.820 ;
        RECT 1911.370 444.760 1911.690 444.820 ;
      LAYER via ;
        RECT 1559.040 444.760 1559.300 445.020 ;
        RECT 1911.400 444.760 1911.660 445.020 ;
      LAYER met2 ;
        RECT 1556.630 960.570 1556.910 964.000 ;
        RECT 1556.630 960.430 1559.240 960.570 ;
        RECT 1556.630 960.000 1556.910 960.430 ;
        RECT 1559.100 445.050 1559.240 960.430 ;
        RECT 1559.040 444.730 1559.300 445.050 ;
        RECT 1911.400 444.730 1911.660 445.050 ;
        RECT 1911.460 7.890 1911.600 444.730 ;
        RECT 1911.460 7.750 1912.060 7.890 ;
        RECT 1911.920 2.400 1912.060 7.750 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.350 458.900 1572.670 458.960 ;
        RECT 1925.170 458.900 1925.490 458.960 ;
        RECT 1572.350 458.760 1925.490 458.900 ;
        RECT 1572.350 458.700 1572.670 458.760 ;
        RECT 1925.170 458.700 1925.490 458.760 ;
      LAYER via ;
        RECT 1572.380 458.700 1572.640 458.960 ;
        RECT 1925.200 458.700 1925.460 458.960 ;
      LAYER met2 ;
        RECT 1569.050 960.570 1569.330 964.000 ;
        RECT 1569.050 960.430 1572.580 960.570 ;
        RECT 1569.050 960.000 1569.330 960.430 ;
        RECT 1572.440 458.990 1572.580 960.430 ;
        RECT 1572.380 458.670 1572.640 458.990 ;
        RECT 1925.200 458.670 1925.460 458.990 ;
        RECT 1925.260 17.410 1925.400 458.670 ;
        RECT 1925.260 17.270 1929.540 17.410 ;
        RECT 1929.400 2.400 1929.540 17.270 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.090 950.540 1581.410 950.600 ;
        RECT 1586.150 950.540 1586.470 950.600 ;
        RECT 1581.090 950.400 1586.470 950.540 ;
        RECT 1581.090 950.340 1581.410 950.400 ;
        RECT 1586.150 950.340 1586.470 950.400 ;
        RECT 1586.150 465.700 1586.470 465.760 ;
        RECT 1945.870 465.700 1946.190 465.760 ;
        RECT 1586.150 465.560 1946.190 465.700 ;
        RECT 1586.150 465.500 1586.470 465.560 ;
        RECT 1945.870 465.500 1946.190 465.560 ;
      LAYER via ;
        RECT 1581.120 950.340 1581.380 950.600 ;
        RECT 1586.180 950.340 1586.440 950.600 ;
        RECT 1586.180 465.500 1586.440 465.760 ;
        RECT 1945.900 465.500 1946.160 465.760 ;
      LAYER met2 ;
        RECT 1581.010 960.500 1581.290 964.000 ;
        RECT 1581.010 960.000 1581.320 960.500 ;
        RECT 1581.180 950.630 1581.320 960.000 ;
        RECT 1581.120 950.310 1581.380 950.630 ;
        RECT 1586.180 950.310 1586.440 950.630 ;
        RECT 1586.240 465.790 1586.380 950.310 ;
        RECT 1586.180 465.470 1586.440 465.790 ;
        RECT 1945.900 465.470 1946.160 465.790 ;
        RECT 1945.960 17.410 1946.100 465.470 ;
        RECT 1945.960 17.270 1947.480 17.410 ;
        RECT 1947.340 2.400 1947.480 17.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 472.500 1593.830 472.560 ;
        RECT 1959.670 472.500 1959.990 472.560 ;
        RECT 1593.510 472.360 1959.990 472.500 ;
        RECT 1593.510 472.300 1593.830 472.360 ;
        RECT 1959.670 472.300 1959.990 472.360 ;
      LAYER via ;
        RECT 1593.540 472.300 1593.800 472.560 ;
        RECT 1959.700 472.300 1959.960 472.560 ;
      LAYER met2 ;
        RECT 1593.430 960.500 1593.710 964.000 ;
        RECT 1593.430 960.000 1593.740 960.500 ;
        RECT 1593.600 472.590 1593.740 960.000 ;
        RECT 1593.540 472.270 1593.800 472.590 ;
        RECT 1959.700 472.270 1959.960 472.590 ;
        RECT 1959.760 17.410 1959.900 472.270 ;
        RECT 1959.760 17.270 1965.420 17.410 ;
        RECT 1965.280 2.400 1965.420 17.270 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1606.850 479.640 1607.170 479.700 ;
        RECT 1980.370 479.640 1980.690 479.700 ;
        RECT 1606.850 479.500 1980.690 479.640 ;
        RECT 1606.850 479.440 1607.170 479.500 ;
        RECT 1980.370 479.440 1980.690 479.500 ;
      LAYER via ;
        RECT 1606.880 479.440 1607.140 479.700 ;
        RECT 1980.400 479.440 1980.660 479.700 ;
      LAYER met2 ;
        RECT 1605.850 960.570 1606.130 964.000 ;
        RECT 1605.850 960.430 1607.080 960.570 ;
        RECT 1605.850 960.000 1606.130 960.430 ;
        RECT 1606.940 479.730 1607.080 960.430 ;
        RECT 1606.880 479.410 1607.140 479.730 ;
        RECT 1980.400 479.410 1980.660 479.730 ;
        RECT 1980.460 17.410 1980.600 479.410 ;
        RECT 1980.460 17.270 1983.360 17.410 ;
        RECT 1983.220 2.400 1983.360 17.270 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1621.110 486.440 1621.430 486.500 ;
        RECT 2001.070 486.440 2001.390 486.500 ;
        RECT 1621.110 486.300 2001.390 486.440 ;
        RECT 1621.110 486.240 1621.430 486.300 ;
        RECT 2001.070 486.240 2001.390 486.300 ;
      LAYER via ;
        RECT 1621.140 486.240 1621.400 486.500 ;
        RECT 2001.100 486.240 2001.360 486.500 ;
      LAYER met2 ;
        RECT 1618.270 960.570 1618.550 964.000 ;
        RECT 1618.270 960.430 1621.340 960.570 ;
        RECT 1618.270 960.000 1618.550 960.430 ;
        RECT 1621.200 486.530 1621.340 960.430 ;
        RECT 1621.140 486.210 1621.400 486.530 ;
        RECT 2001.100 486.210 2001.360 486.530 ;
        RECT 2001.160 2.400 2001.300 486.210 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.450 493.240 1634.770 493.300 ;
        RECT 2014.870 493.240 2015.190 493.300 ;
        RECT 1634.450 493.100 2015.190 493.240 ;
        RECT 1634.450 493.040 1634.770 493.100 ;
        RECT 2014.870 493.040 2015.190 493.100 ;
      LAYER via ;
        RECT 1634.480 493.040 1634.740 493.300 ;
        RECT 2014.900 493.040 2015.160 493.300 ;
      LAYER met2 ;
        RECT 1630.690 960.570 1630.970 964.000 ;
        RECT 1630.690 960.430 1634.680 960.570 ;
        RECT 1630.690 960.000 1630.970 960.430 ;
        RECT 1634.540 493.330 1634.680 960.430 ;
        RECT 1634.480 493.010 1634.740 493.330 ;
        RECT 2014.900 493.010 2015.160 493.330 ;
        RECT 2014.960 17.410 2015.100 493.010 ;
        RECT 2014.960 17.270 2018.780 17.410 ;
        RECT 2018.640 2.400 2018.780 17.270 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1643.190 947.140 1643.510 947.200 ;
        RECT 1648.710 947.140 1649.030 947.200 ;
        RECT 1643.190 947.000 1649.030 947.140 ;
        RECT 1643.190 946.940 1643.510 947.000 ;
        RECT 1648.710 946.940 1649.030 947.000 ;
        RECT 1648.710 500.040 1649.030 500.100 ;
        RECT 2035.570 500.040 2035.890 500.100 ;
        RECT 1648.710 499.900 2035.890 500.040 ;
        RECT 1648.710 499.840 1649.030 499.900 ;
        RECT 2035.570 499.840 2035.890 499.900 ;
      LAYER via ;
        RECT 1643.220 946.940 1643.480 947.200 ;
        RECT 1648.740 946.940 1649.000 947.200 ;
        RECT 1648.740 499.840 1649.000 500.100 ;
        RECT 2035.600 499.840 2035.860 500.100 ;
      LAYER met2 ;
        RECT 1643.110 960.500 1643.390 964.000 ;
        RECT 1643.110 960.000 1643.420 960.500 ;
        RECT 1643.280 947.230 1643.420 960.000 ;
        RECT 1643.220 946.910 1643.480 947.230 ;
        RECT 1648.740 946.910 1649.000 947.230 ;
        RECT 1648.800 500.130 1648.940 946.910 ;
        RECT 1648.740 499.810 1649.000 500.130 ;
        RECT 2035.600 499.810 2035.860 500.130 ;
        RECT 2035.660 17.410 2035.800 499.810 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.150 541.520 1655.470 541.580 ;
        RECT 2049.370 541.520 2049.690 541.580 ;
        RECT 1655.150 541.380 2049.690 541.520 ;
        RECT 1655.150 541.320 1655.470 541.380 ;
        RECT 2049.370 541.320 2049.690 541.380 ;
      LAYER via ;
        RECT 1655.180 541.320 1655.440 541.580 ;
        RECT 2049.400 541.320 2049.660 541.580 ;
      LAYER met2 ;
        RECT 1655.530 960.570 1655.810 964.000 ;
        RECT 1655.240 960.430 1655.810 960.570 ;
        RECT 1655.240 541.610 1655.380 960.430 ;
        RECT 1655.530 960.000 1655.810 960.430 ;
        RECT 1655.180 541.290 1655.440 541.610 ;
        RECT 2049.400 541.290 2049.660 541.610 ;
        RECT 2049.460 17.410 2049.600 541.290 ;
        RECT 2049.460 17.270 2054.660 17.410 ;
        RECT 2054.520 2.400 2054.660 17.270 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.510 17.580 765.830 17.640 ;
        RECT 769.650 17.580 769.970 17.640 ;
        RECT 765.510 17.440 769.970 17.580 ;
        RECT 765.510 17.380 765.830 17.440 ;
        RECT 769.650 17.380 769.970 17.440 ;
      LAYER via ;
        RECT 765.540 17.380 765.800 17.640 ;
        RECT 769.680 17.380 769.940 17.640 ;
      LAYER met2 ;
        RECT 764.970 960.570 765.250 964.000 ;
        RECT 764.970 960.430 765.740 960.570 ;
        RECT 764.970 960.000 765.250 960.430 ;
        RECT 765.600 17.670 765.740 960.430 ;
        RECT 765.540 17.350 765.800 17.670 ;
        RECT 769.680 17.350 769.940 17.670 ;
        RECT 769.740 2.400 769.880 17.350 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.950 548.660 1669.270 548.720 ;
        RECT 2070.070 548.660 2070.390 548.720 ;
        RECT 1668.950 548.520 2070.390 548.660 ;
        RECT 1668.950 548.460 1669.270 548.520 ;
        RECT 2070.070 548.460 2070.390 548.520 ;
      LAYER via ;
        RECT 1668.980 548.460 1669.240 548.720 ;
        RECT 2070.100 548.460 2070.360 548.720 ;
      LAYER met2 ;
        RECT 1667.950 960.570 1668.230 964.000 ;
        RECT 1667.950 960.430 1669.180 960.570 ;
        RECT 1667.950 960.000 1668.230 960.430 ;
        RECT 1669.040 548.750 1669.180 960.430 ;
        RECT 1668.980 548.430 1669.240 548.750 ;
        RECT 2070.100 548.430 2070.360 548.750 ;
        RECT 2070.160 17.410 2070.300 548.430 ;
        RECT 2070.160 17.270 2072.600 17.410 ;
        RECT 2072.460 2.400 2072.600 17.270 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 507.180 1683.530 507.240 ;
        RECT 2083.870 507.180 2084.190 507.240 ;
        RECT 1683.210 507.040 2084.190 507.180 ;
        RECT 1683.210 506.980 1683.530 507.040 ;
        RECT 2083.870 506.980 2084.190 507.040 ;
        RECT 2083.870 16.900 2084.190 16.960 ;
        RECT 2089.850 16.900 2090.170 16.960 ;
        RECT 2083.870 16.760 2090.170 16.900 ;
        RECT 2083.870 16.700 2084.190 16.760 ;
        RECT 2089.850 16.700 2090.170 16.760 ;
      LAYER via ;
        RECT 1683.240 506.980 1683.500 507.240 ;
        RECT 2083.900 506.980 2084.160 507.240 ;
        RECT 2083.900 16.700 2084.160 16.960 ;
        RECT 2089.880 16.700 2090.140 16.960 ;
      LAYER met2 ;
        RECT 1680.370 960.570 1680.650 964.000 ;
        RECT 1680.370 960.430 1683.440 960.570 ;
        RECT 1680.370 960.000 1680.650 960.430 ;
        RECT 1683.300 507.270 1683.440 960.430 ;
        RECT 1683.240 506.950 1683.500 507.270 ;
        RECT 2083.900 506.950 2084.160 507.270 ;
        RECT 2083.960 16.990 2084.100 506.950 ;
        RECT 2083.900 16.670 2084.160 16.990 ;
        RECT 2089.880 16.670 2090.140 16.990 ;
        RECT 2089.940 2.400 2090.080 16.670 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1692.410 945.440 1692.730 945.500 ;
        RECT 1696.550 945.440 1696.870 945.500 ;
        RECT 1692.410 945.300 1696.870 945.440 ;
        RECT 1692.410 945.240 1692.730 945.300 ;
        RECT 1696.550 945.240 1696.870 945.300 ;
        RECT 1696.550 513.980 1696.870 514.040 ;
        RECT 2104.570 513.980 2104.890 514.040 ;
        RECT 1696.550 513.840 2104.890 513.980 ;
        RECT 1696.550 513.780 1696.870 513.840 ;
        RECT 2104.570 513.780 2104.890 513.840 ;
      LAYER via ;
        RECT 1692.440 945.240 1692.700 945.500 ;
        RECT 1696.580 945.240 1696.840 945.500 ;
        RECT 1696.580 513.780 1696.840 514.040 ;
        RECT 2104.600 513.780 2104.860 514.040 ;
      LAYER met2 ;
        RECT 1692.330 960.500 1692.610 964.000 ;
        RECT 1692.330 960.000 1692.640 960.500 ;
        RECT 1692.500 945.530 1692.640 960.000 ;
        RECT 1692.440 945.210 1692.700 945.530 ;
        RECT 1696.580 945.210 1696.840 945.530 ;
        RECT 1696.640 514.070 1696.780 945.210 ;
        RECT 1696.580 513.750 1696.840 514.070 ;
        RECT 2104.600 513.750 2104.860 514.070 ;
        RECT 2104.660 17.410 2104.800 513.750 ;
        RECT 2104.660 17.270 2108.020 17.410 ;
        RECT 2107.880 2.400 2108.020 17.270 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1704.830 949.860 1705.150 949.920 ;
        RECT 1710.350 949.860 1710.670 949.920 ;
        RECT 1704.830 949.720 1710.670 949.860 ;
        RECT 1704.830 949.660 1705.150 949.720 ;
        RECT 1710.350 949.660 1710.670 949.720 ;
        RECT 1710.350 534.720 1710.670 534.780 ;
        RECT 2125.270 534.720 2125.590 534.780 ;
        RECT 1710.350 534.580 2125.590 534.720 ;
        RECT 1710.350 534.520 1710.670 534.580 ;
        RECT 2125.270 534.520 2125.590 534.580 ;
      LAYER via ;
        RECT 1704.860 949.660 1705.120 949.920 ;
        RECT 1710.380 949.660 1710.640 949.920 ;
        RECT 1710.380 534.520 1710.640 534.780 ;
        RECT 2125.300 534.520 2125.560 534.780 ;
      LAYER met2 ;
        RECT 1704.750 960.500 1705.030 964.000 ;
        RECT 1704.750 960.000 1705.060 960.500 ;
        RECT 1704.920 949.950 1705.060 960.000 ;
        RECT 1704.860 949.630 1705.120 949.950 ;
        RECT 1710.380 949.630 1710.640 949.950 ;
        RECT 1710.440 534.810 1710.580 949.630 ;
        RECT 1710.380 534.490 1710.640 534.810 ;
        RECT 2125.300 534.490 2125.560 534.810 ;
        RECT 2125.360 17.410 2125.500 534.490 ;
        RECT 2125.360 17.270 2125.960 17.410 ;
        RECT 2125.820 2.400 2125.960 17.270 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 562.260 1718.030 562.320 ;
        RECT 2139.070 562.260 2139.390 562.320 ;
        RECT 1717.710 562.120 2139.390 562.260 ;
        RECT 1717.710 562.060 1718.030 562.120 ;
        RECT 2139.070 562.060 2139.390 562.120 ;
      LAYER via ;
        RECT 1717.740 562.060 1718.000 562.320 ;
        RECT 2139.100 562.060 2139.360 562.320 ;
      LAYER met2 ;
        RECT 1717.170 960.570 1717.450 964.000 ;
        RECT 1717.170 960.430 1717.940 960.570 ;
        RECT 1717.170 960.000 1717.450 960.430 ;
        RECT 1717.800 562.350 1717.940 960.430 ;
        RECT 1717.740 562.030 1718.000 562.350 ;
        RECT 2139.100 562.030 2139.360 562.350 ;
        RECT 2139.160 17.410 2139.300 562.030 ;
        RECT 2139.160 17.270 2143.900 17.410 ;
        RECT 2143.760 2.400 2143.900 17.270 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.510 251.840 1731.830 251.900 ;
        RECT 2159.770 251.840 2160.090 251.900 ;
        RECT 1731.510 251.700 2160.090 251.840 ;
        RECT 1731.510 251.640 1731.830 251.700 ;
        RECT 2159.770 251.640 2160.090 251.700 ;
      LAYER via ;
        RECT 1731.540 251.640 1731.800 251.900 ;
        RECT 2159.800 251.640 2160.060 251.900 ;
      LAYER met2 ;
        RECT 1729.590 960.570 1729.870 964.000 ;
        RECT 1729.590 960.430 1731.740 960.570 ;
        RECT 1729.590 960.000 1729.870 960.430 ;
        RECT 1731.600 251.930 1731.740 960.430 ;
        RECT 1731.540 251.610 1731.800 251.930 ;
        RECT 2159.800 251.610 2160.060 251.930 ;
        RECT 2159.860 17.410 2160.000 251.610 ;
        RECT 2159.860 17.270 2161.840 17.410 ;
        RECT 2161.700 2.400 2161.840 17.270 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.310 527.920 1745.630 527.980 ;
        RECT 2173.570 527.920 2173.890 527.980 ;
        RECT 1745.310 527.780 2173.890 527.920 ;
        RECT 1745.310 527.720 1745.630 527.780 ;
        RECT 2173.570 527.720 2173.890 527.780 ;
      LAYER via ;
        RECT 1745.340 527.720 1745.600 527.980 ;
        RECT 2173.600 527.720 2173.860 527.980 ;
      LAYER met2 ;
        RECT 1742.010 960.570 1742.290 964.000 ;
        RECT 1742.010 960.430 1745.540 960.570 ;
        RECT 1742.010 960.000 1742.290 960.430 ;
        RECT 1745.400 528.010 1745.540 960.430 ;
        RECT 1745.340 527.690 1745.600 528.010 ;
        RECT 2173.600 527.690 2173.860 528.010 ;
        RECT 2173.660 17.410 2173.800 527.690 ;
        RECT 2173.660 17.270 2179.320 17.410 ;
        RECT 2179.180 2.400 2179.320 17.270 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.510 945.440 1754.830 945.500 ;
        RECT 1758.650 945.440 1758.970 945.500 ;
        RECT 1754.510 945.300 1758.970 945.440 ;
        RECT 1754.510 945.240 1754.830 945.300 ;
        RECT 1758.650 945.240 1758.970 945.300 ;
        RECT 1758.650 569.060 1758.970 569.120 ;
        RECT 2194.270 569.060 2194.590 569.120 ;
        RECT 1758.650 568.920 2194.590 569.060 ;
        RECT 1758.650 568.860 1758.970 568.920 ;
        RECT 2194.270 568.860 2194.590 568.920 ;
      LAYER via ;
        RECT 1754.540 945.240 1754.800 945.500 ;
        RECT 1758.680 945.240 1758.940 945.500 ;
        RECT 1758.680 568.860 1758.940 569.120 ;
        RECT 2194.300 568.860 2194.560 569.120 ;
      LAYER met2 ;
        RECT 1754.430 960.500 1754.710 964.000 ;
        RECT 1754.430 960.000 1754.740 960.500 ;
        RECT 1754.600 945.530 1754.740 960.000 ;
        RECT 1754.540 945.210 1754.800 945.530 ;
        RECT 1758.680 945.210 1758.940 945.530 ;
        RECT 1758.740 569.150 1758.880 945.210 ;
        RECT 1758.680 568.830 1758.940 569.150 ;
        RECT 2194.300 568.830 2194.560 569.150 ;
        RECT 2194.360 17.410 2194.500 568.830 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.930 950.540 1767.250 950.600 ;
        RECT 1772.450 950.540 1772.770 950.600 ;
        RECT 1766.930 950.400 1772.770 950.540 ;
        RECT 1766.930 950.340 1767.250 950.400 ;
        RECT 1772.450 950.340 1772.770 950.400 ;
        RECT 1772.450 831.540 1772.770 831.600 ;
        RECT 2214.970 831.540 2215.290 831.600 ;
        RECT 1772.450 831.400 2215.290 831.540 ;
        RECT 1772.450 831.340 1772.770 831.400 ;
        RECT 2214.970 831.340 2215.290 831.400 ;
      LAYER via ;
        RECT 1766.960 950.340 1767.220 950.600 ;
        RECT 1772.480 950.340 1772.740 950.600 ;
        RECT 1772.480 831.340 1772.740 831.600 ;
        RECT 2215.000 831.340 2215.260 831.600 ;
      LAYER met2 ;
        RECT 1766.850 960.500 1767.130 964.000 ;
        RECT 1766.850 960.000 1767.160 960.500 ;
        RECT 1767.020 950.630 1767.160 960.000 ;
        RECT 1766.960 950.310 1767.220 950.630 ;
        RECT 1772.480 950.310 1772.740 950.630 ;
        RECT 1772.540 831.630 1772.680 950.310 ;
        RECT 1772.480 831.310 1772.740 831.630 ;
        RECT 2215.000 831.310 2215.260 831.630 ;
        RECT 2215.060 2.400 2215.200 831.310 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.910 17.580 2233.230 17.640 ;
        RECT 1787.720 17.440 2233.230 17.580 ;
        RECT 1779.810 17.240 1780.130 17.300 ;
        RECT 1787.720 17.240 1787.860 17.440 ;
        RECT 2232.910 17.380 2233.230 17.440 ;
        RECT 1779.810 17.100 1787.860 17.240 ;
        RECT 1779.810 17.040 1780.130 17.100 ;
      LAYER via ;
        RECT 1779.840 17.040 1780.100 17.300 ;
        RECT 2232.940 17.380 2233.200 17.640 ;
      LAYER met2 ;
        RECT 1779.270 960.570 1779.550 964.000 ;
        RECT 1779.270 960.430 1780.040 960.570 ;
        RECT 1779.270 960.000 1779.550 960.430 ;
        RECT 1779.900 17.330 1780.040 960.430 ;
        RECT 2232.940 17.350 2233.200 17.670 ;
        RECT 1779.840 17.010 1780.100 17.330 ;
        RECT 2233.000 2.400 2233.140 17.350 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 16.560 779.630 16.620 ;
        RECT 787.590 16.560 787.910 16.620 ;
        RECT 779.310 16.420 787.910 16.560 ;
        RECT 779.310 16.360 779.630 16.420 ;
        RECT 787.590 16.360 787.910 16.420 ;
      LAYER via ;
        RECT 779.340 16.360 779.600 16.620 ;
        RECT 787.620 16.360 787.880 16.620 ;
      LAYER met2 ;
        RECT 776.930 960.570 777.210 964.000 ;
        RECT 776.930 960.430 779.540 960.570 ;
        RECT 776.930 960.000 777.210 960.430 ;
        RECT 779.400 16.650 779.540 960.430 ;
        RECT 779.340 16.330 779.600 16.650 ;
        RECT 787.620 16.330 787.880 16.650 ;
        RECT 787.680 2.400 787.820 16.330 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 17.240 1793.930 17.300 ;
        RECT 2250.850 17.240 2251.170 17.300 ;
        RECT 1793.610 17.100 2251.170 17.240 ;
        RECT 1793.610 17.040 1793.930 17.100 ;
        RECT 2250.850 17.040 2251.170 17.100 ;
      LAYER via ;
        RECT 1793.640 17.040 1793.900 17.300 ;
        RECT 2250.880 17.040 2251.140 17.300 ;
      LAYER met2 ;
        RECT 1791.690 960.570 1791.970 964.000 ;
        RECT 1791.690 960.430 1793.840 960.570 ;
        RECT 1791.690 960.000 1791.970 960.430 ;
        RECT 1793.700 17.330 1793.840 960.430 ;
        RECT 1793.640 17.010 1793.900 17.330 ;
        RECT 2250.880 17.010 2251.140 17.330 ;
        RECT 2250.940 2.400 2251.080 17.010 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.410 20.640 1807.730 20.700 ;
        RECT 2268.330 20.640 2268.650 20.700 ;
        RECT 1807.410 20.500 2268.650 20.640 ;
        RECT 1807.410 20.440 1807.730 20.500 ;
        RECT 2268.330 20.440 2268.650 20.500 ;
      LAYER via ;
        RECT 1807.440 20.440 1807.700 20.700 ;
        RECT 2268.360 20.440 2268.620 20.700 ;
      LAYER met2 ;
        RECT 1803.650 960.570 1803.930 964.000 ;
        RECT 1803.650 960.430 1807.640 960.570 ;
        RECT 1803.650 960.000 1803.930 960.430 ;
        RECT 1807.500 20.730 1807.640 960.430 ;
        RECT 1807.440 20.410 1807.700 20.730 ;
        RECT 2268.360 20.410 2268.620 20.730 ;
        RECT 2268.420 2.400 2268.560 20.410 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1816.150 945.440 1816.470 945.500 ;
        RECT 1821.210 945.440 1821.530 945.500 ;
        RECT 1816.150 945.300 1821.530 945.440 ;
        RECT 1816.150 945.240 1816.470 945.300 ;
        RECT 1821.210 945.240 1821.530 945.300 ;
        RECT 1821.210 20.300 1821.530 20.360 ;
        RECT 2286.270 20.300 2286.590 20.360 ;
        RECT 1821.210 20.160 2286.590 20.300 ;
        RECT 1821.210 20.100 1821.530 20.160 ;
        RECT 2286.270 20.100 2286.590 20.160 ;
      LAYER via ;
        RECT 1816.180 945.240 1816.440 945.500 ;
        RECT 1821.240 945.240 1821.500 945.500 ;
        RECT 1821.240 20.100 1821.500 20.360 ;
        RECT 2286.300 20.100 2286.560 20.360 ;
      LAYER met2 ;
        RECT 1816.070 960.500 1816.350 964.000 ;
        RECT 1816.070 960.000 1816.380 960.500 ;
        RECT 1816.240 945.530 1816.380 960.000 ;
        RECT 1816.180 945.210 1816.440 945.530 ;
        RECT 1821.240 945.210 1821.500 945.530 ;
        RECT 1821.300 20.390 1821.440 945.210 ;
        RECT 1821.240 20.070 1821.500 20.390 ;
        RECT 2286.300 20.070 2286.560 20.390 ;
        RECT 2286.360 2.400 2286.500 20.070 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.570 946.460 1828.890 946.520 ;
        RECT 1835.010 946.460 1835.330 946.520 ;
        RECT 1828.570 946.320 1835.330 946.460 ;
        RECT 1828.570 946.260 1828.890 946.320 ;
        RECT 1835.010 946.260 1835.330 946.320 ;
        RECT 1835.010 19.960 1835.330 20.020 ;
        RECT 2304.210 19.960 2304.530 20.020 ;
        RECT 1835.010 19.820 2304.530 19.960 ;
        RECT 1835.010 19.760 1835.330 19.820 ;
        RECT 2304.210 19.760 2304.530 19.820 ;
      LAYER via ;
        RECT 1828.600 946.260 1828.860 946.520 ;
        RECT 1835.040 946.260 1835.300 946.520 ;
        RECT 1835.040 19.760 1835.300 20.020 ;
        RECT 2304.240 19.760 2304.500 20.020 ;
      LAYER met2 ;
        RECT 1828.490 960.500 1828.770 964.000 ;
        RECT 1828.490 960.000 1828.800 960.500 ;
        RECT 1828.660 946.550 1828.800 960.000 ;
        RECT 1828.600 946.230 1828.860 946.550 ;
        RECT 1835.040 946.230 1835.300 946.550 ;
        RECT 1835.100 20.050 1835.240 946.230 ;
        RECT 1835.040 19.730 1835.300 20.050 ;
        RECT 2304.240 19.730 2304.500 20.050 ;
        RECT 2304.300 2.400 2304.440 19.730 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1841.910 19.620 1842.230 19.680 ;
        RECT 2322.150 19.620 2322.470 19.680 ;
        RECT 1841.910 19.480 2322.470 19.620 ;
        RECT 1841.910 19.420 1842.230 19.480 ;
        RECT 2322.150 19.420 2322.470 19.480 ;
      LAYER via ;
        RECT 1841.940 19.420 1842.200 19.680 ;
        RECT 2322.180 19.420 2322.440 19.680 ;
      LAYER met2 ;
        RECT 1840.910 960.570 1841.190 964.000 ;
        RECT 1840.910 960.430 1842.140 960.570 ;
        RECT 1840.910 960.000 1841.190 960.430 ;
        RECT 1842.000 19.710 1842.140 960.430 ;
        RECT 1841.940 19.390 1842.200 19.710 ;
        RECT 2322.180 19.390 2322.440 19.710 ;
        RECT 2322.240 2.400 2322.380 19.390 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.710 18.940 1856.030 19.000 ;
        RECT 2339.170 18.940 2339.490 19.000 ;
        RECT 1855.710 18.800 2339.490 18.940 ;
        RECT 1855.710 18.740 1856.030 18.800 ;
        RECT 2339.170 18.740 2339.490 18.800 ;
      LAYER via ;
        RECT 1855.740 18.740 1856.000 19.000 ;
        RECT 2339.200 18.740 2339.460 19.000 ;
      LAYER met2 ;
        RECT 1853.330 960.570 1853.610 964.000 ;
        RECT 1853.330 960.430 1855.940 960.570 ;
        RECT 1853.330 960.000 1853.610 960.430 ;
        RECT 1855.800 19.030 1855.940 960.430 ;
        RECT 1855.740 18.710 1856.000 19.030 ;
        RECT 2339.200 18.710 2339.460 19.030 ;
        RECT 2339.260 16.050 2339.400 18.710 ;
        RECT 2339.260 15.910 2339.860 16.050 ;
        RECT 2339.720 2.400 2339.860 15.910 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1865.830 949.860 1866.150 949.920 ;
        RECT 1869.510 949.860 1869.830 949.920 ;
        RECT 1865.830 949.720 1869.830 949.860 ;
        RECT 1865.830 949.660 1866.150 949.720 ;
        RECT 1869.510 949.660 1869.830 949.720 ;
        RECT 1869.510 19.280 1869.830 19.340 ;
        RECT 2357.570 19.280 2357.890 19.340 ;
        RECT 1869.510 19.140 2357.890 19.280 ;
        RECT 1869.510 19.080 1869.830 19.140 ;
        RECT 2357.570 19.080 2357.890 19.140 ;
      LAYER via ;
        RECT 1865.860 949.660 1866.120 949.920 ;
        RECT 1869.540 949.660 1869.800 949.920 ;
        RECT 1869.540 19.080 1869.800 19.340 ;
        RECT 2357.600 19.080 2357.860 19.340 ;
      LAYER met2 ;
        RECT 1865.750 960.500 1866.030 964.000 ;
        RECT 1865.750 960.000 1866.060 960.500 ;
        RECT 1865.920 949.950 1866.060 960.000 ;
        RECT 1865.860 949.630 1866.120 949.950 ;
        RECT 1869.540 949.630 1869.800 949.950 ;
        RECT 1869.600 19.370 1869.740 949.630 ;
        RECT 1869.540 19.050 1869.800 19.370 ;
        RECT 2357.600 19.050 2357.860 19.370 ;
        RECT 2357.660 2.400 2357.800 19.050 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1878.250 951.220 1878.570 951.280 ;
        RECT 1883.310 951.220 1883.630 951.280 ;
        RECT 1878.250 951.080 1883.630 951.220 ;
        RECT 1878.250 951.020 1878.570 951.080 ;
        RECT 1883.310 951.020 1883.630 951.080 ;
        RECT 1883.310 18.260 1883.630 18.320 ;
        RECT 2375.510 18.260 2375.830 18.320 ;
        RECT 1883.310 18.120 2375.830 18.260 ;
        RECT 1883.310 18.060 1883.630 18.120 ;
        RECT 2375.510 18.060 2375.830 18.120 ;
      LAYER via ;
        RECT 1878.280 951.020 1878.540 951.280 ;
        RECT 1883.340 951.020 1883.600 951.280 ;
        RECT 1883.340 18.060 1883.600 18.320 ;
        RECT 2375.540 18.060 2375.800 18.320 ;
      LAYER met2 ;
        RECT 1878.170 960.500 1878.450 964.000 ;
        RECT 1878.170 960.000 1878.480 960.500 ;
        RECT 1878.340 951.310 1878.480 960.000 ;
        RECT 1878.280 950.990 1878.540 951.310 ;
        RECT 1883.340 950.990 1883.600 951.310 ;
        RECT 1883.400 18.350 1883.540 950.990 ;
        RECT 1883.340 18.030 1883.600 18.350 ;
        RECT 2375.540 18.030 2375.800 18.350 ;
        RECT 2375.600 2.400 2375.740 18.030 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1890.670 946.460 1890.990 946.520 ;
        RECT 1897.110 946.460 1897.430 946.520 ;
        RECT 1890.670 946.320 1897.430 946.460 ;
        RECT 1890.670 946.260 1890.990 946.320 ;
        RECT 1897.110 946.260 1897.430 946.320 ;
        RECT 1897.110 18.600 1897.430 18.660 ;
        RECT 2393.450 18.600 2393.770 18.660 ;
        RECT 1897.110 18.460 2393.770 18.600 ;
        RECT 1897.110 18.400 1897.430 18.460 ;
        RECT 2393.450 18.400 2393.770 18.460 ;
      LAYER via ;
        RECT 1890.700 946.260 1890.960 946.520 ;
        RECT 1897.140 946.260 1897.400 946.520 ;
        RECT 1897.140 18.400 1897.400 18.660 ;
        RECT 2393.480 18.400 2393.740 18.660 ;
      LAYER met2 ;
        RECT 1890.590 960.500 1890.870 964.000 ;
        RECT 1890.590 960.000 1890.900 960.500 ;
        RECT 1890.760 946.550 1890.900 960.000 ;
        RECT 1890.700 946.230 1890.960 946.550 ;
        RECT 1897.140 946.230 1897.400 946.550 ;
        RECT 1897.200 18.690 1897.340 946.230 ;
        RECT 1897.140 18.370 1897.400 18.690 ;
        RECT 2393.480 18.370 2393.740 18.690 ;
        RECT 2393.540 2.400 2393.680 18.370 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 17.920 1904.330 17.980 ;
        RECT 2411.390 17.920 2411.710 17.980 ;
        RECT 1904.010 17.780 2411.710 17.920 ;
        RECT 1904.010 17.720 1904.330 17.780 ;
        RECT 2411.390 17.720 2411.710 17.780 ;
      LAYER via ;
        RECT 1904.040 17.720 1904.300 17.980 ;
        RECT 2411.420 17.720 2411.680 17.980 ;
      LAYER met2 ;
        RECT 1903.010 960.570 1903.290 964.000 ;
        RECT 1903.010 960.430 1904.240 960.570 ;
        RECT 1903.010 960.000 1903.290 960.430 ;
        RECT 1904.100 18.010 1904.240 960.430 ;
        RECT 1904.040 17.690 1904.300 18.010 ;
        RECT 2411.420 17.690 2411.680 18.010 ;
        RECT 2411.480 2.400 2411.620 17.690 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 789.430 945.440 789.750 945.500 ;
        RECT 793.110 945.440 793.430 945.500 ;
        RECT 789.430 945.300 793.430 945.440 ;
        RECT 789.430 945.240 789.750 945.300 ;
        RECT 793.110 945.240 793.430 945.300 ;
        RECT 793.110 17.240 793.430 17.300 ;
        RECT 805.530 17.240 805.850 17.300 ;
        RECT 793.110 17.100 805.850 17.240 ;
        RECT 793.110 17.040 793.430 17.100 ;
        RECT 805.530 17.040 805.850 17.100 ;
      LAYER via ;
        RECT 789.460 945.240 789.720 945.500 ;
        RECT 793.140 945.240 793.400 945.500 ;
        RECT 793.140 17.040 793.400 17.300 ;
        RECT 805.560 17.040 805.820 17.300 ;
      LAYER met2 ;
        RECT 789.350 960.500 789.630 964.000 ;
        RECT 789.350 960.000 789.660 960.500 ;
        RECT 789.520 945.530 789.660 960.000 ;
        RECT 789.460 945.210 789.720 945.530 ;
        RECT 793.140 945.210 793.400 945.530 ;
        RECT 793.200 17.330 793.340 945.210 ;
        RECT 793.140 17.010 793.400 17.330 ;
        RECT 805.560 17.010 805.820 17.330 ;
        RECT 805.620 2.400 805.760 17.010 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 655.570 17.240 655.890 17.300 ;
        RECT 2.830 17.100 655.890 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 655.570 17.040 655.890 17.100 ;
      LAYER via ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 655.600 17.040 655.860 17.300 ;
      LAYER met2 ;
        RECT 661.930 960.570 662.210 964.000 ;
        RECT 655.660 960.430 662.210 960.570 ;
        RECT 655.660 17.330 655.800 960.430 ;
        RECT 661.930 960.000 662.210 960.430 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 655.600 17.010 655.860 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 662.470 17.580 662.790 17.640 ;
        RECT 8.350 17.440 662.790 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 662.470 17.380 662.790 17.440 ;
      LAYER via ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 662.500 17.380 662.760 17.640 ;
      LAYER met2 ;
        RECT 665.610 960.570 665.890 964.000 ;
        RECT 662.560 960.430 665.890 960.570 ;
        RECT 662.560 17.670 662.700 960.430 ;
        RECT 665.610 960.000 665.890 960.430 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 662.500 17.350 662.760 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.580 -14.220 -16.580 3533.900 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.420 7.020 3529.100 ;
        RECT 22.020 -19.020 25.020 3538.700 ;
        RECT 184.020 -9.420 187.020 3529.100 ;
        RECT 202.020 -19.020 205.020 3538.700 ;
        RECT 364.020 -9.420 367.020 3529.100 ;
        RECT 382.020 -19.020 385.020 3538.700 ;
        RECT 544.020 -9.420 547.020 3529.100 ;
        RECT 562.020 -19.020 565.020 3538.700 ;
        RECT 724.020 2562.185 727.020 3529.100 ;
        RECT 742.020 2562.185 745.020 3538.700 ;
        RECT 904.020 2562.185 907.020 3529.100 ;
        RECT 922.020 2562.185 925.020 3538.700 ;
        RECT 1084.020 2562.185 1087.020 3529.100 ;
        RECT 1102.020 2562.185 1105.020 3538.700 ;
        RECT 1264.020 2562.185 1267.020 3529.100 ;
        RECT 1282.020 2562.185 1285.020 3538.700 ;
        RECT 1444.020 2562.185 1447.020 3529.100 ;
        RECT 1462.020 2562.185 1465.020 3538.700 ;
        RECT 1624.020 2562.185 1627.020 3529.100 ;
        RECT 1642.020 2562.185 1645.020 3538.700 ;
        RECT 1804.020 2562.185 1807.020 3529.100 ;
        RECT 1822.020 2562.185 1825.020 3538.700 ;
        RECT 1984.020 2562.185 1987.020 3529.100 ;
        RECT 2002.020 2562.185 2005.020 3538.700 ;
        RECT 2164.020 2562.185 2167.020 3529.100 ;
        RECT 2182.020 2562.185 2185.020 3538.700 ;
        RECT 681.040 970.640 682.640 2551.440 ;
        RECT 724.020 -9.420 727.020 960.000 ;
        RECT 742.020 -19.020 745.020 960.000 ;
        RECT 904.020 -9.420 907.020 960.000 ;
        RECT 922.020 -19.020 925.020 960.000 ;
        RECT 1084.020 -9.420 1087.020 960.000 ;
        RECT 1102.020 -19.020 1105.020 960.000 ;
        RECT 1264.020 -9.420 1267.020 960.000 ;
        RECT 1282.020 -19.020 1285.020 960.000 ;
        RECT 1444.020 -9.420 1447.020 960.000 ;
        RECT 1462.020 -19.020 1465.020 960.000 ;
        RECT 1624.020 -9.420 1627.020 960.000 ;
        RECT 1642.020 -19.020 1645.020 960.000 ;
        RECT 1804.020 -9.420 1807.020 960.000 ;
        RECT 1822.020 -19.020 1825.020 960.000 ;
        RECT 1984.020 -9.420 1987.020 960.000 ;
        RECT 2002.020 -19.020 2005.020 960.000 ;
        RECT 2164.020 -9.420 2167.020 960.000 ;
        RECT 2182.020 -19.020 2185.020 960.000 ;
        RECT 2344.020 -9.420 2347.020 3529.100 ;
        RECT 2362.020 -19.020 2365.020 3538.700 ;
        RECT 2524.020 -9.420 2527.020 3529.100 ;
        RECT 2542.020 -19.020 2545.020 3538.700 ;
        RECT 2704.020 -9.420 2707.020 3529.100 ;
        RECT 2722.020 -19.020 2725.020 3538.700 ;
        RECT 2884.020 -9.420 2887.020 3529.100 ;
        RECT 2902.020 -19.020 2905.020 3538.700 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.200 -14.220 2939.200 3533.900 ;
      LAYER via4 ;
        RECT -18.670 3532.610 -17.490 3533.790 ;
        RECT -18.670 3531.010 -17.490 3532.190 ;
        RECT 22.930 3532.610 24.110 3533.790 ;
        RECT 22.930 3531.010 24.110 3532.190 ;
        RECT -18.670 3449.090 -17.490 3450.270 ;
        RECT -18.670 3447.490 -17.490 3448.670 ;
        RECT -18.670 3269.090 -17.490 3270.270 ;
        RECT -18.670 3267.490 -17.490 3268.670 ;
        RECT -18.670 3089.090 -17.490 3090.270 ;
        RECT -18.670 3087.490 -17.490 3088.670 ;
        RECT -18.670 2909.090 -17.490 2910.270 ;
        RECT -18.670 2907.490 -17.490 2908.670 ;
        RECT -18.670 2729.090 -17.490 2730.270 ;
        RECT -18.670 2727.490 -17.490 2728.670 ;
        RECT -18.670 2549.090 -17.490 2550.270 ;
        RECT -18.670 2547.490 -17.490 2548.670 ;
        RECT -18.670 2369.090 -17.490 2370.270 ;
        RECT -18.670 2367.490 -17.490 2368.670 ;
        RECT -18.670 2189.090 -17.490 2190.270 ;
        RECT -18.670 2187.490 -17.490 2188.670 ;
        RECT -18.670 2009.090 -17.490 2010.270 ;
        RECT -18.670 2007.490 -17.490 2008.670 ;
        RECT -18.670 1829.090 -17.490 1830.270 ;
        RECT -18.670 1827.490 -17.490 1828.670 ;
        RECT -18.670 1649.090 -17.490 1650.270 ;
        RECT -18.670 1647.490 -17.490 1648.670 ;
        RECT -18.670 1469.090 -17.490 1470.270 ;
        RECT -18.670 1467.490 -17.490 1468.670 ;
        RECT -18.670 1289.090 -17.490 1290.270 ;
        RECT -18.670 1287.490 -17.490 1288.670 ;
        RECT -18.670 1109.090 -17.490 1110.270 ;
        RECT -18.670 1107.490 -17.490 1108.670 ;
        RECT -18.670 929.090 -17.490 930.270 ;
        RECT -18.670 927.490 -17.490 928.670 ;
        RECT -18.670 749.090 -17.490 750.270 ;
        RECT -18.670 747.490 -17.490 748.670 ;
        RECT -18.670 569.090 -17.490 570.270 ;
        RECT -18.670 567.490 -17.490 568.670 ;
        RECT -18.670 389.090 -17.490 390.270 ;
        RECT -18.670 387.490 -17.490 388.670 ;
        RECT -18.670 209.090 -17.490 210.270 ;
        RECT -18.670 207.490 -17.490 208.670 ;
        RECT -18.670 29.090 -17.490 30.270 ;
        RECT -18.670 27.490 -17.490 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 202.930 3532.610 204.110 3533.790 ;
        RECT 202.930 3531.010 204.110 3532.190 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.670 -12.510 -17.490 -11.330 ;
        RECT -18.670 -14.110 -17.490 -12.930 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 382.930 3532.610 384.110 3533.790 ;
        RECT 382.930 3531.010 384.110 3532.190 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 22.930 -12.510 24.110 -11.330 ;
        RECT 22.930 -14.110 24.110 -12.930 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 562.930 3532.610 564.110 3533.790 ;
        RECT 562.930 3531.010 564.110 3532.190 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 202.930 -12.510 204.110 -11.330 ;
        RECT 202.930 -14.110 204.110 -12.930 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 742.930 3532.610 744.110 3533.790 ;
        RECT 742.930 3531.010 744.110 3532.190 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 922.930 3532.610 924.110 3533.790 ;
        RECT 922.930 3531.010 924.110 3532.190 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 1102.930 3532.610 1104.110 3533.790 ;
        RECT 1102.930 3531.010 1104.110 3532.190 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1282.930 3532.610 1284.110 3533.790 ;
        RECT 1282.930 3531.010 1284.110 3532.190 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1462.930 3532.610 1464.110 3533.790 ;
        RECT 1462.930 3531.010 1464.110 3532.190 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1642.930 3532.610 1644.110 3533.790 ;
        RECT 1642.930 3531.010 1644.110 3532.190 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1822.930 3532.610 1824.110 3533.790 ;
        RECT 1822.930 3531.010 1824.110 3532.190 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 2002.930 3532.610 2004.110 3533.790 ;
        RECT 2002.930 3531.010 2004.110 3532.190 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 2182.930 3532.610 2184.110 3533.790 ;
        RECT 2182.930 3531.010 2184.110 3532.190 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2362.930 3532.610 2364.110 3533.790 ;
        RECT 2362.930 3531.010 2364.110 3532.190 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 681.250 2549.090 682.430 2550.270 ;
        RECT 681.250 2547.490 682.430 2548.670 ;
        RECT 681.250 2531.090 682.430 2532.270 ;
        RECT 681.250 2529.490 682.430 2530.670 ;
        RECT 681.250 2369.090 682.430 2370.270 ;
        RECT 681.250 2367.490 682.430 2368.670 ;
        RECT 681.250 2351.090 682.430 2352.270 ;
        RECT 681.250 2349.490 682.430 2350.670 ;
        RECT 681.250 2189.090 682.430 2190.270 ;
        RECT 681.250 2187.490 682.430 2188.670 ;
        RECT 681.250 2171.090 682.430 2172.270 ;
        RECT 681.250 2169.490 682.430 2170.670 ;
        RECT 681.250 2009.090 682.430 2010.270 ;
        RECT 681.250 2007.490 682.430 2008.670 ;
        RECT 681.250 1991.090 682.430 1992.270 ;
        RECT 681.250 1989.490 682.430 1990.670 ;
        RECT 681.250 1829.090 682.430 1830.270 ;
        RECT 681.250 1827.490 682.430 1828.670 ;
        RECT 681.250 1811.090 682.430 1812.270 ;
        RECT 681.250 1809.490 682.430 1810.670 ;
        RECT 681.250 1649.090 682.430 1650.270 ;
        RECT 681.250 1647.490 682.430 1648.670 ;
        RECT 681.250 1631.090 682.430 1632.270 ;
        RECT 681.250 1629.490 682.430 1630.670 ;
        RECT 681.250 1469.090 682.430 1470.270 ;
        RECT 681.250 1467.490 682.430 1468.670 ;
        RECT 681.250 1451.090 682.430 1452.270 ;
        RECT 681.250 1449.490 682.430 1450.670 ;
        RECT 681.250 1289.090 682.430 1290.270 ;
        RECT 681.250 1287.490 682.430 1288.670 ;
        RECT 681.250 1271.090 682.430 1272.270 ;
        RECT 681.250 1269.490 682.430 1270.670 ;
        RECT 681.250 1109.090 682.430 1110.270 ;
        RECT 681.250 1107.490 682.430 1108.670 ;
        RECT 681.250 1091.090 682.430 1092.270 ;
        RECT 681.250 1089.490 682.430 1090.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 382.930 -12.510 384.110 -11.330 ;
        RECT 382.930 -14.110 384.110 -12.930 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 562.930 -12.510 564.110 -11.330 ;
        RECT 562.930 -14.110 564.110 -12.930 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 742.930 -12.510 744.110 -11.330 ;
        RECT 742.930 -14.110 744.110 -12.930 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 922.930 -12.510 924.110 -11.330 ;
        RECT 922.930 -14.110 924.110 -12.930 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1102.930 -12.510 1104.110 -11.330 ;
        RECT 1102.930 -14.110 1104.110 -12.930 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1282.930 -12.510 1284.110 -11.330 ;
        RECT 1282.930 -14.110 1284.110 -12.930 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1462.930 -12.510 1464.110 -11.330 ;
        RECT 1462.930 -14.110 1464.110 -12.930 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1642.930 -12.510 1644.110 -11.330 ;
        RECT 1642.930 -14.110 1644.110 -12.930 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 1822.930 -12.510 1824.110 -11.330 ;
        RECT 1822.930 -14.110 1824.110 -12.930 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2002.930 -12.510 2004.110 -11.330 ;
        RECT 2002.930 -14.110 2004.110 -12.930 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2542.930 3532.610 2544.110 3533.790 ;
        RECT 2542.930 3531.010 2544.110 3532.190 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2182.930 -12.510 2184.110 -11.330 ;
        RECT 2182.930 -14.110 2184.110 -12.930 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2722.930 3532.610 2724.110 3533.790 ;
        RECT 2722.930 3531.010 2724.110 3532.190 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2362.930 -12.510 2364.110 -11.330 ;
        RECT 2362.930 -14.110 2364.110 -12.930 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2902.930 3532.610 2904.110 3533.790 ;
        RECT 2902.930 3531.010 2904.110 3532.190 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2542.930 -12.510 2544.110 -11.330 ;
        RECT 2542.930 -14.110 2544.110 -12.930 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2937.110 3532.610 2938.290 3533.790 ;
        RECT 2937.110 3531.010 2938.290 3532.190 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2722.930 -12.510 2724.110 -11.330 ;
        RECT 2722.930 -14.110 2724.110 -12.930 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2937.110 3449.090 2938.290 3450.270 ;
        RECT 2937.110 3447.490 2938.290 3448.670 ;
        RECT 2937.110 3269.090 2938.290 3270.270 ;
        RECT 2937.110 3267.490 2938.290 3268.670 ;
        RECT 2937.110 3089.090 2938.290 3090.270 ;
        RECT 2937.110 3087.490 2938.290 3088.670 ;
        RECT 2937.110 2909.090 2938.290 2910.270 ;
        RECT 2937.110 2907.490 2938.290 2908.670 ;
        RECT 2937.110 2729.090 2938.290 2730.270 ;
        RECT 2937.110 2727.490 2938.290 2728.670 ;
        RECT 2937.110 2549.090 2938.290 2550.270 ;
        RECT 2937.110 2547.490 2938.290 2548.670 ;
        RECT 2937.110 2369.090 2938.290 2370.270 ;
        RECT 2937.110 2367.490 2938.290 2368.670 ;
        RECT 2937.110 2189.090 2938.290 2190.270 ;
        RECT 2937.110 2187.490 2938.290 2188.670 ;
        RECT 2937.110 2009.090 2938.290 2010.270 ;
        RECT 2937.110 2007.490 2938.290 2008.670 ;
        RECT 2937.110 1829.090 2938.290 1830.270 ;
        RECT 2937.110 1827.490 2938.290 1828.670 ;
        RECT 2937.110 1649.090 2938.290 1650.270 ;
        RECT 2937.110 1647.490 2938.290 1648.670 ;
        RECT 2937.110 1469.090 2938.290 1470.270 ;
        RECT 2937.110 1467.490 2938.290 1468.670 ;
        RECT 2937.110 1289.090 2938.290 1290.270 ;
        RECT 2937.110 1287.490 2938.290 1288.670 ;
        RECT 2937.110 1109.090 2938.290 1110.270 ;
        RECT 2937.110 1107.490 2938.290 1108.670 ;
        RECT 2937.110 929.090 2938.290 930.270 ;
        RECT 2937.110 927.490 2938.290 928.670 ;
        RECT 2937.110 749.090 2938.290 750.270 ;
        RECT 2937.110 747.490 2938.290 748.670 ;
        RECT 2937.110 569.090 2938.290 570.270 ;
        RECT 2937.110 567.490 2938.290 568.670 ;
        RECT 2937.110 389.090 2938.290 390.270 ;
        RECT 2937.110 387.490 2938.290 388.670 ;
        RECT 2937.110 209.090 2938.290 210.270 ;
        RECT 2937.110 207.490 2938.290 208.670 ;
        RECT 2937.110 29.090 2938.290 30.270 ;
        RECT 2937.110 27.490 2938.290 28.670 ;
        RECT 2902.930 -12.510 2904.110 -11.330 ;
        RECT 2902.930 -14.110 2904.110 -12.930 ;
        RECT 2937.110 -12.510 2938.290 -11.330 ;
        RECT 2937.110 -14.110 2938.290 -12.930 ;
      LAYER met5 ;
        RECT -19.580 3533.900 -16.580 3533.910 ;
        RECT 22.020 3533.900 25.020 3533.910 ;
        RECT 202.020 3533.900 205.020 3533.910 ;
        RECT 382.020 3533.900 385.020 3533.910 ;
        RECT 562.020 3533.900 565.020 3533.910 ;
        RECT 742.020 3533.900 745.020 3533.910 ;
        RECT 922.020 3533.900 925.020 3533.910 ;
        RECT 1102.020 3533.900 1105.020 3533.910 ;
        RECT 1282.020 3533.900 1285.020 3533.910 ;
        RECT 1462.020 3533.900 1465.020 3533.910 ;
        RECT 1642.020 3533.900 1645.020 3533.910 ;
        RECT 1822.020 3533.900 1825.020 3533.910 ;
        RECT 2002.020 3533.900 2005.020 3533.910 ;
        RECT 2182.020 3533.900 2185.020 3533.910 ;
        RECT 2362.020 3533.900 2365.020 3533.910 ;
        RECT 2542.020 3533.900 2545.020 3533.910 ;
        RECT 2722.020 3533.900 2725.020 3533.910 ;
        RECT 2902.020 3533.900 2905.020 3533.910 ;
        RECT 2936.200 3533.900 2939.200 3533.910 ;
        RECT -19.580 3530.900 2939.200 3533.900 ;
        RECT -19.580 3530.890 -16.580 3530.900 ;
        RECT 22.020 3530.890 25.020 3530.900 ;
        RECT 202.020 3530.890 205.020 3530.900 ;
        RECT 382.020 3530.890 385.020 3530.900 ;
        RECT 562.020 3530.890 565.020 3530.900 ;
        RECT 742.020 3530.890 745.020 3530.900 ;
        RECT 922.020 3530.890 925.020 3530.900 ;
        RECT 1102.020 3530.890 1105.020 3530.900 ;
        RECT 1282.020 3530.890 1285.020 3530.900 ;
        RECT 1462.020 3530.890 1465.020 3530.900 ;
        RECT 1642.020 3530.890 1645.020 3530.900 ;
        RECT 1822.020 3530.890 1825.020 3530.900 ;
        RECT 2002.020 3530.890 2005.020 3530.900 ;
        RECT 2182.020 3530.890 2185.020 3530.900 ;
        RECT 2362.020 3530.890 2365.020 3530.900 ;
        RECT 2542.020 3530.890 2545.020 3530.900 ;
        RECT 2722.020 3530.890 2725.020 3530.900 ;
        RECT 2902.020 3530.890 2905.020 3530.900 ;
        RECT 2936.200 3530.890 2939.200 3530.900 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -19.580 3450.380 -16.580 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.200 3450.380 2939.200 3450.390 ;
        RECT -24.380 3447.380 2944.000 3450.380 ;
        RECT -19.580 3447.370 -16.580 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.200 3447.370 2939.200 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.780 3429.380 2934.400 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -19.580 3270.380 -16.580 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.200 3270.380 2939.200 3270.390 ;
        RECT -24.380 3267.380 2944.000 3270.380 ;
        RECT -19.580 3267.370 -16.580 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.200 3267.370 2939.200 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.780 3249.380 2934.400 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -19.580 3090.380 -16.580 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.200 3090.380 2939.200 3090.390 ;
        RECT -24.380 3087.380 2944.000 3090.380 ;
        RECT -19.580 3087.370 -16.580 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.200 3087.370 2939.200 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.780 3069.380 2934.400 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -19.580 2910.380 -16.580 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.200 2910.380 2939.200 2910.390 ;
        RECT -24.380 2907.380 2944.000 2910.380 ;
        RECT -19.580 2907.370 -16.580 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.200 2907.370 2939.200 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.780 2889.380 2934.400 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -19.580 2730.380 -16.580 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.200 2730.380 2939.200 2730.390 ;
        RECT -24.380 2727.380 2944.000 2730.380 ;
        RECT -19.580 2727.370 -16.580 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.200 2727.370 2939.200 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.780 2709.380 2934.400 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -19.580 2550.380 -16.580 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 681.040 2550.380 682.640 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.200 2550.380 2939.200 2550.390 ;
        RECT -24.380 2547.380 2944.000 2550.380 ;
        RECT -19.580 2547.370 -16.580 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 681.040 2547.370 682.640 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.200 2547.370 2939.200 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 681.040 2532.380 682.640 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.780 2529.380 2934.400 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 681.040 2529.370 682.640 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -19.580 2370.380 -16.580 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 681.040 2370.380 682.640 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.200 2370.380 2939.200 2370.390 ;
        RECT -24.380 2367.380 2944.000 2370.380 ;
        RECT -19.580 2367.370 -16.580 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 681.040 2367.370 682.640 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.200 2367.370 2939.200 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 681.040 2352.380 682.640 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.780 2349.380 2934.400 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 681.040 2349.370 682.640 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -19.580 2190.380 -16.580 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 681.040 2190.380 682.640 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.200 2190.380 2939.200 2190.390 ;
        RECT -24.380 2187.380 2944.000 2190.380 ;
        RECT -19.580 2187.370 -16.580 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 681.040 2187.370 682.640 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.200 2187.370 2939.200 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 681.040 2172.380 682.640 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.780 2169.380 2934.400 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 681.040 2169.370 682.640 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -19.580 2010.380 -16.580 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 681.040 2010.380 682.640 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.200 2010.380 2939.200 2010.390 ;
        RECT -24.380 2007.380 2944.000 2010.380 ;
        RECT -19.580 2007.370 -16.580 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 681.040 2007.370 682.640 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.200 2007.370 2939.200 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 681.040 1992.380 682.640 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.780 1989.380 2934.400 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 681.040 1989.370 682.640 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -19.580 1830.380 -16.580 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 681.040 1830.380 682.640 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.200 1830.380 2939.200 1830.390 ;
        RECT -24.380 1827.380 2944.000 1830.380 ;
        RECT -19.580 1827.370 -16.580 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 681.040 1827.370 682.640 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.200 1827.370 2939.200 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 681.040 1812.380 682.640 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.780 1809.380 2934.400 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 681.040 1809.370 682.640 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -19.580 1650.380 -16.580 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 681.040 1650.380 682.640 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.200 1650.380 2939.200 1650.390 ;
        RECT -24.380 1647.380 2944.000 1650.380 ;
        RECT -19.580 1647.370 -16.580 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 681.040 1647.370 682.640 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.200 1647.370 2939.200 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 681.040 1632.380 682.640 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.780 1629.380 2934.400 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 681.040 1629.370 682.640 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -19.580 1470.380 -16.580 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 681.040 1470.380 682.640 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.200 1470.380 2939.200 1470.390 ;
        RECT -24.380 1467.380 2944.000 1470.380 ;
        RECT -19.580 1467.370 -16.580 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 681.040 1467.370 682.640 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.200 1467.370 2939.200 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 681.040 1452.380 682.640 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.780 1449.380 2934.400 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 681.040 1449.370 682.640 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -19.580 1290.380 -16.580 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 681.040 1290.380 682.640 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.200 1290.380 2939.200 1290.390 ;
        RECT -24.380 1287.380 2944.000 1290.380 ;
        RECT -19.580 1287.370 -16.580 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 681.040 1287.370 682.640 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.200 1287.370 2939.200 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 681.040 1272.380 682.640 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.780 1269.380 2934.400 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 681.040 1269.370 682.640 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -19.580 1110.380 -16.580 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 681.040 1110.380 682.640 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.200 1110.380 2939.200 1110.390 ;
        RECT -24.380 1107.380 2944.000 1110.380 ;
        RECT -19.580 1107.370 -16.580 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 681.040 1107.370 682.640 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.200 1107.370 2939.200 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 681.040 1092.380 682.640 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.780 1089.380 2934.400 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 681.040 1089.370 682.640 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -19.580 930.380 -16.580 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.200 930.380 2939.200 930.390 ;
        RECT -24.380 927.380 2944.000 930.380 ;
        RECT -19.580 927.370 -16.580 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.200 927.370 2939.200 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.780 909.380 2934.400 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -19.580 750.380 -16.580 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.200 750.380 2939.200 750.390 ;
        RECT -24.380 747.380 2944.000 750.380 ;
        RECT -19.580 747.370 -16.580 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.200 747.370 2939.200 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.780 729.380 2934.400 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -19.580 570.380 -16.580 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.200 570.380 2939.200 570.390 ;
        RECT -24.380 567.380 2944.000 570.380 ;
        RECT -19.580 567.370 -16.580 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.200 567.370 2939.200 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.780 549.380 2934.400 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -19.580 390.380 -16.580 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.200 390.380 2939.200 390.390 ;
        RECT -24.380 387.380 2944.000 390.380 ;
        RECT -19.580 387.370 -16.580 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.200 387.370 2939.200 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.780 369.380 2934.400 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -19.580 210.380 -16.580 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.200 210.380 2939.200 210.390 ;
        RECT -24.380 207.380 2944.000 210.380 ;
        RECT -19.580 207.370 -16.580 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.200 207.370 2939.200 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.780 189.380 2934.400 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -19.580 30.380 -16.580 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.200 30.380 2939.200 30.390 ;
        RECT -24.380 27.380 2944.000 30.380 ;
        RECT -19.580 27.370 -16.580 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.200 27.370 2939.200 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.780 9.380 2934.400 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.580 -11.220 -16.580 -11.210 ;
        RECT 22.020 -11.220 25.020 -11.210 ;
        RECT 202.020 -11.220 205.020 -11.210 ;
        RECT 382.020 -11.220 385.020 -11.210 ;
        RECT 562.020 -11.220 565.020 -11.210 ;
        RECT 742.020 -11.220 745.020 -11.210 ;
        RECT 922.020 -11.220 925.020 -11.210 ;
        RECT 1102.020 -11.220 1105.020 -11.210 ;
        RECT 1282.020 -11.220 1285.020 -11.210 ;
        RECT 1462.020 -11.220 1465.020 -11.210 ;
        RECT 1642.020 -11.220 1645.020 -11.210 ;
        RECT 1822.020 -11.220 1825.020 -11.210 ;
        RECT 2002.020 -11.220 2005.020 -11.210 ;
        RECT 2182.020 -11.220 2185.020 -11.210 ;
        RECT 2362.020 -11.220 2365.020 -11.210 ;
        RECT 2542.020 -11.220 2545.020 -11.210 ;
        RECT 2722.020 -11.220 2725.020 -11.210 ;
        RECT 2902.020 -11.220 2905.020 -11.210 ;
        RECT 2936.200 -11.220 2939.200 -11.210 ;
        RECT -19.580 -14.220 2939.200 -11.220 ;
        RECT -19.580 -14.230 -16.580 -14.220 ;
        RECT 22.020 -14.230 25.020 -14.220 ;
        RECT 202.020 -14.230 205.020 -14.220 ;
        RECT 382.020 -14.230 385.020 -14.220 ;
        RECT 562.020 -14.230 565.020 -14.220 ;
        RECT 742.020 -14.230 745.020 -14.220 ;
        RECT 922.020 -14.230 925.020 -14.220 ;
        RECT 1102.020 -14.230 1105.020 -14.220 ;
        RECT 1282.020 -14.230 1285.020 -14.220 ;
        RECT 1462.020 -14.230 1465.020 -14.220 ;
        RECT 1642.020 -14.230 1645.020 -14.220 ;
        RECT 1822.020 -14.230 1825.020 -14.220 ;
        RECT 2002.020 -14.230 2005.020 -14.220 ;
        RECT 2182.020 -14.230 2185.020 -14.220 ;
        RECT 2362.020 -14.230 2365.020 -14.220 ;
        RECT 2542.020 -14.230 2545.020 -14.220 ;
        RECT 2722.020 -14.230 2725.020 -14.220 ;
        RECT 2902.020 -14.230 2905.020 -14.220 ;
        RECT 2936.200 -14.230 2939.200 -14.220 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.380 -19.020 -21.380 3538.700 ;
        RECT -14.780 -9.420 -11.780 3529.100 ;
        RECT 94.020 -9.420 97.020 3529.100 ;
        RECT 112.020 -19.020 115.020 3538.700 ;
        RECT 274.020 -9.420 277.020 3529.100 ;
        RECT 292.020 -19.020 295.020 3538.700 ;
        RECT 454.020 -9.420 457.020 3529.100 ;
        RECT 472.020 -19.020 475.020 3538.700 ;
        RECT 634.020 -9.420 637.020 3529.100 ;
        RECT 652.020 -19.020 655.020 3538.700 ;
        RECT 814.020 2562.185 817.020 3529.100 ;
        RECT 832.020 2562.185 835.020 3538.700 ;
        RECT 994.020 2562.185 997.020 3529.100 ;
        RECT 1012.020 2562.185 1015.020 3538.700 ;
        RECT 1174.020 2562.185 1177.020 3529.100 ;
        RECT 1192.020 2562.185 1195.020 3538.700 ;
        RECT 1354.020 2562.185 1357.020 3529.100 ;
        RECT 1372.020 2562.185 1375.020 3538.700 ;
        RECT 1534.020 2562.185 1537.020 3529.100 ;
        RECT 1552.020 2562.185 1555.020 3538.700 ;
        RECT 1714.020 2562.185 1717.020 3529.100 ;
        RECT 1732.020 2562.185 1735.020 3538.700 ;
        RECT 1894.020 2562.185 1897.020 3529.100 ;
        RECT 1912.020 2562.185 1915.020 3538.700 ;
        RECT 2074.020 2562.185 2077.020 3529.100 ;
        RECT 2092.020 2562.185 2095.020 3538.700 ;
        RECT 757.840 970.640 759.440 2551.440 ;
        RECT 814.020 -9.420 817.020 960.000 ;
        RECT 832.020 -19.020 835.020 960.000 ;
        RECT 994.020 -9.420 997.020 960.000 ;
        RECT 1012.020 -19.020 1015.020 960.000 ;
        RECT 1174.020 -9.420 1177.020 960.000 ;
        RECT 1192.020 -19.020 1195.020 960.000 ;
        RECT 1354.020 -9.420 1357.020 960.000 ;
        RECT 1372.020 -19.020 1375.020 960.000 ;
        RECT 1534.020 -9.420 1537.020 960.000 ;
        RECT 1552.020 -19.020 1555.020 960.000 ;
        RECT 1714.020 -9.420 1717.020 960.000 ;
        RECT 1732.020 -19.020 1735.020 960.000 ;
        RECT 1894.020 -9.420 1897.020 960.000 ;
        RECT 1912.020 -19.020 1915.020 960.000 ;
        RECT 2074.020 -9.420 2077.020 960.000 ;
        RECT 2092.020 -19.020 2095.020 960.000 ;
        RECT 2254.020 -9.420 2257.020 3529.100 ;
        RECT 2272.020 -19.020 2275.020 3538.700 ;
        RECT 2434.020 -9.420 2437.020 3529.100 ;
        RECT 2452.020 -19.020 2455.020 3538.700 ;
        RECT 2614.020 -9.420 2617.020 3529.100 ;
        RECT 2632.020 -19.020 2635.020 3538.700 ;
        RECT 2794.020 -9.420 2797.020 3529.100 ;
        RECT 2812.020 -19.020 2815.020 3538.700 ;
        RECT 2931.400 -9.420 2934.400 3529.100 ;
        RECT 2941.000 -19.020 2944.000 3538.700 ;
      LAYER via4 ;
        RECT -23.470 3537.410 -22.290 3538.590 ;
        RECT -23.470 3535.810 -22.290 3536.990 ;
        RECT 112.930 3537.410 114.110 3538.590 ;
        RECT 112.930 3535.810 114.110 3536.990 ;
        RECT -23.470 3359.090 -22.290 3360.270 ;
        RECT -23.470 3357.490 -22.290 3358.670 ;
        RECT -23.470 3179.090 -22.290 3180.270 ;
        RECT -23.470 3177.490 -22.290 3178.670 ;
        RECT -23.470 2999.090 -22.290 3000.270 ;
        RECT -23.470 2997.490 -22.290 2998.670 ;
        RECT -23.470 2819.090 -22.290 2820.270 ;
        RECT -23.470 2817.490 -22.290 2818.670 ;
        RECT -23.470 2639.090 -22.290 2640.270 ;
        RECT -23.470 2637.490 -22.290 2638.670 ;
        RECT -23.470 2459.090 -22.290 2460.270 ;
        RECT -23.470 2457.490 -22.290 2458.670 ;
        RECT -23.470 2279.090 -22.290 2280.270 ;
        RECT -23.470 2277.490 -22.290 2278.670 ;
        RECT -23.470 2099.090 -22.290 2100.270 ;
        RECT -23.470 2097.490 -22.290 2098.670 ;
        RECT -23.470 1919.090 -22.290 1920.270 ;
        RECT -23.470 1917.490 -22.290 1918.670 ;
        RECT -23.470 1739.090 -22.290 1740.270 ;
        RECT -23.470 1737.490 -22.290 1738.670 ;
        RECT -23.470 1559.090 -22.290 1560.270 ;
        RECT -23.470 1557.490 -22.290 1558.670 ;
        RECT -23.470 1379.090 -22.290 1380.270 ;
        RECT -23.470 1377.490 -22.290 1378.670 ;
        RECT -23.470 1199.090 -22.290 1200.270 ;
        RECT -23.470 1197.490 -22.290 1198.670 ;
        RECT -23.470 1019.090 -22.290 1020.270 ;
        RECT -23.470 1017.490 -22.290 1018.670 ;
        RECT -23.470 839.090 -22.290 840.270 ;
        RECT -23.470 837.490 -22.290 838.670 ;
        RECT -23.470 659.090 -22.290 660.270 ;
        RECT -23.470 657.490 -22.290 658.670 ;
        RECT -23.470 479.090 -22.290 480.270 ;
        RECT -23.470 477.490 -22.290 478.670 ;
        RECT -23.470 299.090 -22.290 300.270 ;
        RECT -23.470 297.490 -22.290 298.670 ;
        RECT -23.470 119.090 -22.290 120.270 ;
        RECT -23.470 117.490 -22.290 118.670 ;
        RECT -13.870 3527.810 -12.690 3528.990 ;
        RECT -13.870 3526.210 -12.690 3527.390 ;
        RECT -13.870 3341.090 -12.690 3342.270 ;
        RECT -13.870 3339.490 -12.690 3340.670 ;
        RECT -13.870 3161.090 -12.690 3162.270 ;
        RECT -13.870 3159.490 -12.690 3160.670 ;
        RECT -13.870 2981.090 -12.690 2982.270 ;
        RECT -13.870 2979.490 -12.690 2980.670 ;
        RECT -13.870 2801.090 -12.690 2802.270 ;
        RECT -13.870 2799.490 -12.690 2800.670 ;
        RECT -13.870 2621.090 -12.690 2622.270 ;
        RECT -13.870 2619.490 -12.690 2620.670 ;
        RECT -13.870 2441.090 -12.690 2442.270 ;
        RECT -13.870 2439.490 -12.690 2440.670 ;
        RECT -13.870 2261.090 -12.690 2262.270 ;
        RECT -13.870 2259.490 -12.690 2260.670 ;
        RECT -13.870 2081.090 -12.690 2082.270 ;
        RECT -13.870 2079.490 -12.690 2080.670 ;
        RECT -13.870 1901.090 -12.690 1902.270 ;
        RECT -13.870 1899.490 -12.690 1900.670 ;
        RECT -13.870 1721.090 -12.690 1722.270 ;
        RECT -13.870 1719.490 -12.690 1720.670 ;
        RECT -13.870 1541.090 -12.690 1542.270 ;
        RECT -13.870 1539.490 -12.690 1540.670 ;
        RECT -13.870 1361.090 -12.690 1362.270 ;
        RECT -13.870 1359.490 -12.690 1360.670 ;
        RECT -13.870 1181.090 -12.690 1182.270 ;
        RECT -13.870 1179.490 -12.690 1180.670 ;
        RECT -13.870 1001.090 -12.690 1002.270 ;
        RECT -13.870 999.490 -12.690 1000.670 ;
        RECT -13.870 821.090 -12.690 822.270 ;
        RECT -13.870 819.490 -12.690 820.670 ;
        RECT -13.870 641.090 -12.690 642.270 ;
        RECT -13.870 639.490 -12.690 640.670 ;
        RECT -13.870 461.090 -12.690 462.270 ;
        RECT -13.870 459.490 -12.690 460.670 ;
        RECT -13.870 281.090 -12.690 282.270 ;
        RECT -13.870 279.490 -12.690 280.670 ;
        RECT -13.870 101.090 -12.690 102.270 ;
        RECT -13.870 99.490 -12.690 100.670 ;
        RECT -13.870 -7.710 -12.690 -6.530 ;
        RECT -13.870 -9.310 -12.690 -8.130 ;
        RECT 94.930 3527.810 96.110 3528.990 ;
        RECT 94.930 3526.210 96.110 3527.390 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.710 96.110 -6.530 ;
        RECT 94.930 -9.310 96.110 -8.130 ;
        RECT 292.930 3537.410 294.110 3538.590 ;
        RECT 292.930 3535.810 294.110 3536.990 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.470 -17.310 -22.290 -16.130 ;
        RECT -23.470 -18.910 -22.290 -17.730 ;
        RECT 274.930 3527.810 276.110 3528.990 ;
        RECT 274.930 3526.210 276.110 3527.390 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.710 276.110 -6.530 ;
        RECT 274.930 -9.310 276.110 -8.130 ;
        RECT 472.930 3537.410 474.110 3538.590 ;
        RECT 472.930 3535.810 474.110 3536.990 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 112.930 -17.310 114.110 -16.130 ;
        RECT 112.930 -18.910 114.110 -17.730 ;
        RECT 454.930 3527.810 456.110 3528.990 ;
        RECT 454.930 3526.210 456.110 3527.390 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.710 456.110 -6.530 ;
        RECT 454.930 -9.310 456.110 -8.130 ;
        RECT 652.930 3537.410 654.110 3538.590 ;
        RECT 652.930 3535.810 654.110 3536.990 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 292.930 -17.310 294.110 -16.130 ;
        RECT 292.930 -18.910 294.110 -17.730 ;
        RECT 634.930 3527.810 636.110 3528.990 ;
        RECT 634.930 3526.210 636.110 3527.390 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.710 636.110 -6.530 ;
        RECT 634.930 -9.310 636.110 -8.130 ;
        RECT 832.930 3537.410 834.110 3538.590 ;
        RECT 832.930 3535.810 834.110 3536.990 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 814.930 3527.810 816.110 3528.990 ;
        RECT 814.930 3526.210 816.110 3527.390 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 1012.930 3537.410 1014.110 3538.590 ;
        RECT 1012.930 3535.810 1014.110 3536.990 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 994.930 3527.810 996.110 3528.990 ;
        RECT 994.930 3526.210 996.110 3527.390 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 1192.930 3537.410 1194.110 3538.590 ;
        RECT 1192.930 3535.810 1194.110 3536.990 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1174.930 3527.810 1176.110 3528.990 ;
        RECT 1174.930 3526.210 1176.110 3527.390 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1372.930 3537.410 1374.110 3538.590 ;
        RECT 1372.930 3535.810 1374.110 3536.990 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1354.930 3527.810 1356.110 3528.990 ;
        RECT 1354.930 3526.210 1356.110 3527.390 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1552.930 3537.410 1554.110 3538.590 ;
        RECT 1552.930 3535.810 1554.110 3536.990 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1534.930 3527.810 1536.110 3528.990 ;
        RECT 1534.930 3526.210 1536.110 3527.390 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1732.930 3537.410 1734.110 3538.590 ;
        RECT 1732.930 3535.810 1734.110 3536.990 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1714.930 3527.810 1716.110 3528.990 ;
        RECT 1714.930 3526.210 1716.110 3527.390 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1912.930 3537.410 1914.110 3538.590 ;
        RECT 1912.930 3535.810 1914.110 3536.990 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1894.930 3527.810 1896.110 3528.990 ;
        RECT 1894.930 3526.210 1896.110 3527.390 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 2092.930 3537.410 2094.110 3538.590 ;
        RECT 2092.930 3535.810 2094.110 3536.990 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 2074.930 3527.810 2076.110 3528.990 ;
        RECT 2074.930 3526.210 2076.110 3527.390 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2272.930 3537.410 2274.110 3538.590 ;
        RECT 2272.930 3535.810 2274.110 3536.990 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2254.930 3527.810 2256.110 3528.990 ;
        RECT 2254.930 3526.210 2256.110 3527.390 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 758.050 2459.090 759.230 2460.270 ;
        RECT 758.050 2457.490 759.230 2458.670 ;
        RECT 758.050 2441.090 759.230 2442.270 ;
        RECT 758.050 2439.490 759.230 2440.670 ;
        RECT 758.050 2279.090 759.230 2280.270 ;
        RECT 758.050 2277.490 759.230 2278.670 ;
        RECT 758.050 2261.090 759.230 2262.270 ;
        RECT 758.050 2259.490 759.230 2260.670 ;
        RECT 758.050 2099.090 759.230 2100.270 ;
        RECT 758.050 2097.490 759.230 2098.670 ;
        RECT 758.050 2081.090 759.230 2082.270 ;
        RECT 758.050 2079.490 759.230 2080.670 ;
        RECT 758.050 1919.090 759.230 1920.270 ;
        RECT 758.050 1917.490 759.230 1918.670 ;
        RECT 758.050 1901.090 759.230 1902.270 ;
        RECT 758.050 1899.490 759.230 1900.670 ;
        RECT 758.050 1739.090 759.230 1740.270 ;
        RECT 758.050 1737.490 759.230 1738.670 ;
        RECT 758.050 1721.090 759.230 1722.270 ;
        RECT 758.050 1719.490 759.230 1720.670 ;
        RECT 758.050 1559.090 759.230 1560.270 ;
        RECT 758.050 1557.490 759.230 1558.670 ;
        RECT 758.050 1541.090 759.230 1542.270 ;
        RECT 758.050 1539.490 759.230 1540.670 ;
        RECT 758.050 1379.090 759.230 1380.270 ;
        RECT 758.050 1377.490 759.230 1378.670 ;
        RECT 758.050 1361.090 759.230 1362.270 ;
        RECT 758.050 1359.490 759.230 1360.670 ;
        RECT 758.050 1199.090 759.230 1200.270 ;
        RECT 758.050 1197.490 759.230 1198.670 ;
        RECT 758.050 1181.090 759.230 1182.270 ;
        RECT 758.050 1179.490 759.230 1180.670 ;
        RECT 758.050 1019.090 759.230 1020.270 ;
        RECT 758.050 1017.490 759.230 1018.670 ;
        RECT 758.050 1001.090 759.230 1002.270 ;
        RECT 758.050 999.490 759.230 1000.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 472.930 -17.310 474.110 -16.130 ;
        RECT 472.930 -18.910 474.110 -17.730 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.710 816.110 -6.530 ;
        RECT 814.930 -9.310 816.110 -8.130 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 652.930 -17.310 654.110 -16.130 ;
        RECT 652.930 -18.910 654.110 -17.730 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.710 996.110 -6.530 ;
        RECT 994.930 -9.310 996.110 -8.130 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 832.930 -17.310 834.110 -16.130 ;
        RECT 832.930 -18.910 834.110 -17.730 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.710 1176.110 -6.530 ;
        RECT 1174.930 -9.310 1176.110 -8.130 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1012.930 -17.310 1014.110 -16.130 ;
        RECT 1012.930 -18.910 1014.110 -17.730 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.710 1356.110 -6.530 ;
        RECT 1354.930 -9.310 1356.110 -8.130 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1192.930 -17.310 1194.110 -16.130 ;
        RECT 1192.930 -18.910 1194.110 -17.730 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.710 1536.110 -6.530 ;
        RECT 1534.930 -9.310 1536.110 -8.130 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1372.930 -17.310 1374.110 -16.130 ;
        RECT 1372.930 -18.910 1374.110 -17.730 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.710 1716.110 -6.530 ;
        RECT 1714.930 -9.310 1716.110 -8.130 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1552.930 -17.310 1554.110 -16.130 ;
        RECT 1552.930 -18.910 1554.110 -17.730 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.710 1896.110 -6.530 ;
        RECT 1894.930 -9.310 1896.110 -8.130 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1732.930 -17.310 1734.110 -16.130 ;
        RECT 1732.930 -18.910 1734.110 -17.730 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.710 2076.110 -6.530 ;
        RECT 2074.930 -9.310 2076.110 -8.130 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 1912.930 -17.310 1914.110 -16.130 ;
        RECT 1912.930 -18.910 1914.110 -17.730 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.710 2256.110 -6.530 ;
        RECT 2254.930 -9.310 2256.110 -8.130 ;
        RECT 2452.930 3537.410 2454.110 3538.590 ;
        RECT 2452.930 3535.810 2454.110 3536.990 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2092.930 -17.310 2094.110 -16.130 ;
        RECT 2092.930 -18.910 2094.110 -17.730 ;
        RECT 2434.930 3527.810 2436.110 3528.990 ;
        RECT 2434.930 3526.210 2436.110 3527.390 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.710 2436.110 -6.530 ;
        RECT 2434.930 -9.310 2436.110 -8.130 ;
        RECT 2632.930 3537.410 2634.110 3538.590 ;
        RECT 2632.930 3535.810 2634.110 3536.990 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2272.930 -17.310 2274.110 -16.130 ;
        RECT 2272.930 -18.910 2274.110 -17.730 ;
        RECT 2614.930 3527.810 2616.110 3528.990 ;
        RECT 2614.930 3526.210 2616.110 3527.390 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.710 2616.110 -6.530 ;
        RECT 2614.930 -9.310 2616.110 -8.130 ;
        RECT 2812.930 3537.410 2814.110 3538.590 ;
        RECT 2812.930 3535.810 2814.110 3536.990 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2452.930 -17.310 2454.110 -16.130 ;
        RECT 2452.930 -18.910 2454.110 -17.730 ;
        RECT 2794.930 3527.810 2796.110 3528.990 ;
        RECT 2794.930 3526.210 2796.110 3527.390 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.710 2796.110 -6.530 ;
        RECT 2794.930 -9.310 2796.110 -8.130 ;
        RECT 2941.910 3537.410 2943.090 3538.590 ;
        RECT 2941.910 3535.810 2943.090 3536.990 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2632.930 -17.310 2634.110 -16.130 ;
        RECT 2632.930 -18.910 2634.110 -17.730 ;
        RECT 2932.310 3527.810 2933.490 3528.990 ;
        RECT 2932.310 3526.210 2933.490 3527.390 ;
        RECT 2932.310 3341.090 2933.490 3342.270 ;
        RECT 2932.310 3339.490 2933.490 3340.670 ;
        RECT 2932.310 3161.090 2933.490 3162.270 ;
        RECT 2932.310 3159.490 2933.490 3160.670 ;
        RECT 2932.310 2981.090 2933.490 2982.270 ;
        RECT 2932.310 2979.490 2933.490 2980.670 ;
        RECT 2932.310 2801.090 2933.490 2802.270 ;
        RECT 2932.310 2799.490 2933.490 2800.670 ;
        RECT 2932.310 2621.090 2933.490 2622.270 ;
        RECT 2932.310 2619.490 2933.490 2620.670 ;
        RECT 2932.310 2441.090 2933.490 2442.270 ;
        RECT 2932.310 2439.490 2933.490 2440.670 ;
        RECT 2932.310 2261.090 2933.490 2262.270 ;
        RECT 2932.310 2259.490 2933.490 2260.670 ;
        RECT 2932.310 2081.090 2933.490 2082.270 ;
        RECT 2932.310 2079.490 2933.490 2080.670 ;
        RECT 2932.310 1901.090 2933.490 1902.270 ;
        RECT 2932.310 1899.490 2933.490 1900.670 ;
        RECT 2932.310 1721.090 2933.490 1722.270 ;
        RECT 2932.310 1719.490 2933.490 1720.670 ;
        RECT 2932.310 1541.090 2933.490 1542.270 ;
        RECT 2932.310 1539.490 2933.490 1540.670 ;
        RECT 2932.310 1361.090 2933.490 1362.270 ;
        RECT 2932.310 1359.490 2933.490 1360.670 ;
        RECT 2932.310 1181.090 2933.490 1182.270 ;
        RECT 2932.310 1179.490 2933.490 1180.670 ;
        RECT 2932.310 1001.090 2933.490 1002.270 ;
        RECT 2932.310 999.490 2933.490 1000.670 ;
        RECT 2932.310 821.090 2933.490 822.270 ;
        RECT 2932.310 819.490 2933.490 820.670 ;
        RECT 2932.310 641.090 2933.490 642.270 ;
        RECT 2932.310 639.490 2933.490 640.670 ;
        RECT 2932.310 461.090 2933.490 462.270 ;
        RECT 2932.310 459.490 2933.490 460.670 ;
        RECT 2932.310 281.090 2933.490 282.270 ;
        RECT 2932.310 279.490 2933.490 280.670 ;
        RECT 2932.310 101.090 2933.490 102.270 ;
        RECT 2932.310 99.490 2933.490 100.670 ;
        RECT 2932.310 -7.710 2933.490 -6.530 ;
        RECT 2932.310 -9.310 2933.490 -8.130 ;
        RECT 2941.910 3359.090 2943.090 3360.270 ;
        RECT 2941.910 3357.490 2943.090 3358.670 ;
        RECT 2941.910 3179.090 2943.090 3180.270 ;
        RECT 2941.910 3177.490 2943.090 3178.670 ;
        RECT 2941.910 2999.090 2943.090 3000.270 ;
        RECT 2941.910 2997.490 2943.090 2998.670 ;
        RECT 2941.910 2819.090 2943.090 2820.270 ;
        RECT 2941.910 2817.490 2943.090 2818.670 ;
        RECT 2941.910 2639.090 2943.090 2640.270 ;
        RECT 2941.910 2637.490 2943.090 2638.670 ;
        RECT 2941.910 2459.090 2943.090 2460.270 ;
        RECT 2941.910 2457.490 2943.090 2458.670 ;
        RECT 2941.910 2279.090 2943.090 2280.270 ;
        RECT 2941.910 2277.490 2943.090 2278.670 ;
        RECT 2941.910 2099.090 2943.090 2100.270 ;
        RECT 2941.910 2097.490 2943.090 2098.670 ;
        RECT 2941.910 1919.090 2943.090 1920.270 ;
        RECT 2941.910 1917.490 2943.090 1918.670 ;
        RECT 2941.910 1739.090 2943.090 1740.270 ;
        RECT 2941.910 1737.490 2943.090 1738.670 ;
        RECT 2941.910 1559.090 2943.090 1560.270 ;
        RECT 2941.910 1557.490 2943.090 1558.670 ;
        RECT 2941.910 1379.090 2943.090 1380.270 ;
        RECT 2941.910 1377.490 2943.090 1378.670 ;
        RECT 2941.910 1199.090 2943.090 1200.270 ;
        RECT 2941.910 1197.490 2943.090 1198.670 ;
        RECT 2941.910 1019.090 2943.090 1020.270 ;
        RECT 2941.910 1017.490 2943.090 1018.670 ;
        RECT 2941.910 839.090 2943.090 840.270 ;
        RECT 2941.910 837.490 2943.090 838.670 ;
        RECT 2941.910 659.090 2943.090 660.270 ;
        RECT 2941.910 657.490 2943.090 658.670 ;
        RECT 2941.910 479.090 2943.090 480.270 ;
        RECT 2941.910 477.490 2943.090 478.670 ;
        RECT 2941.910 299.090 2943.090 300.270 ;
        RECT 2941.910 297.490 2943.090 298.670 ;
        RECT 2941.910 119.090 2943.090 120.270 ;
        RECT 2941.910 117.490 2943.090 118.670 ;
        RECT 2812.930 -17.310 2814.110 -16.130 ;
        RECT 2812.930 -18.910 2814.110 -17.730 ;
        RECT 2941.910 -17.310 2943.090 -16.130 ;
        RECT 2941.910 -18.910 2943.090 -17.730 ;
      LAYER met5 ;
        RECT -24.380 3538.700 -21.380 3538.710 ;
        RECT 112.020 3538.700 115.020 3538.710 ;
        RECT 292.020 3538.700 295.020 3538.710 ;
        RECT 472.020 3538.700 475.020 3538.710 ;
        RECT 652.020 3538.700 655.020 3538.710 ;
        RECT 832.020 3538.700 835.020 3538.710 ;
        RECT 1012.020 3538.700 1015.020 3538.710 ;
        RECT 1192.020 3538.700 1195.020 3538.710 ;
        RECT 1372.020 3538.700 1375.020 3538.710 ;
        RECT 1552.020 3538.700 1555.020 3538.710 ;
        RECT 1732.020 3538.700 1735.020 3538.710 ;
        RECT 1912.020 3538.700 1915.020 3538.710 ;
        RECT 2092.020 3538.700 2095.020 3538.710 ;
        RECT 2272.020 3538.700 2275.020 3538.710 ;
        RECT 2452.020 3538.700 2455.020 3538.710 ;
        RECT 2632.020 3538.700 2635.020 3538.710 ;
        RECT 2812.020 3538.700 2815.020 3538.710 ;
        RECT 2941.000 3538.700 2944.000 3538.710 ;
        RECT -24.380 3535.700 2944.000 3538.700 ;
        RECT -24.380 3535.690 -21.380 3535.700 ;
        RECT 112.020 3535.690 115.020 3535.700 ;
        RECT 292.020 3535.690 295.020 3535.700 ;
        RECT 472.020 3535.690 475.020 3535.700 ;
        RECT 652.020 3535.690 655.020 3535.700 ;
        RECT 832.020 3535.690 835.020 3535.700 ;
        RECT 1012.020 3535.690 1015.020 3535.700 ;
        RECT 1192.020 3535.690 1195.020 3535.700 ;
        RECT 1372.020 3535.690 1375.020 3535.700 ;
        RECT 1552.020 3535.690 1555.020 3535.700 ;
        RECT 1732.020 3535.690 1735.020 3535.700 ;
        RECT 1912.020 3535.690 1915.020 3535.700 ;
        RECT 2092.020 3535.690 2095.020 3535.700 ;
        RECT 2272.020 3535.690 2275.020 3535.700 ;
        RECT 2452.020 3535.690 2455.020 3535.700 ;
        RECT 2632.020 3535.690 2635.020 3535.700 ;
        RECT 2812.020 3535.690 2815.020 3535.700 ;
        RECT 2941.000 3535.690 2944.000 3535.700 ;
        RECT -14.780 3529.100 -11.780 3529.110 ;
        RECT 94.020 3529.100 97.020 3529.110 ;
        RECT 274.020 3529.100 277.020 3529.110 ;
        RECT 454.020 3529.100 457.020 3529.110 ;
        RECT 634.020 3529.100 637.020 3529.110 ;
        RECT 814.020 3529.100 817.020 3529.110 ;
        RECT 994.020 3529.100 997.020 3529.110 ;
        RECT 1174.020 3529.100 1177.020 3529.110 ;
        RECT 1354.020 3529.100 1357.020 3529.110 ;
        RECT 1534.020 3529.100 1537.020 3529.110 ;
        RECT 1714.020 3529.100 1717.020 3529.110 ;
        RECT 1894.020 3529.100 1897.020 3529.110 ;
        RECT 2074.020 3529.100 2077.020 3529.110 ;
        RECT 2254.020 3529.100 2257.020 3529.110 ;
        RECT 2434.020 3529.100 2437.020 3529.110 ;
        RECT 2614.020 3529.100 2617.020 3529.110 ;
        RECT 2794.020 3529.100 2797.020 3529.110 ;
        RECT 2931.400 3529.100 2934.400 3529.110 ;
        RECT -14.780 3526.100 2934.400 3529.100 ;
        RECT -14.780 3526.090 -11.780 3526.100 ;
        RECT 94.020 3526.090 97.020 3526.100 ;
        RECT 274.020 3526.090 277.020 3526.100 ;
        RECT 454.020 3526.090 457.020 3526.100 ;
        RECT 634.020 3526.090 637.020 3526.100 ;
        RECT 814.020 3526.090 817.020 3526.100 ;
        RECT 994.020 3526.090 997.020 3526.100 ;
        RECT 1174.020 3526.090 1177.020 3526.100 ;
        RECT 1354.020 3526.090 1357.020 3526.100 ;
        RECT 1534.020 3526.090 1537.020 3526.100 ;
        RECT 1714.020 3526.090 1717.020 3526.100 ;
        RECT 1894.020 3526.090 1897.020 3526.100 ;
        RECT 2074.020 3526.090 2077.020 3526.100 ;
        RECT 2254.020 3526.090 2257.020 3526.100 ;
        RECT 2434.020 3526.090 2437.020 3526.100 ;
        RECT 2614.020 3526.090 2617.020 3526.100 ;
        RECT 2794.020 3526.090 2797.020 3526.100 ;
        RECT 2931.400 3526.090 2934.400 3526.100 ;
        RECT -24.380 3360.380 -21.380 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2941.000 3360.380 2944.000 3360.390 ;
        RECT -24.380 3357.380 2944.000 3360.380 ;
        RECT -24.380 3357.370 -21.380 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2941.000 3357.370 2944.000 3357.380 ;
        RECT -14.780 3342.380 -11.780 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.400 3342.380 2934.400 3342.390 ;
        RECT -14.780 3339.380 2934.400 3342.380 ;
        RECT -14.780 3339.370 -11.780 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.400 3339.370 2934.400 3339.380 ;
        RECT -24.380 3180.380 -21.380 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2941.000 3180.380 2944.000 3180.390 ;
        RECT -24.380 3177.380 2944.000 3180.380 ;
        RECT -24.380 3177.370 -21.380 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2941.000 3177.370 2944.000 3177.380 ;
        RECT -14.780 3162.380 -11.780 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.400 3162.380 2934.400 3162.390 ;
        RECT -14.780 3159.380 2934.400 3162.380 ;
        RECT -14.780 3159.370 -11.780 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.400 3159.370 2934.400 3159.380 ;
        RECT -24.380 3000.380 -21.380 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2941.000 3000.380 2944.000 3000.390 ;
        RECT -24.380 2997.380 2944.000 3000.380 ;
        RECT -24.380 2997.370 -21.380 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2941.000 2997.370 2944.000 2997.380 ;
        RECT -14.780 2982.380 -11.780 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.400 2982.380 2934.400 2982.390 ;
        RECT -14.780 2979.380 2934.400 2982.380 ;
        RECT -14.780 2979.370 -11.780 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.400 2979.370 2934.400 2979.380 ;
        RECT -24.380 2820.380 -21.380 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2941.000 2820.380 2944.000 2820.390 ;
        RECT -24.380 2817.380 2944.000 2820.380 ;
        RECT -24.380 2817.370 -21.380 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2941.000 2817.370 2944.000 2817.380 ;
        RECT -14.780 2802.380 -11.780 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.400 2802.380 2934.400 2802.390 ;
        RECT -14.780 2799.380 2934.400 2802.380 ;
        RECT -14.780 2799.370 -11.780 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.400 2799.370 2934.400 2799.380 ;
        RECT -24.380 2640.380 -21.380 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2941.000 2640.380 2944.000 2640.390 ;
        RECT -24.380 2637.380 2944.000 2640.380 ;
        RECT -24.380 2637.370 -21.380 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2941.000 2637.370 2944.000 2637.380 ;
        RECT -14.780 2622.380 -11.780 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.400 2622.380 2934.400 2622.390 ;
        RECT -14.780 2619.380 2934.400 2622.380 ;
        RECT -14.780 2619.370 -11.780 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.400 2619.370 2934.400 2619.380 ;
        RECT -24.380 2460.380 -21.380 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 757.840 2460.380 759.440 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2941.000 2460.380 2944.000 2460.390 ;
        RECT -24.380 2457.380 2944.000 2460.380 ;
        RECT -24.380 2457.370 -21.380 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 757.840 2457.370 759.440 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2941.000 2457.370 2944.000 2457.380 ;
        RECT -14.780 2442.380 -11.780 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 757.840 2442.380 759.440 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.400 2442.380 2934.400 2442.390 ;
        RECT -14.780 2439.380 2934.400 2442.380 ;
        RECT -14.780 2439.370 -11.780 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 757.840 2439.370 759.440 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.400 2439.370 2934.400 2439.380 ;
        RECT -24.380 2280.380 -21.380 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 757.840 2280.380 759.440 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2941.000 2280.380 2944.000 2280.390 ;
        RECT -24.380 2277.380 2944.000 2280.380 ;
        RECT -24.380 2277.370 -21.380 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 757.840 2277.370 759.440 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2941.000 2277.370 2944.000 2277.380 ;
        RECT -14.780 2262.380 -11.780 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 757.840 2262.380 759.440 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.400 2262.380 2934.400 2262.390 ;
        RECT -14.780 2259.380 2934.400 2262.380 ;
        RECT -14.780 2259.370 -11.780 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 757.840 2259.370 759.440 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.400 2259.370 2934.400 2259.380 ;
        RECT -24.380 2100.380 -21.380 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 757.840 2100.380 759.440 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2941.000 2100.380 2944.000 2100.390 ;
        RECT -24.380 2097.380 2944.000 2100.380 ;
        RECT -24.380 2097.370 -21.380 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 757.840 2097.370 759.440 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2941.000 2097.370 2944.000 2097.380 ;
        RECT -14.780 2082.380 -11.780 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 757.840 2082.380 759.440 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.400 2082.380 2934.400 2082.390 ;
        RECT -14.780 2079.380 2934.400 2082.380 ;
        RECT -14.780 2079.370 -11.780 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 757.840 2079.370 759.440 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.400 2079.370 2934.400 2079.380 ;
        RECT -24.380 1920.380 -21.380 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 757.840 1920.380 759.440 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2941.000 1920.380 2944.000 1920.390 ;
        RECT -24.380 1917.380 2944.000 1920.380 ;
        RECT -24.380 1917.370 -21.380 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 757.840 1917.370 759.440 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2941.000 1917.370 2944.000 1917.380 ;
        RECT -14.780 1902.380 -11.780 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 757.840 1902.380 759.440 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.400 1902.380 2934.400 1902.390 ;
        RECT -14.780 1899.380 2934.400 1902.380 ;
        RECT -14.780 1899.370 -11.780 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 757.840 1899.370 759.440 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.400 1899.370 2934.400 1899.380 ;
        RECT -24.380 1740.380 -21.380 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 757.840 1740.380 759.440 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2941.000 1740.380 2944.000 1740.390 ;
        RECT -24.380 1737.380 2944.000 1740.380 ;
        RECT -24.380 1737.370 -21.380 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 757.840 1737.370 759.440 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2941.000 1737.370 2944.000 1737.380 ;
        RECT -14.780 1722.380 -11.780 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 757.840 1722.380 759.440 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.400 1722.380 2934.400 1722.390 ;
        RECT -14.780 1719.380 2934.400 1722.380 ;
        RECT -14.780 1719.370 -11.780 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 757.840 1719.370 759.440 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.400 1719.370 2934.400 1719.380 ;
        RECT -24.380 1560.380 -21.380 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 757.840 1560.380 759.440 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2941.000 1560.380 2944.000 1560.390 ;
        RECT -24.380 1557.380 2944.000 1560.380 ;
        RECT -24.380 1557.370 -21.380 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 757.840 1557.370 759.440 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2941.000 1557.370 2944.000 1557.380 ;
        RECT -14.780 1542.380 -11.780 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 757.840 1542.380 759.440 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.400 1542.380 2934.400 1542.390 ;
        RECT -14.780 1539.380 2934.400 1542.380 ;
        RECT -14.780 1539.370 -11.780 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 757.840 1539.370 759.440 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.400 1539.370 2934.400 1539.380 ;
        RECT -24.380 1380.380 -21.380 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 757.840 1380.380 759.440 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2941.000 1380.380 2944.000 1380.390 ;
        RECT -24.380 1377.380 2944.000 1380.380 ;
        RECT -24.380 1377.370 -21.380 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 757.840 1377.370 759.440 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2941.000 1377.370 2944.000 1377.380 ;
        RECT -14.780 1362.380 -11.780 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 757.840 1362.380 759.440 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.400 1362.380 2934.400 1362.390 ;
        RECT -14.780 1359.380 2934.400 1362.380 ;
        RECT -14.780 1359.370 -11.780 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 757.840 1359.370 759.440 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.400 1359.370 2934.400 1359.380 ;
        RECT -24.380 1200.380 -21.380 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 757.840 1200.380 759.440 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2941.000 1200.380 2944.000 1200.390 ;
        RECT -24.380 1197.380 2944.000 1200.380 ;
        RECT -24.380 1197.370 -21.380 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 757.840 1197.370 759.440 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2941.000 1197.370 2944.000 1197.380 ;
        RECT -14.780 1182.380 -11.780 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 757.840 1182.380 759.440 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.400 1182.380 2934.400 1182.390 ;
        RECT -14.780 1179.380 2934.400 1182.380 ;
        RECT -14.780 1179.370 -11.780 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 757.840 1179.370 759.440 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.400 1179.370 2934.400 1179.380 ;
        RECT -24.380 1020.380 -21.380 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 757.840 1020.380 759.440 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2941.000 1020.380 2944.000 1020.390 ;
        RECT -24.380 1017.380 2944.000 1020.380 ;
        RECT -24.380 1017.370 -21.380 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 757.840 1017.370 759.440 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2941.000 1017.370 2944.000 1017.380 ;
        RECT -14.780 1002.380 -11.780 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 757.840 1002.380 759.440 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.400 1002.380 2934.400 1002.390 ;
        RECT -14.780 999.380 2934.400 1002.380 ;
        RECT -14.780 999.370 -11.780 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 757.840 999.370 759.440 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.400 999.370 2934.400 999.380 ;
        RECT -24.380 840.380 -21.380 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2941.000 840.380 2944.000 840.390 ;
        RECT -24.380 837.380 2944.000 840.380 ;
        RECT -24.380 837.370 -21.380 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2941.000 837.370 2944.000 837.380 ;
        RECT -14.780 822.380 -11.780 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.400 822.380 2934.400 822.390 ;
        RECT -14.780 819.380 2934.400 822.380 ;
        RECT -14.780 819.370 -11.780 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.400 819.370 2934.400 819.380 ;
        RECT -24.380 660.380 -21.380 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2941.000 660.380 2944.000 660.390 ;
        RECT -24.380 657.380 2944.000 660.380 ;
        RECT -24.380 657.370 -21.380 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2941.000 657.370 2944.000 657.380 ;
        RECT -14.780 642.380 -11.780 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.400 642.380 2934.400 642.390 ;
        RECT -14.780 639.380 2934.400 642.380 ;
        RECT -14.780 639.370 -11.780 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.400 639.370 2934.400 639.380 ;
        RECT -24.380 480.380 -21.380 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2941.000 480.380 2944.000 480.390 ;
        RECT -24.380 477.380 2944.000 480.380 ;
        RECT -24.380 477.370 -21.380 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2941.000 477.370 2944.000 477.380 ;
        RECT -14.780 462.380 -11.780 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.400 462.380 2934.400 462.390 ;
        RECT -14.780 459.380 2934.400 462.380 ;
        RECT -14.780 459.370 -11.780 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.400 459.370 2934.400 459.380 ;
        RECT -24.380 300.380 -21.380 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2941.000 300.380 2944.000 300.390 ;
        RECT -24.380 297.380 2944.000 300.380 ;
        RECT -24.380 297.370 -21.380 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2941.000 297.370 2944.000 297.380 ;
        RECT -14.780 282.380 -11.780 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.400 282.380 2934.400 282.390 ;
        RECT -14.780 279.380 2934.400 282.380 ;
        RECT -14.780 279.370 -11.780 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.400 279.370 2934.400 279.380 ;
        RECT -24.380 120.380 -21.380 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2941.000 120.380 2944.000 120.390 ;
        RECT -24.380 117.380 2944.000 120.380 ;
        RECT -24.380 117.370 -21.380 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2941.000 117.370 2944.000 117.380 ;
        RECT -14.780 102.380 -11.780 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.400 102.380 2934.400 102.390 ;
        RECT -14.780 99.380 2934.400 102.380 ;
        RECT -14.780 99.370 -11.780 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.400 99.370 2934.400 99.380 ;
        RECT -14.780 -6.420 -11.780 -6.410 ;
        RECT 94.020 -6.420 97.020 -6.410 ;
        RECT 274.020 -6.420 277.020 -6.410 ;
        RECT 454.020 -6.420 457.020 -6.410 ;
        RECT 634.020 -6.420 637.020 -6.410 ;
        RECT 814.020 -6.420 817.020 -6.410 ;
        RECT 994.020 -6.420 997.020 -6.410 ;
        RECT 1174.020 -6.420 1177.020 -6.410 ;
        RECT 1354.020 -6.420 1357.020 -6.410 ;
        RECT 1534.020 -6.420 1537.020 -6.410 ;
        RECT 1714.020 -6.420 1717.020 -6.410 ;
        RECT 1894.020 -6.420 1897.020 -6.410 ;
        RECT 2074.020 -6.420 2077.020 -6.410 ;
        RECT 2254.020 -6.420 2257.020 -6.410 ;
        RECT 2434.020 -6.420 2437.020 -6.410 ;
        RECT 2614.020 -6.420 2617.020 -6.410 ;
        RECT 2794.020 -6.420 2797.020 -6.410 ;
        RECT 2931.400 -6.420 2934.400 -6.410 ;
        RECT -14.780 -9.420 2934.400 -6.420 ;
        RECT -14.780 -9.430 -11.780 -9.420 ;
        RECT 94.020 -9.430 97.020 -9.420 ;
        RECT 274.020 -9.430 277.020 -9.420 ;
        RECT 454.020 -9.430 457.020 -9.420 ;
        RECT 634.020 -9.430 637.020 -9.420 ;
        RECT 814.020 -9.430 817.020 -9.420 ;
        RECT 994.020 -9.430 997.020 -9.420 ;
        RECT 1174.020 -9.430 1177.020 -9.420 ;
        RECT 1354.020 -9.430 1357.020 -9.420 ;
        RECT 1534.020 -9.430 1537.020 -9.420 ;
        RECT 1714.020 -9.430 1717.020 -9.420 ;
        RECT 1894.020 -9.430 1897.020 -9.420 ;
        RECT 2074.020 -9.430 2077.020 -9.420 ;
        RECT 2254.020 -9.430 2257.020 -9.420 ;
        RECT 2434.020 -9.430 2437.020 -9.420 ;
        RECT 2614.020 -9.430 2617.020 -9.420 ;
        RECT 2794.020 -9.430 2797.020 -9.420 ;
        RECT 2931.400 -9.430 2934.400 -9.420 ;
        RECT -24.380 -16.020 -21.380 -16.010 ;
        RECT 112.020 -16.020 115.020 -16.010 ;
        RECT 292.020 -16.020 295.020 -16.010 ;
        RECT 472.020 -16.020 475.020 -16.010 ;
        RECT 652.020 -16.020 655.020 -16.010 ;
        RECT 832.020 -16.020 835.020 -16.010 ;
        RECT 1012.020 -16.020 1015.020 -16.010 ;
        RECT 1192.020 -16.020 1195.020 -16.010 ;
        RECT 1372.020 -16.020 1375.020 -16.010 ;
        RECT 1552.020 -16.020 1555.020 -16.010 ;
        RECT 1732.020 -16.020 1735.020 -16.010 ;
        RECT 1912.020 -16.020 1915.020 -16.010 ;
        RECT 2092.020 -16.020 2095.020 -16.010 ;
        RECT 2272.020 -16.020 2275.020 -16.010 ;
        RECT 2452.020 -16.020 2455.020 -16.010 ;
        RECT 2632.020 -16.020 2635.020 -16.010 ;
        RECT 2812.020 -16.020 2815.020 -16.010 ;
        RECT 2941.000 -16.020 2944.000 -16.010 ;
        RECT -24.380 -19.020 2944.000 -16.020 ;
        RECT -24.380 -19.030 -21.380 -19.020 ;
        RECT 112.020 -19.030 115.020 -19.020 ;
        RECT 292.020 -19.030 295.020 -19.020 ;
        RECT 472.020 -19.030 475.020 -19.020 ;
        RECT 652.020 -19.030 655.020 -19.020 ;
        RECT 832.020 -19.030 835.020 -19.020 ;
        RECT 1012.020 -19.030 1015.020 -19.020 ;
        RECT 1192.020 -19.030 1195.020 -19.020 ;
        RECT 1372.020 -19.030 1375.020 -19.020 ;
        RECT 1552.020 -19.030 1555.020 -19.020 ;
        RECT 1732.020 -19.030 1735.020 -19.020 ;
        RECT 1912.020 -19.030 1915.020 -19.020 ;
        RECT 2092.020 -19.030 2095.020 -19.020 ;
        RECT 2272.020 -19.030 2275.020 -19.020 ;
        RECT 2452.020 -19.030 2455.020 -19.020 ;
        RECT 2632.020 -19.030 2635.020 -19.020 ;
        RECT 2812.020 -19.030 2815.020 -19.020 ;
        RECT 2941.000 -19.030 2944.000 -19.020 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 665.520 970.795 2245.620 2551.285 ;
      LAYER met1 ;
        RECT 661.910 969.560 2245.620 2551.440 ;
      LAYER met2 ;
        RECT 661.940 2557.905 689.250 2558.185 ;
        RECT 690.090 2557.905 748.130 2558.185 ;
        RECT 748.970 2557.905 807.010 2558.185 ;
        RECT 807.850 2557.905 865.890 2558.185 ;
        RECT 866.730 2557.905 924.770 2558.185 ;
        RECT 925.610 2557.905 983.650 2558.185 ;
        RECT 984.490 2557.905 1042.530 2558.185 ;
        RECT 1043.370 2557.905 1101.870 2558.185 ;
        RECT 1102.710 2557.905 1160.750 2558.185 ;
        RECT 1161.590 2557.905 1219.630 2558.185 ;
        RECT 1220.470 2557.905 1278.510 2558.185 ;
        RECT 1279.350 2557.905 1337.390 2558.185 ;
        RECT 1338.230 2557.905 1396.270 2558.185 ;
        RECT 1397.110 2557.905 1455.150 2558.185 ;
        RECT 1455.990 2557.905 1514.490 2558.185 ;
        RECT 1515.330 2557.905 1573.370 2558.185 ;
        RECT 1574.210 2557.905 1632.250 2558.185 ;
        RECT 1633.090 2557.905 1691.130 2558.185 ;
        RECT 1691.970 2557.905 1750.010 2558.185 ;
        RECT 1750.850 2557.905 1808.890 2558.185 ;
        RECT 1809.730 2557.905 1867.770 2558.185 ;
        RECT 1868.610 2557.905 1927.110 2558.185 ;
        RECT 1927.950 2557.905 1985.990 2558.185 ;
        RECT 1986.830 2557.905 2044.870 2558.185 ;
        RECT 2045.710 2557.905 2103.750 2558.185 ;
        RECT 2104.590 2557.905 2162.630 2558.185 ;
        RECT 2163.470 2557.905 2221.510 2558.185 ;
        RECT 2222.350 2557.905 2245.520 2558.185 ;
        RECT 661.940 964.280 2245.520 2557.905 ;
        RECT 662.490 964.000 665.330 964.280 ;
        RECT 666.170 964.000 669.470 964.280 ;
        RECT 670.310 964.000 673.610 964.280 ;
        RECT 674.450 964.000 677.750 964.280 ;
        RECT 678.590 964.000 681.890 964.280 ;
        RECT 682.730 964.000 686.030 964.280 ;
        RECT 686.870 964.000 690.170 964.280 ;
        RECT 691.010 964.000 694.310 964.280 ;
        RECT 695.150 964.000 698.450 964.280 ;
        RECT 699.290 964.000 702.590 964.280 ;
        RECT 703.430 964.000 706.730 964.280 ;
        RECT 707.570 964.000 710.870 964.280 ;
        RECT 711.710 964.000 715.010 964.280 ;
        RECT 715.850 964.000 719.150 964.280 ;
        RECT 719.990 964.000 723.290 964.280 ;
        RECT 724.130 964.000 727.430 964.280 ;
        RECT 728.270 964.000 731.570 964.280 ;
        RECT 732.410 964.000 735.710 964.280 ;
        RECT 736.550 964.000 739.850 964.280 ;
        RECT 740.690 964.000 743.990 964.280 ;
        RECT 744.830 964.000 748.130 964.280 ;
        RECT 748.970 964.000 752.270 964.280 ;
        RECT 753.110 964.000 756.410 964.280 ;
        RECT 757.250 964.000 760.550 964.280 ;
        RECT 761.390 964.000 764.690 964.280 ;
        RECT 765.530 964.000 768.830 964.280 ;
        RECT 769.670 964.000 772.970 964.280 ;
        RECT 773.810 964.000 776.650 964.280 ;
        RECT 777.490 964.000 780.790 964.280 ;
        RECT 781.630 964.000 784.930 964.280 ;
        RECT 785.770 964.000 789.070 964.280 ;
        RECT 789.910 964.000 793.210 964.280 ;
        RECT 794.050 964.000 797.350 964.280 ;
        RECT 798.190 964.000 801.490 964.280 ;
        RECT 802.330 964.000 805.630 964.280 ;
        RECT 806.470 964.000 809.770 964.280 ;
        RECT 810.610 964.000 813.910 964.280 ;
        RECT 814.750 964.000 818.050 964.280 ;
        RECT 818.890 964.000 822.190 964.280 ;
        RECT 823.030 964.000 826.330 964.280 ;
        RECT 827.170 964.000 830.470 964.280 ;
        RECT 831.310 964.000 834.610 964.280 ;
        RECT 835.450 964.000 838.750 964.280 ;
        RECT 839.590 964.000 842.890 964.280 ;
        RECT 843.730 964.000 847.030 964.280 ;
        RECT 847.870 964.000 851.170 964.280 ;
        RECT 852.010 964.000 855.310 964.280 ;
        RECT 856.150 964.000 859.450 964.280 ;
        RECT 860.290 964.000 863.590 964.280 ;
        RECT 864.430 964.000 867.730 964.280 ;
        RECT 868.570 964.000 871.870 964.280 ;
        RECT 872.710 964.000 876.010 964.280 ;
        RECT 876.850 964.000 880.150 964.280 ;
        RECT 880.990 964.000 884.290 964.280 ;
        RECT 885.130 964.000 888.430 964.280 ;
        RECT 889.270 964.000 892.110 964.280 ;
        RECT 892.950 964.000 896.250 964.280 ;
        RECT 897.090 964.000 900.390 964.280 ;
        RECT 901.230 964.000 904.530 964.280 ;
        RECT 905.370 964.000 908.670 964.280 ;
        RECT 909.510 964.000 912.810 964.280 ;
        RECT 913.650 964.000 916.950 964.280 ;
        RECT 917.790 964.000 921.090 964.280 ;
        RECT 921.930 964.000 925.230 964.280 ;
        RECT 926.070 964.000 929.370 964.280 ;
        RECT 930.210 964.000 933.510 964.280 ;
        RECT 934.350 964.000 937.650 964.280 ;
        RECT 938.490 964.000 941.790 964.280 ;
        RECT 942.630 964.000 945.930 964.280 ;
        RECT 946.770 964.000 950.070 964.280 ;
        RECT 950.910 964.000 954.210 964.280 ;
        RECT 955.050 964.000 958.350 964.280 ;
        RECT 959.190 964.000 962.490 964.280 ;
        RECT 963.330 964.000 966.630 964.280 ;
        RECT 967.470 964.000 970.770 964.280 ;
        RECT 971.610 964.000 974.910 964.280 ;
        RECT 975.750 964.000 979.050 964.280 ;
        RECT 979.890 964.000 983.190 964.280 ;
        RECT 984.030 964.000 987.330 964.280 ;
        RECT 988.170 964.000 991.470 964.280 ;
        RECT 992.310 964.000 995.610 964.280 ;
        RECT 996.450 964.000 999.750 964.280 ;
        RECT 1000.590 964.000 1003.430 964.280 ;
        RECT 1004.270 964.000 1007.570 964.280 ;
        RECT 1008.410 964.000 1011.710 964.280 ;
        RECT 1012.550 964.000 1015.850 964.280 ;
        RECT 1016.690 964.000 1019.990 964.280 ;
        RECT 1020.830 964.000 1024.130 964.280 ;
        RECT 1024.970 964.000 1028.270 964.280 ;
        RECT 1029.110 964.000 1032.410 964.280 ;
        RECT 1033.250 964.000 1036.550 964.280 ;
        RECT 1037.390 964.000 1040.690 964.280 ;
        RECT 1041.530 964.000 1044.830 964.280 ;
        RECT 1045.670 964.000 1048.970 964.280 ;
        RECT 1049.810 964.000 1053.110 964.280 ;
        RECT 1053.950 964.000 1057.250 964.280 ;
        RECT 1058.090 964.000 1061.390 964.280 ;
        RECT 1062.230 964.000 1065.530 964.280 ;
        RECT 1066.370 964.000 1069.670 964.280 ;
        RECT 1070.510 964.000 1073.810 964.280 ;
        RECT 1074.650 964.000 1077.950 964.280 ;
        RECT 1078.790 964.000 1082.090 964.280 ;
        RECT 1082.930 964.000 1086.230 964.280 ;
        RECT 1087.070 964.000 1090.370 964.280 ;
        RECT 1091.210 964.000 1094.510 964.280 ;
        RECT 1095.350 964.000 1098.650 964.280 ;
        RECT 1099.490 964.000 1102.790 964.280 ;
        RECT 1103.630 964.000 1106.930 964.280 ;
        RECT 1107.770 964.000 1111.070 964.280 ;
        RECT 1111.910 964.000 1115.210 964.280 ;
        RECT 1116.050 964.000 1118.890 964.280 ;
        RECT 1119.730 964.000 1123.030 964.280 ;
        RECT 1123.870 964.000 1127.170 964.280 ;
        RECT 1128.010 964.000 1131.310 964.280 ;
        RECT 1132.150 964.000 1135.450 964.280 ;
        RECT 1136.290 964.000 1139.590 964.280 ;
        RECT 1140.430 964.000 1143.730 964.280 ;
        RECT 1144.570 964.000 1147.870 964.280 ;
        RECT 1148.710 964.000 1152.010 964.280 ;
        RECT 1152.850 964.000 1156.150 964.280 ;
        RECT 1156.990 964.000 1160.290 964.280 ;
        RECT 1161.130 964.000 1164.430 964.280 ;
        RECT 1165.270 964.000 1168.570 964.280 ;
        RECT 1169.410 964.000 1172.710 964.280 ;
        RECT 1173.550 964.000 1176.850 964.280 ;
        RECT 1177.690 964.000 1180.990 964.280 ;
        RECT 1181.830 964.000 1185.130 964.280 ;
        RECT 1185.970 964.000 1189.270 964.280 ;
        RECT 1190.110 964.000 1193.410 964.280 ;
        RECT 1194.250 964.000 1197.550 964.280 ;
        RECT 1198.390 964.000 1201.690 964.280 ;
        RECT 1202.530 964.000 1205.830 964.280 ;
        RECT 1206.670 964.000 1209.970 964.280 ;
        RECT 1210.810 964.000 1214.110 964.280 ;
        RECT 1214.950 964.000 1218.250 964.280 ;
        RECT 1219.090 964.000 1222.390 964.280 ;
        RECT 1223.230 964.000 1226.530 964.280 ;
        RECT 1227.370 964.000 1230.210 964.280 ;
        RECT 1231.050 964.000 1234.350 964.280 ;
        RECT 1235.190 964.000 1238.490 964.280 ;
        RECT 1239.330 964.000 1242.630 964.280 ;
        RECT 1243.470 964.000 1246.770 964.280 ;
        RECT 1247.610 964.000 1250.910 964.280 ;
        RECT 1251.750 964.000 1255.050 964.280 ;
        RECT 1255.890 964.000 1259.190 964.280 ;
        RECT 1260.030 964.000 1263.330 964.280 ;
        RECT 1264.170 964.000 1267.470 964.280 ;
        RECT 1268.310 964.000 1271.610 964.280 ;
        RECT 1272.450 964.000 1275.750 964.280 ;
        RECT 1276.590 964.000 1279.890 964.280 ;
        RECT 1280.730 964.000 1284.030 964.280 ;
        RECT 1284.870 964.000 1288.170 964.280 ;
        RECT 1289.010 964.000 1292.310 964.280 ;
        RECT 1293.150 964.000 1296.450 964.280 ;
        RECT 1297.290 964.000 1300.590 964.280 ;
        RECT 1301.430 964.000 1304.730 964.280 ;
        RECT 1305.570 964.000 1308.870 964.280 ;
        RECT 1309.710 964.000 1313.010 964.280 ;
        RECT 1313.850 964.000 1317.150 964.280 ;
        RECT 1317.990 964.000 1321.290 964.280 ;
        RECT 1322.130 964.000 1325.430 964.280 ;
        RECT 1326.270 964.000 1329.570 964.280 ;
        RECT 1330.410 964.000 1333.710 964.280 ;
        RECT 1334.550 964.000 1337.850 964.280 ;
        RECT 1338.690 964.000 1341.990 964.280 ;
        RECT 1342.830 964.000 1345.670 964.280 ;
        RECT 1346.510 964.000 1349.810 964.280 ;
        RECT 1350.650 964.000 1353.950 964.280 ;
        RECT 1354.790 964.000 1358.090 964.280 ;
        RECT 1358.930 964.000 1362.230 964.280 ;
        RECT 1363.070 964.000 1366.370 964.280 ;
        RECT 1367.210 964.000 1370.510 964.280 ;
        RECT 1371.350 964.000 1374.650 964.280 ;
        RECT 1375.490 964.000 1378.790 964.280 ;
        RECT 1379.630 964.000 1382.930 964.280 ;
        RECT 1383.770 964.000 1387.070 964.280 ;
        RECT 1387.910 964.000 1391.210 964.280 ;
        RECT 1392.050 964.000 1395.350 964.280 ;
        RECT 1396.190 964.000 1399.490 964.280 ;
        RECT 1400.330 964.000 1403.630 964.280 ;
        RECT 1404.470 964.000 1407.770 964.280 ;
        RECT 1408.610 964.000 1411.910 964.280 ;
        RECT 1412.750 964.000 1416.050 964.280 ;
        RECT 1416.890 964.000 1420.190 964.280 ;
        RECT 1421.030 964.000 1424.330 964.280 ;
        RECT 1425.170 964.000 1428.470 964.280 ;
        RECT 1429.310 964.000 1432.610 964.280 ;
        RECT 1433.450 964.000 1436.750 964.280 ;
        RECT 1437.590 964.000 1440.890 964.280 ;
        RECT 1441.730 964.000 1445.030 964.280 ;
        RECT 1445.870 964.000 1449.170 964.280 ;
        RECT 1450.010 964.000 1453.310 964.280 ;
        RECT 1454.150 964.000 1457.450 964.280 ;
        RECT 1458.290 964.000 1461.130 964.280 ;
        RECT 1461.970 964.000 1465.270 964.280 ;
        RECT 1466.110 964.000 1469.410 964.280 ;
        RECT 1470.250 964.000 1473.550 964.280 ;
        RECT 1474.390 964.000 1477.690 964.280 ;
        RECT 1478.530 964.000 1481.830 964.280 ;
        RECT 1482.670 964.000 1485.970 964.280 ;
        RECT 1486.810 964.000 1490.110 964.280 ;
        RECT 1490.950 964.000 1494.250 964.280 ;
        RECT 1495.090 964.000 1498.390 964.280 ;
        RECT 1499.230 964.000 1502.530 964.280 ;
        RECT 1503.370 964.000 1506.670 964.280 ;
        RECT 1507.510 964.000 1510.810 964.280 ;
        RECT 1511.650 964.000 1514.950 964.280 ;
        RECT 1515.790 964.000 1519.090 964.280 ;
        RECT 1519.930 964.000 1523.230 964.280 ;
        RECT 1524.070 964.000 1527.370 964.280 ;
        RECT 1528.210 964.000 1531.510 964.280 ;
        RECT 1532.350 964.000 1535.650 964.280 ;
        RECT 1536.490 964.000 1539.790 964.280 ;
        RECT 1540.630 964.000 1543.930 964.280 ;
        RECT 1544.770 964.000 1548.070 964.280 ;
        RECT 1548.910 964.000 1552.210 964.280 ;
        RECT 1553.050 964.000 1556.350 964.280 ;
        RECT 1557.190 964.000 1560.490 964.280 ;
        RECT 1561.330 964.000 1564.630 964.280 ;
        RECT 1565.470 964.000 1568.770 964.280 ;
        RECT 1569.610 964.000 1572.450 964.280 ;
        RECT 1573.290 964.000 1576.590 964.280 ;
        RECT 1577.430 964.000 1580.730 964.280 ;
        RECT 1581.570 964.000 1584.870 964.280 ;
        RECT 1585.710 964.000 1589.010 964.280 ;
        RECT 1589.850 964.000 1593.150 964.280 ;
        RECT 1593.990 964.000 1597.290 964.280 ;
        RECT 1598.130 964.000 1601.430 964.280 ;
        RECT 1602.270 964.000 1605.570 964.280 ;
        RECT 1606.410 964.000 1609.710 964.280 ;
        RECT 1610.550 964.000 1613.850 964.280 ;
        RECT 1614.690 964.000 1617.990 964.280 ;
        RECT 1618.830 964.000 1622.130 964.280 ;
        RECT 1622.970 964.000 1626.270 964.280 ;
        RECT 1627.110 964.000 1630.410 964.280 ;
        RECT 1631.250 964.000 1634.550 964.280 ;
        RECT 1635.390 964.000 1638.690 964.280 ;
        RECT 1639.530 964.000 1642.830 964.280 ;
        RECT 1643.670 964.000 1646.970 964.280 ;
        RECT 1647.810 964.000 1651.110 964.280 ;
        RECT 1651.950 964.000 1655.250 964.280 ;
        RECT 1656.090 964.000 1659.390 964.280 ;
        RECT 1660.230 964.000 1663.530 964.280 ;
        RECT 1664.370 964.000 1667.670 964.280 ;
        RECT 1668.510 964.000 1671.810 964.280 ;
        RECT 1672.650 964.000 1675.950 964.280 ;
        RECT 1676.790 964.000 1680.090 964.280 ;
        RECT 1680.930 964.000 1684.230 964.280 ;
        RECT 1685.070 964.000 1687.910 964.280 ;
        RECT 1688.750 964.000 1692.050 964.280 ;
        RECT 1692.890 964.000 1696.190 964.280 ;
        RECT 1697.030 964.000 1700.330 964.280 ;
        RECT 1701.170 964.000 1704.470 964.280 ;
        RECT 1705.310 964.000 1708.610 964.280 ;
        RECT 1709.450 964.000 1712.750 964.280 ;
        RECT 1713.590 964.000 1716.890 964.280 ;
        RECT 1717.730 964.000 1721.030 964.280 ;
        RECT 1721.870 964.000 1725.170 964.280 ;
        RECT 1726.010 964.000 1729.310 964.280 ;
        RECT 1730.150 964.000 1733.450 964.280 ;
        RECT 1734.290 964.000 1737.590 964.280 ;
        RECT 1738.430 964.000 1741.730 964.280 ;
        RECT 1742.570 964.000 1745.870 964.280 ;
        RECT 1746.710 964.000 1750.010 964.280 ;
        RECT 1750.850 964.000 1754.150 964.280 ;
        RECT 1754.990 964.000 1758.290 964.280 ;
        RECT 1759.130 964.000 1762.430 964.280 ;
        RECT 1763.270 964.000 1766.570 964.280 ;
        RECT 1767.410 964.000 1770.710 964.280 ;
        RECT 1771.550 964.000 1774.850 964.280 ;
        RECT 1775.690 964.000 1778.990 964.280 ;
        RECT 1779.830 964.000 1783.130 964.280 ;
        RECT 1783.970 964.000 1787.270 964.280 ;
        RECT 1788.110 964.000 1791.410 964.280 ;
        RECT 1792.250 964.000 1795.550 964.280 ;
        RECT 1796.390 964.000 1799.230 964.280 ;
        RECT 1800.070 964.000 1803.370 964.280 ;
        RECT 1804.210 964.000 1807.510 964.280 ;
        RECT 1808.350 964.000 1811.650 964.280 ;
        RECT 1812.490 964.000 1815.790 964.280 ;
        RECT 1816.630 964.000 1819.930 964.280 ;
        RECT 1820.770 964.000 1824.070 964.280 ;
        RECT 1824.910 964.000 1828.210 964.280 ;
        RECT 1829.050 964.000 1832.350 964.280 ;
        RECT 1833.190 964.000 1836.490 964.280 ;
        RECT 1837.330 964.000 1840.630 964.280 ;
        RECT 1841.470 964.000 1844.770 964.280 ;
        RECT 1845.610 964.000 1848.910 964.280 ;
        RECT 1849.750 964.000 1853.050 964.280 ;
        RECT 1853.890 964.000 1857.190 964.280 ;
        RECT 1858.030 964.000 1861.330 964.280 ;
        RECT 1862.170 964.000 1865.470 964.280 ;
        RECT 1866.310 964.000 1869.610 964.280 ;
        RECT 1870.450 964.000 1873.750 964.280 ;
        RECT 1874.590 964.000 1877.890 964.280 ;
        RECT 1878.730 964.000 1882.030 964.280 ;
        RECT 1882.870 964.000 1886.170 964.280 ;
        RECT 1887.010 964.000 1890.310 964.280 ;
        RECT 1891.150 964.000 1894.450 964.280 ;
        RECT 1895.290 964.000 1898.590 964.280 ;
        RECT 1899.430 964.000 1902.730 964.280 ;
        RECT 1903.570 964.000 1906.870 964.280 ;
        RECT 1907.710 964.000 1911.010 964.280 ;
        RECT 1911.850 964.000 1914.690 964.280 ;
        RECT 1915.530 964.000 1918.830 964.280 ;
        RECT 1919.670 964.000 1922.970 964.280 ;
        RECT 1923.810 964.000 1927.110 964.280 ;
        RECT 1927.950 964.000 1931.250 964.280 ;
        RECT 1932.090 964.000 1935.390 964.280 ;
        RECT 1936.230 964.000 1939.530 964.280 ;
        RECT 1940.370 964.000 1943.670 964.280 ;
        RECT 1944.510 964.000 1947.810 964.280 ;
        RECT 1948.650 964.000 1951.950 964.280 ;
        RECT 1952.790 964.000 1956.090 964.280 ;
        RECT 1956.930 964.000 1960.230 964.280 ;
        RECT 1961.070 964.000 1964.370 964.280 ;
        RECT 1965.210 964.000 1968.510 964.280 ;
        RECT 1969.350 964.000 1972.650 964.280 ;
        RECT 1973.490 964.000 1976.790 964.280 ;
        RECT 1977.630 964.000 1980.930 964.280 ;
        RECT 1981.770 964.000 1985.070 964.280 ;
        RECT 1985.910 964.000 1989.210 964.280 ;
        RECT 1990.050 964.000 1993.350 964.280 ;
        RECT 1994.190 964.000 1997.490 964.280 ;
        RECT 1998.330 964.000 2001.630 964.280 ;
        RECT 2002.470 964.000 2005.770 964.280 ;
        RECT 2006.610 964.000 2009.910 964.280 ;
        RECT 2010.750 964.000 2014.050 964.280 ;
        RECT 2014.890 964.000 2018.190 964.280 ;
        RECT 2019.030 964.000 2022.330 964.280 ;
        RECT 2023.170 964.000 2026.010 964.280 ;
        RECT 2026.850 964.000 2030.150 964.280 ;
        RECT 2030.990 964.000 2034.290 964.280 ;
        RECT 2035.130 964.000 2038.430 964.280 ;
        RECT 2039.270 964.000 2042.570 964.280 ;
        RECT 2043.410 964.000 2046.710 964.280 ;
        RECT 2047.550 964.000 2050.850 964.280 ;
        RECT 2051.690 964.000 2054.990 964.280 ;
        RECT 2055.830 964.000 2059.130 964.280 ;
        RECT 2059.970 964.000 2063.270 964.280 ;
        RECT 2064.110 964.000 2067.410 964.280 ;
        RECT 2068.250 964.000 2071.550 964.280 ;
        RECT 2072.390 964.000 2075.690 964.280 ;
        RECT 2076.530 964.000 2079.830 964.280 ;
        RECT 2080.670 964.000 2083.970 964.280 ;
        RECT 2084.810 964.000 2088.110 964.280 ;
        RECT 2088.950 964.000 2092.250 964.280 ;
        RECT 2093.090 964.000 2096.390 964.280 ;
        RECT 2097.230 964.000 2100.530 964.280 ;
        RECT 2101.370 964.000 2104.670 964.280 ;
        RECT 2105.510 964.000 2108.810 964.280 ;
        RECT 2109.650 964.000 2112.950 964.280 ;
        RECT 2113.790 964.000 2117.090 964.280 ;
        RECT 2117.930 964.000 2121.230 964.280 ;
        RECT 2122.070 964.000 2125.370 964.280 ;
        RECT 2126.210 964.000 2129.510 964.280 ;
        RECT 2130.350 964.000 2133.650 964.280 ;
        RECT 2134.490 964.000 2137.790 964.280 ;
        RECT 2138.630 964.000 2141.470 964.280 ;
        RECT 2142.310 964.000 2145.610 964.280 ;
        RECT 2146.450 964.000 2149.750 964.280 ;
        RECT 2150.590 964.000 2153.890 964.280 ;
        RECT 2154.730 964.000 2158.030 964.280 ;
        RECT 2158.870 964.000 2162.170 964.280 ;
        RECT 2163.010 964.000 2166.310 964.280 ;
        RECT 2167.150 964.000 2170.450 964.280 ;
        RECT 2171.290 964.000 2174.590 964.280 ;
        RECT 2175.430 964.000 2178.730 964.280 ;
        RECT 2179.570 964.000 2182.870 964.280 ;
        RECT 2183.710 964.000 2187.010 964.280 ;
        RECT 2187.850 964.000 2191.150 964.280 ;
        RECT 2191.990 964.000 2195.290 964.280 ;
        RECT 2196.130 964.000 2199.430 964.280 ;
        RECT 2200.270 964.000 2203.570 964.280 ;
        RECT 2204.410 964.000 2207.710 964.280 ;
        RECT 2208.550 964.000 2211.850 964.280 ;
        RECT 2212.690 964.000 2215.990 964.280 ;
        RECT 2216.830 964.000 2220.130 964.280 ;
        RECT 2220.970 964.000 2224.270 964.280 ;
        RECT 2225.110 964.000 2228.410 964.280 ;
        RECT 2229.250 964.000 2232.550 964.280 ;
        RECT 2233.390 964.000 2236.690 964.280 ;
        RECT 2237.530 964.000 2240.830 964.280 ;
        RECT 2241.670 964.000 2244.970 964.280 ;
      LAYER met3 ;
        RECT 663.990 2544.760 2247.610 2551.365 ;
        RECT 663.990 2543.400 2247.065 2544.760 ;
        RECT 664.400 2543.360 2247.065 2543.400 ;
        RECT 664.400 2542.000 2247.610 2543.360 ;
        RECT 663.990 2509.400 2247.610 2542.000 ;
        RECT 663.990 2508.000 2247.065 2509.400 ;
        RECT 663.990 2505.320 2247.610 2508.000 ;
        RECT 664.400 2503.920 2247.610 2505.320 ;
        RECT 663.990 2473.360 2247.610 2503.920 ;
        RECT 663.990 2471.960 2247.065 2473.360 ;
        RECT 663.990 2467.240 2247.610 2471.960 ;
        RECT 664.400 2465.840 2247.610 2467.240 ;
        RECT 663.990 2438.000 2247.610 2465.840 ;
        RECT 663.990 2436.600 2247.065 2438.000 ;
        RECT 663.990 2429.160 2247.610 2436.600 ;
        RECT 664.400 2427.760 2247.610 2429.160 ;
        RECT 663.990 2402.640 2247.610 2427.760 ;
        RECT 663.990 2401.240 2247.065 2402.640 ;
        RECT 663.990 2391.080 2247.610 2401.240 ;
        RECT 664.400 2389.680 2247.610 2391.080 ;
        RECT 663.990 2366.600 2247.610 2389.680 ;
        RECT 663.990 2365.200 2247.065 2366.600 ;
        RECT 663.990 2353.000 2247.610 2365.200 ;
        RECT 664.400 2351.600 2247.610 2353.000 ;
        RECT 663.990 2331.240 2247.610 2351.600 ;
        RECT 663.990 2329.840 2247.065 2331.240 ;
        RECT 663.990 2314.920 2247.610 2329.840 ;
        RECT 664.400 2313.520 2247.610 2314.920 ;
        RECT 663.990 2295.880 2247.610 2313.520 ;
        RECT 663.990 2294.480 2247.065 2295.880 ;
        RECT 663.990 2276.840 2247.610 2294.480 ;
        RECT 664.400 2275.440 2247.610 2276.840 ;
        RECT 663.990 2259.840 2247.610 2275.440 ;
        RECT 663.990 2258.440 2247.065 2259.840 ;
        RECT 663.990 2238.760 2247.610 2258.440 ;
        RECT 664.400 2237.360 2247.610 2238.760 ;
        RECT 663.990 2224.480 2247.610 2237.360 ;
        RECT 663.990 2223.080 2247.065 2224.480 ;
        RECT 663.990 2200.680 2247.610 2223.080 ;
        RECT 664.400 2199.280 2247.610 2200.680 ;
        RECT 663.990 2189.120 2247.610 2199.280 ;
        RECT 663.990 2187.720 2247.065 2189.120 ;
        RECT 663.990 2161.920 2247.610 2187.720 ;
        RECT 664.400 2160.520 2247.610 2161.920 ;
        RECT 663.990 2153.080 2247.610 2160.520 ;
        RECT 663.990 2151.680 2247.065 2153.080 ;
        RECT 663.990 2123.840 2247.610 2151.680 ;
        RECT 664.400 2122.440 2247.610 2123.840 ;
        RECT 663.990 2117.720 2247.610 2122.440 ;
        RECT 663.990 2116.320 2247.065 2117.720 ;
        RECT 663.990 2085.760 2247.610 2116.320 ;
        RECT 664.400 2084.360 2247.610 2085.760 ;
        RECT 663.990 2082.360 2247.610 2084.360 ;
        RECT 663.990 2080.960 2247.065 2082.360 ;
        RECT 663.990 2047.680 2247.610 2080.960 ;
        RECT 664.400 2046.320 2247.610 2047.680 ;
        RECT 664.400 2046.280 2247.065 2046.320 ;
        RECT 663.990 2044.920 2247.065 2046.280 ;
        RECT 663.990 2010.960 2247.610 2044.920 ;
        RECT 663.990 2009.600 2247.065 2010.960 ;
        RECT 664.400 2009.560 2247.065 2009.600 ;
        RECT 664.400 2008.200 2247.610 2009.560 ;
        RECT 663.990 1974.920 2247.610 2008.200 ;
        RECT 663.990 1973.520 2247.065 1974.920 ;
        RECT 663.990 1971.520 2247.610 1973.520 ;
        RECT 664.400 1970.120 2247.610 1971.520 ;
        RECT 663.990 1939.560 2247.610 1970.120 ;
        RECT 663.990 1938.160 2247.065 1939.560 ;
        RECT 663.990 1933.440 2247.610 1938.160 ;
        RECT 664.400 1932.040 2247.610 1933.440 ;
        RECT 663.990 1904.200 2247.610 1932.040 ;
        RECT 663.990 1902.800 2247.065 1904.200 ;
        RECT 663.990 1895.360 2247.610 1902.800 ;
        RECT 664.400 1893.960 2247.610 1895.360 ;
        RECT 663.990 1868.160 2247.610 1893.960 ;
        RECT 663.990 1866.760 2247.065 1868.160 ;
        RECT 663.990 1857.280 2247.610 1866.760 ;
        RECT 664.400 1855.880 2247.610 1857.280 ;
        RECT 663.990 1832.800 2247.610 1855.880 ;
        RECT 663.990 1831.400 2247.065 1832.800 ;
        RECT 663.990 1819.200 2247.610 1831.400 ;
        RECT 664.400 1817.800 2247.610 1819.200 ;
        RECT 663.990 1797.440 2247.610 1817.800 ;
        RECT 663.990 1796.040 2247.065 1797.440 ;
        RECT 663.990 1781.120 2247.610 1796.040 ;
        RECT 664.400 1779.720 2247.610 1781.120 ;
        RECT 663.990 1761.400 2247.610 1779.720 ;
        RECT 663.990 1760.000 2247.065 1761.400 ;
        RECT 663.990 1742.360 2247.610 1760.000 ;
        RECT 664.400 1740.960 2247.610 1742.360 ;
        RECT 663.990 1726.040 2247.610 1740.960 ;
        RECT 663.990 1724.640 2247.065 1726.040 ;
        RECT 663.990 1704.280 2247.610 1724.640 ;
        RECT 664.400 1702.880 2247.610 1704.280 ;
        RECT 663.990 1690.680 2247.610 1702.880 ;
        RECT 663.990 1689.280 2247.065 1690.680 ;
        RECT 663.990 1666.200 2247.610 1689.280 ;
        RECT 664.400 1664.800 2247.610 1666.200 ;
        RECT 663.990 1654.640 2247.610 1664.800 ;
        RECT 663.990 1653.240 2247.065 1654.640 ;
        RECT 663.990 1628.120 2247.610 1653.240 ;
        RECT 664.400 1626.720 2247.610 1628.120 ;
        RECT 663.990 1619.280 2247.610 1626.720 ;
        RECT 663.990 1617.880 2247.065 1619.280 ;
        RECT 663.990 1590.040 2247.610 1617.880 ;
        RECT 664.400 1588.640 2247.610 1590.040 ;
        RECT 663.990 1583.920 2247.610 1588.640 ;
        RECT 663.990 1582.520 2247.065 1583.920 ;
        RECT 663.990 1551.960 2247.610 1582.520 ;
        RECT 664.400 1550.560 2247.610 1551.960 ;
        RECT 663.990 1547.880 2247.610 1550.560 ;
        RECT 663.990 1546.480 2247.065 1547.880 ;
        RECT 663.990 1513.880 2247.610 1546.480 ;
        RECT 664.400 1512.520 2247.610 1513.880 ;
        RECT 664.400 1512.480 2247.065 1512.520 ;
        RECT 663.990 1511.120 2247.065 1512.480 ;
        RECT 663.990 1476.480 2247.610 1511.120 ;
        RECT 663.990 1475.800 2247.065 1476.480 ;
        RECT 664.400 1475.080 2247.065 1475.800 ;
        RECT 664.400 1474.400 2247.610 1475.080 ;
        RECT 663.990 1441.120 2247.610 1474.400 ;
        RECT 663.990 1439.720 2247.065 1441.120 ;
        RECT 663.990 1437.720 2247.610 1439.720 ;
        RECT 664.400 1436.320 2247.610 1437.720 ;
        RECT 663.990 1405.760 2247.610 1436.320 ;
        RECT 663.990 1404.360 2247.065 1405.760 ;
        RECT 663.990 1399.640 2247.610 1404.360 ;
        RECT 664.400 1398.240 2247.610 1399.640 ;
        RECT 663.990 1369.720 2247.610 1398.240 ;
        RECT 663.990 1368.320 2247.065 1369.720 ;
        RECT 663.990 1360.880 2247.610 1368.320 ;
        RECT 664.400 1359.480 2247.610 1360.880 ;
        RECT 663.990 1334.360 2247.610 1359.480 ;
        RECT 663.990 1332.960 2247.065 1334.360 ;
        RECT 663.990 1322.800 2247.610 1332.960 ;
        RECT 664.400 1321.400 2247.610 1322.800 ;
        RECT 663.990 1299.000 2247.610 1321.400 ;
        RECT 663.990 1297.600 2247.065 1299.000 ;
        RECT 663.990 1284.720 2247.610 1297.600 ;
        RECT 664.400 1283.320 2247.610 1284.720 ;
        RECT 663.990 1262.960 2247.610 1283.320 ;
        RECT 663.990 1261.560 2247.065 1262.960 ;
        RECT 663.990 1246.640 2247.610 1261.560 ;
        RECT 664.400 1245.240 2247.610 1246.640 ;
        RECT 663.990 1227.600 2247.610 1245.240 ;
        RECT 663.990 1226.200 2247.065 1227.600 ;
        RECT 663.990 1208.560 2247.610 1226.200 ;
        RECT 664.400 1207.160 2247.610 1208.560 ;
        RECT 663.990 1192.240 2247.610 1207.160 ;
        RECT 663.990 1190.840 2247.065 1192.240 ;
        RECT 663.990 1170.480 2247.610 1190.840 ;
        RECT 664.400 1169.080 2247.610 1170.480 ;
        RECT 663.990 1156.200 2247.610 1169.080 ;
        RECT 663.990 1154.800 2247.065 1156.200 ;
        RECT 663.990 1132.400 2247.610 1154.800 ;
        RECT 664.400 1131.000 2247.610 1132.400 ;
        RECT 663.990 1120.840 2247.610 1131.000 ;
        RECT 663.990 1119.440 2247.065 1120.840 ;
        RECT 663.990 1094.320 2247.610 1119.440 ;
        RECT 664.400 1092.920 2247.610 1094.320 ;
        RECT 663.990 1085.480 2247.610 1092.920 ;
        RECT 663.990 1084.080 2247.065 1085.480 ;
        RECT 663.990 1056.240 2247.610 1084.080 ;
        RECT 664.400 1054.840 2247.610 1056.240 ;
        RECT 663.990 1049.440 2247.610 1054.840 ;
        RECT 663.990 1048.040 2247.065 1049.440 ;
        RECT 663.990 1018.160 2247.610 1048.040 ;
        RECT 664.400 1016.760 2247.610 1018.160 ;
        RECT 663.990 1014.080 2247.610 1016.760 ;
        RECT 663.990 1012.680 2247.065 1014.080 ;
        RECT 663.990 980.080 2247.610 1012.680 ;
        RECT 664.400 978.720 2247.610 980.080 ;
        RECT 664.400 978.680 2247.065 978.720 ;
        RECT 663.990 977.320 2247.065 978.680 ;
        RECT 663.990 964.255 2247.610 977.320 ;
      LAYER met4 ;
        RECT 678.695 970.640 680.640 2551.440 ;
        RECT 683.040 970.640 757.440 2551.440 ;
        RECT 759.840 970.640 2218.640 2551.440 ;
  END
END user_project_wrapper
END LIBRARY

