magic
tech sky130A
magscale 1 2
timestamp 1611548290
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 412649 683247 412683 692733
rect 218989 666587 219023 676141
rect 413017 666587 413051 683077
rect 429577 666587 429611 683077
rect 494069 666587 494103 676141
rect 542737 666587 542771 683077
rect 559297 666587 559331 683077
rect 72985 647275 73019 656829
rect 219265 647275 219299 656829
rect 73077 616879 73111 626501
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 412833 601715 412867 608549
rect 429393 601715 429427 608549
rect 542553 601715 542587 608549
rect 559113 601715 559147 608549
rect 72893 589339 72927 598893
rect 219173 589339 219207 598893
rect 413017 589339 413051 598893
rect 429577 589339 429611 598893
rect 542737 589339 542771 598893
rect 559297 589339 559331 598893
rect 8033 579751 8067 589237
rect 137753 579751 137787 589237
rect 154313 579751 154347 589237
rect 284033 579751 284067 589237
rect 347789 579683 347823 589237
rect 364349 579683 364383 589237
rect 477509 579683 477543 589237
rect 72617 569959 72651 579581
rect 137569 569959 137603 579581
rect 218897 569959 218931 579581
rect 347881 563091 347915 569857
rect 364441 563091 364475 569857
rect 477601 563091 477635 569857
rect 494161 563091 494195 569857
rect 72709 550647 72743 560201
rect 137661 550647 137695 560201
rect 218989 550647 219023 560201
rect 412741 550647 412775 560201
rect 429301 550647 429335 560201
rect 542461 550647 542495 560201
rect 559021 550647 559055 560201
rect 8033 543779 8067 550545
rect 154313 543779 154347 550545
rect 284033 543779 284067 550545
rect 72801 521679 72835 524433
rect 137753 521679 137787 524433
rect 219081 521679 219115 524433
rect 135361 77299 135395 86921
rect 135361 70295 135395 77129
rect 135545 48331 135579 57885
rect 135545 29019 135579 38573
rect 135637 12291 135671 19261
rect 212549 3995 212583 4097
rect 213101 3111 213135 3757
rect 217333 3723 217367 4097
rect 214515 3621 214665 3655
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 412649 692733 412683 692767
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 412649 683213 412683 683247
rect 284033 676209 284067 676243
rect 413017 683077 413051 683111
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 413017 666553 413051 666587
rect 429577 683077 429611 683111
rect 542737 683077 542771 683111
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 542737 666553 542771 666587
rect 559297 683077 559331 683111
rect 559297 666553 559331 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 73077 626501 73111 626535
rect 73077 616845 73111 616879
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 412833 608549 412867 608583
rect 412833 601681 412867 601715
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 542553 608549 542587 608583
rect 542553 601681 542587 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 219265 601545 219299 601579
rect 72893 598893 72927 598927
rect 72893 589305 72927 589339
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 413017 598893 413051 598927
rect 413017 589305 413051 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 542737 598893 542771 598927
rect 542737 589305 542771 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 8033 589237 8067 589271
rect 8033 579717 8067 579751
rect 137753 589237 137787 589271
rect 137753 579717 137787 579751
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 284033 589237 284067 589271
rect 284033 579717 284067 579751
rect 347789 589237 347823 589271
rect 347789 579649 347823 579683
rect 364349 589237 364383 589271
rect 364349 579649 364383 579683
rect 477509 589237 477543 589271
rect 477509 579649 477543 579683
rect 72617 579581 72651 579615
rect 72617 569925 72651 569959
rect 137569 579581 137603 579615
rect 137569 569925 137603 569959
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 347881 569857 347915 569891
rect 347881 563057 347915 563091
rect 364441 569857 364475 569891
rect 364441 563057 364475 563091
rect 477601 569857 477635 569891
rect 477601 563057 477635 563091
rect 494161 569857 494195 569891
rect 494161 563057 494195 563091
rect 72709 560201 72743 560235
rect 72709 550613 72743 550647
rect 137661 560201 137695 560235
rect 137661 550613 137695 550647
rect 218989 560201 219023 560235
rect 218989 550613 219023 550647
rect 412741 560201 412775 560235
rect 412741 550613 412775 550647
rect 429301 560201 429335 560235
rect 429301 550613 429335 550647
rect 542461 560201 542495 560235
rect 542461 550613 542495 550647
rect 559021 560201 559055 560235
rect 559021 550613 559055 550647
rect 8033 550545 8067 550579
rect 8033 543745 8067 543779
rect 154313 550545 154347 550579
rect 154313 543745 154347 543779
rect 284033 550545 284067 550579
rect 284033 543745 284067 543779
rect 72801 524433 72835 524467
rect 72801 521645 72835 521679
rect 137753 524433 137787 524467
rect 137753 521645 137787 521679
rect 219081 524433 219115 524467
rect 219081 521645 219115 521679
rect 135361 86921 135395 86955
rect 135361 77265 135395 77299
rect 135361 77129 135395 77163
rect 135361 70261 135395 70295
rect 135545 57885 135579 57919
rect 135545 48297 135579 48331
rect 135545 38573 135579 38607
rect 135545 28985 135579 29019
rect 135637 19261 135671 19295
rect 135637 12257 135671 12291
rect 212549 4097 212583 4131
rect 212549 3961 212583 3995
rect 217333 4097 217367 4131
rect 213101 3757 213135 3791
rect 217333 3689 217367 3723
rect 214481 3621 214515 3655
rect 214665 3621 214699 3655
rect 213101 3077 213135 3111
<< metal1 >>
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 413002 698232 413008 698284
rect 413060 698272 413066 698284
rect 413738 698272 413744 698284
rect 413060 698244 413744 698272
rect 413060 698232 413066 698244
rect 413738 698232 413744 698244
rect 413796 698232 413802 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 331214 697552 331220 697604
rect 331272 697592 331278 697604
rect 332502 697592 332508 697604
rect 331272 697564 332508 697592
rect 331272 697552 331278 697564
rect 332502 697552 332508 697564
rect 332560 697552 332566 697604
rect 472618 696940 472624 696992
rect 472676 696980 472682 696992
rect 580166 696980 580172 696992
rect 472676 696952 580172 696980
rect 472676 696940 472682 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 412818 694084 412824 694136
rect 412876 694124 412882 694136
rect 413002 694124 413008 694136
rect 412876 694096 413008 694124
rect 412876 694084 412882 694096
rect 413002 694084 413008 694096
rect 413060 694084 413066 694136
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 347774 692792 347780 692844
rect 347832 692832 347838 692844
rect 348878 692832 348884 692844
rect 347832 692804 348884 692832
rect 347832 692792 347838 692804
rect 348878 692792 348884 692804
rect 348936 692792 348942 692844
rect 364334 692792 364340 692844
rect 364392 692832 364398 692844
rect 365070 692832 365076 692844
rect 364392 692804 365076 692832
rect 364392 692792 364398 692804
rect 365070 692792 365076 692804
rect 365128 692792 365134 692844
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 412637 692767 412695 692773
rect 412637 692733 412649 692767
rect 412683 692764 412695 692767
rect 412818 692764 412824 692776
rect 412683 692736 412824 692764
rect 412683 692733 412695 692736
rect 412637 692727 412695 692733
rect 412818 692724 412824 692736
rect 412876 692724 412882 692776
rect 542538 692724 542544 692776
rect 542596 692764 542602 692776
rect 542722 692764 542728 692776
rect 542596 692736 542728 692764
rect 542596 692724 542602 692736
rect 542722 692724 542728 692736
rect 542780 692724 542786 692776
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 494238 685856 494244 685908
rect 494296 685896 494302 685908
rect 494882 685896 494888 685908
rect 494296 685868 494888 685896
rect 494296 685856 494302 685868
rect 494882 685856 494888 685868
rect 494940 685856 494946 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 429194 684428 429200 684480
rect 429252 684468 429258 684480
rect 429838 684468 429844 684480
rect 429252 684440 429844 684468
rect 429252 684428 429258 684440
rect 429838 684428 429844 684440
rect 429896 684428 429902 684480
rect 558914 684428 558920 684480
rect 558972 684468 558978 684480
rect 559650 684468 559656 684480
rect 558972 684440 559656 684468
rect 558972 684428 558978 684440
rect 559650 684428 559656 684440
rect 559708 684428 559714 684480
rect 412634 683204 412640 683256
rect 412692 683244 412698 683256
rect 412692 683216 412737 683244
rect 412692 683204 412698 683216
rect 412634 683068 412640 683120
rect 412692 683108 412698 683120
rect 413005 683111 413063 683117
rect 413005 683108 413017 683111
rect 412692 683080 413017 683108
rect 412692 683068 412698 683080
rect 413005 683077 413017 683080
rect 413051 683077 413063 683111
rect 413005 683071 413063 683077
rect 429194 683068 429200 683120
rect 429252 683108 429258 683120
rect 429565 683111 429623 683117
rect 429565 683108 429577 683111
rect 429252 683080 429577 683108
rect 429252 683068 429258 683080
rect 429565 683077 429577 683080
rect 429611 683077 429623 683111
rect 429565 683071 429623 683077
rect 542354 683068 542360 683120
rect 542412 683108 542418 683120
rect 542725 683111 542783 683117
rect 542725 683108 542737 683111
rect 542412 683080 542737 683108
rect 542412 683068 542418 683080
rect 542725 683077 542737 683080
rect 542771 683077 542783 683111
rect 542725 683071 542783 683077
rect 558914 683068 558920 683120
rect 558972 683108 558978 683120
rect 559285 683111 559343 683117
rect 559285 683108 559297 683111
rect 558972 683080 559297 683108
rect 558972 683068 558978 683080
rect 559285 683077 559297 683080
rect 559331 683077 559343 683111
rect 559285 683071 559343 683077
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 8938 681748 8944 681760
rect 3568 681720 8944 681748
rect 3568 681708 3574 681720
rect 8938 681708 8944 681720
rect 8996 681708 9002 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 347774 673480 347780 673532
rect 347832 673520 347838 673532
rect 347958 673520 347964 673532
rect 347832 673492 347964 673520
rect 347832 673480 347838 673492
rect 347958 673480 347964 673492
rect 348016 673480 348022 673532
rect 364334 673480 364340 673532
rect 364392 673520 364398 673532
rect 364518 673520 364524 673532
rect 364392 673492 364524 673520
rect 364392 673480 364398 673492
rect 364518 673480 364524 673492
rect 364576 673480 364582 673532
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 490558 673480 490564 673532
rect 490616 673520 490622 673532
rect 580166 673520 580172 673532
rect 490616 673492 580172 673520
rect 490616 673480 490622 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 17218 667944 17224 667956
rect 3476 667916 17224 667944
rect 3476 667904 3482 667916
rect 17218 667904 17224 667916
rect 17276 667904 17282 667956
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 413005 666587 413063 666593
rect 413005 666553 413017 666587
rect 413051 666584 413063 666587
rect 413094 666584 413100 666596
rect 413051 666556 413100 666584
rect 413051 666553 413063 666556
rect 413005 666547 413063 666553
rect 413094 666544 413100 666556
rect 413152 666544 413158 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 284018 654100 284024 654152
rect 284076 654140 284082 654152
rect 284202 654140 284208 654152
rect 284076 654112 284208 654140
rect 284076 654100 284082 654112
rect 284202 654100 284208 654112
rect 284260 654100 284266 654152
rect 347774 654100 347780 654152
rect 347832 654140 347838 654152
rect 347958 654140 347964 654152
rect 347832 654112 347964 654140
rect 347832 654100 347838 654112
rect 347958 654100 347964 654112
rect 348016 654100 348022 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 14458 652780 14464 652792
rect 3108 652752 14464 652780
rect 3108 652740 3114 652752
rect 14458 652740 14464 652752
rect 14516 652740 14522 652792
rect 471238 650020 471244 650072
rect 471296 650060 471302 650072
rect 580166 650060 580172 650072
rect 471296 650032 580172 650060
rect 471296 650020 471302 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 412818 647232 412824 647284
rect 412876 647272 412882 647284
rect 412910 647272 412916 647284
rect 412876 647244 412916 647272
rect 412876 647232 412882 647244
rect 412910 647232 412916 647244
rect 412968 647232 412974 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 412818 640364 412824 640416
rect 412876 640404 412882 640416
rect 412910 640404 412916 640416
rect 412876 640376 412916 640404
rect 412876 640364 412882 640376
rect 412910 640364 412916 640376
rect 412968 640364 412974 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 72786 637508 72792 637560
rect 72844 637548 72850 637560
rect 72878 637548 72884 637560
rect 72844 637520 72884 637548
rect 72844 637508 72850 637520
rect 72878 637508 72884 637520
rect 72936 637508 72942 637560
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 137738 634788 137744 634840
rect 137796 634828 137802 634840
rect 137922 634828 137928 634840
rect 137796 634800 137928 634828
rect 137796 634788 137802 634800
rect 137922 634788 137928 634800
rect 137980 634788 137986 634840
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 284018 634788 284024 634840
rect 284076 634828 284082 634840
rect 284202 634828 284208 634840
rect 284076 634800 284208 634828
rect 284076 634788 284082 634800
rect 284202 634788 284208 634800
rect 284260 634788 284266 634840
rect 347774 634788 347780 634840
rect 347832 634828 347838 634840
rect 347958 634828 347964 634840
rect 347832 634800 347964 634828
rect 347832 634788 347838 634800
rect 347958 634788 347964 634800
rect 348016 634788 348022 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 412726 630640 412732 630692
rect 412784 630680 412790 630692
rect 412910 630680 412916 630692
rect 412784 630652 412916 630680
rect 412784 630640 412790 630652
rect 412910 630640 412916 630652
rect 412968 630640 412974 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 479518 626560 479524 626612
rect 479576 626600 479582 626612
rect 580166 626600 580172 626612
rect 479576 626572 580172 626600
rect 479576 626560 479582 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 73062 626532 73068 626544
rect 73023 626504 73068 626532
rect 73062 626492 73068 626504
rect 73120 626492 73126 626544
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 10318 623812 10324 623824
rect 3476 623784 10324 623812
rect 3476 623772 3482 623784
rect 10318 623772 10324 623784
rect 10376 623772 10382 623824
rect 73062 616876 73068 616888
rect 73023 616848 73068 616876
rect 73062 616836 73068 616848
rect 73120 616836 73126 616888
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 137738 615476 137744 615528
rect 137796 615516 137802 615528
rect 137922 615516 137928 615528
rect 137796 615488 137928 615516
rect 137796 615476 137802 615488
rect 137922 615476 137928 615488
rect 137980 615476 137986 615528
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 284018 615476 284024 615528
rect 284076 615516 284082 615528
rect 284202 615516 284208 615528
rect 284076 615488 284208 615516
rect 284076 615476 284082 615488
rect 284202 615476 284208 615488
rect 284260 615476 284266 615528
rect 347774 615476 347780 615528
rect 347832 615516 347838 615528
rect 347958 615516 347964 615528
rect 347832 615488 347964 615516
rect 347832 615476 347838 615488
rect 347958 615476 347964 615488
rect 348016 615476 348022 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 477494 615476 477500 615528
rect 477552 615516 477558 615528
rect 477678 615516 477684 615528
rect 477552 615488 477684 615516
rect 477552 615476 477558 615488
rect 477678 615476 477684 615488
rect 477736 615476 477742 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 73062 611436 73068 611448
rect 72896 611408 73068 611436
rect 72896 611312 72924 611408
rect 73062 611396 73068 611408
rect 73120 611396 73126 611448
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 412726 611328 412732 611380
rect 412784 611368 412790 611380
rect 412910 611368 412916 611380
rect 412784 611340 412916 611368
rect 412784 611328 412790 611340
rect 412910 611328 412916 611340
rect 412968 611328 412974 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 72878 611260 72884 611312
rect 72936 611260 72942 611312
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 19978 610008 19984 610020
rect 3476 609980 19984 610008
rect 3476 609968 3482 609980
rect 19978 609968 19984 609980
rect 20036 609968 20042 610020
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 412818 608580 412824 608592
rect 412779 608552 412824 608580
rect 219253 608543 219311 608549
rect 412818 608540 412824 608552
rect 412876 608540 412882 608592
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 542538 608580 542544 608592
rect 542499 608552 542544 608580
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 467098 603100 467104 603152
rect 467156 603140 467162 603152
rect 580166 603140 580172 603152
rect 467156 603112 580172 603140
rect 467156 603100 467162 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 412821 601715 412879 601721
rect 412821 601681 412833 601715
rect 412867 601712 412879 601715
rect 413002 601712 413008 601724
rect 412867 601684 413008 601712
rect 412867 601681 412879 601684
rect 412821 601675 412879 601681
rect 413002 601672 413008 601684
rect 413060 601672 413066 601724
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 542541 601715 542599 601721
rect 542541 601681 542553 601715
rect 542587 601712 542599 601715
rect 542722 601712 542728 601724
rect 542587 601684 542728 601712
rect 542587 601681 542599 601684
rect 542541 601675 542599 601681
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 72970 601536 72976 601588
rect 73028 601576 73034 601588
rect 73154 601576 73160 601588
rect 73028 601548 73160 601576
rect 73028 601536 73034 601548
rect 73154 601536 73160 601548
rect 73212 601536 73218 601588
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 72881 598927 72939 598933
rect 72881 598893 72893 598927
rect 72927 598924 72939 598927
rect 72970 598924 72976 598936
rect 72927 598896 72976 598924
rect 72927 598893 72939 598896
rect 72881 598887 72939 598893
rect 72970 598884 72976 598896
rect 73028 598884 73034 598936
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 413002 598924 413008 598936
rect 412963 598896 413008 598924
rect 413002 598884 413008 598896
rect 413060 598884 413066 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 542722 598924 542728 598936
rect 542683 598896 542728 598924
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 137738 596164 137744 596216
rect 137796 596204 137802 596216
rect 137922 596204 137928 596216
rect 137796 596176 137928 596204
rect 137796 596164 137802 596176
rect 137922 596164 137928 596176
rect 137980 596164 137986 596216
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 284018 596164 284024 596216
rect 284076 596204 284082 596216
rect 284202 596204 284208 596216
rect 284076 596176 284208 596204
rect 284076 596164 284082 596176
rect 284202 596164 284208 596176
rect 284260 596164 284266 596216
rect 347774 596164 347780 596216
rect 347832 596204 347838 596216
rect 347958 596204 347964 596216
rect 347832 596176 347964 596204
rect 347832 596164 347838 596176
rect 347958 596164 347964 596176
rect 348016 596164 348022 596216
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 477494 596164 477500 596216
rect 477552 596204 477558 596216
rect 477678 596204 477684 596216
rect 477552 596176 477684 596204
rect 477552 596164 477558 596176
rect 477678 596164 477684 596176
rect 477736 596164 477742 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 13078 594844 13084 594856
rect 3292 594816 13084 594844
rect 3292 594804 3298 594816
rect 13078 594804 13084 594816
rect 13136 594804 13142 594856
rect 476758 592016 476764 592068
rect 476816 592056 476822 592068
rect 579890 592056 579896 592068
rect 476816 592028 579896 592056
rect 476816 592016 476822 592028
rect 579890 592016 579896 592028
rect 579948 592016 579954 592068
rect 72878 589336 72884 589348
rect 72839 589308 72884 589336
rect 72878 589296 72884 589308
rect 72936 589296 72942 589348
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 413005 589339 413063 589345
rect 413005 589305 413017 589339
rect 413051 589336 413063 589339
rect 413094 589336 413100 589348
rect 413051 589308 413100 589336
rect 413051 589305 413063 589308
rect 413005 589299 413063 589305
rect 413094 589296 413100 589308
rect 413152 589296 413158 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 542725 589339 542783 589345
rect 542725 589305 542737 589339
rect 542771 589336 542783 589339
rect 542814 589336 542820 589348
rect 542771 589308 542820 589336
rect 542771 589305 542783 589308
rect 542725 589299 542783 589305
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 8018 589268 8024 589280
rect 7979 589240 8024 589268
rect 8018 589228 8024 589240
rect 8076 589228 8082 589280
rect 137738 589268 137744 589280
rect 137699 589240 137744 589268
rect 137738 589228 137744 589240
rect 137796 589228 137802 589280
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 284018 589268 284024 589280
rect 283979 589240 284024 589268
rect 284018 589228 284024 589240
rect 284076 589228 284082 589280
rect 347777 589271 347835 589277
rect 347777 589237 347789 589271
rect 347823 589268 347835 589271
rect 347866 589268 347872 589280
rect 347823 589240 347872 589268
rect 347823 589237 347835 589240
rect 347777 589231 347835 589237
rect 347866 589228 347872 589240
rect 347924 589228 347930 589280
rect 364337 589271 364395 589277
rect 364337 589237 364349 589271
rect 364383 589268 364395 589271
rect 364426 589268 364432 589280
rect 364383 589240 364432 589268
rect 364383 589237 364395 589240
rect 364337 589231 364395 589237
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 477497 589271 477555 589277
rect 477497 589237 477509 589271
rect 477543 589268 477555 589271
rect 477586 589268 477592 589280
rect 477543 589240 477592 589268
rect 477543 589237 477555 589240
rect 477497 589231 477555 589237
rect 477586 589228 477592 589240
rect 477644 589228 477650 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 413094 582468 413100 582480
rect 413020 582440 413100 582468
rect 72694 582360 72700 582412
rect 72752 582400 72758 582412
rect 72878 582400 72884 582412
rect 72752 582372 72884 582400
rect 72752 582360 72758 582372
rect 72878 582360 72884 582372
rect 72936 582360 72942 582412
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 413020 582344 413048 582440
rect 413094 582428 413100 582440
rect 413152 582428 413158 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 413002 582292 413008 582344
rect 413060 582292 413066 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 8018 579748 8024 579760
rect 7979 579720 8024 579748
rect 8018 579708 8024 579720
rect 8076 579708 8082 579760
rect 137738 579748 137744 579760
rect 137699 579720 137744 579748
rect 137738 579708 137744 579720
rect 137796 579708 137802 579760
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 284018 579748 284024 579760
rect 283979 579720 284024 579748
rect 284018 579708 284024 579720
rect 284076 579708 284082 579760
rect 347774 579640 347780 579692
rect 347832 579680 347838 579692
rect 364334 579680 364340 579692
rect 347832 579652 347877 579680
rect 364295 579652 364340 579680
rect 347832 579640 347838 579652
rect 364334 579640 364340 579652
rect 364392 579640 364398 579692
rect 477494 579680 477500 579692
rect 477455 579652 477500 579680
rect 477494 579640 477500 579652
rect 477552 579640 477558 579692
rect 489178 579640 489184 579692
rect 489236 579680 489242 579692
rect 580166 579680 580172 579692
rect 489236 579652 580172 579680
rect 489236 579640 489242 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 7926 579572 7932 579624
rect 7984 579612 7990 579624
rect 8110 579612 8116 579624
rect 7984 579584 8116 579612
rect 7984 579572 7990 579584
rect 8110 579572 8116 579584
rect 8168 579572 8174 579624
rect 72605 579615 72663 579621
rect 72605 579581 72617 579615
rect 72651 579612 72663 579615
rect 72694 579612 72700 579624
rect 72651 579584 72700 579612
rect 72651 579581 72663 579584
rect 72605 579575 72663 579581
rect 72694 579572 72700 579584
rect 72752 579572 72758 579624
rect 137557 579615 137615 579621
rect 137557 579581 137569 579615
rect 137603 579612 137615 579615
rect 137646 579612 137652 579624
rect 137603 579584 137652 579612
rect 137603 579581 137615 579584
rect 137557 579575 137615 579581
rect 137646 579572 137652 579584
rect 137704 579572 137710 579624
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 283926 579572 283932 579624
rect 283984 579612 283990 579624
rect 284110 579612 284116 579624
rect 283984 579584 284116 579612
rect 283984 579572 283990 579584
rect 284110 579572 284116 579584
rect 284168 579572 284174 579624
rect 72602 569956 72608 569968
rect 72563 569928 72608 569956
rect 72602 569916 72608 569928
rect 72660 569916 72666 569968
rect 137554 569956 137560 569968
rect 137515 569928 137560 569956
rect 137554 569916 137560 569928
rect 137612 569916 137618 569968
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 347866 569888 347872 569900
rect 347827 569860 347872 569888
rect 347866 569848 347872 569860
rect 347924 569848 347930 569900
rect 364426 569888 364432 569900
rect 364387 569860 364432 569888
rect 364426 569848 364432 569860
rect 364484 569848 364490 569900
rect 477586 569888 477592 569900
rect 477547 569860 477592 569888
rect 477586 569848 477592 569860
rect 477644 569848 477650 569900
rect 494146 569888 494152 569900
rect 494107 569860 494152 569888
rect 494146 569848 494152 569860
rect 494204 569848 494210 569900
rect 13078 567808 13084 567860
rect 13136 567848 13142 567860
rect 128998 567848 129004 567860
rect 13136 567820 129004 567848
rect 13136 567808 13142 567820
rect 128998 567808 129004 567820
rect 129056 567808 129062 567860
rect 4062 567264 4068 567316
rect 4120 567304 4126 567316
rect 11698 567304 11704 567316
rect 4120 567276 11704 567304
rect 4120 567264 4126 567276
rect 11698 567264 11704 567276
rect 11756 567264 11762 567316
rect 412726 563116 412732 563168
rect 412784 563116 412790 563168
rect 429286 563116 429292 563168
rect 429344 563116 429350 563168
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 72602 563048 72608 563100
rect 72660 563048 72666 563100
rect 137554 563048 137560 563100
rect 137612 563048 137618 563100
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 347869 563091 347927 563097
rect 347869 563057 347881 563091
rect 347915 563088 347927 563091
rect 348050 563088 348056 563100
rect 347915 563060 348056 563088
rect 347915 563057 347927 563060
rect 347869 563051 347927 563057
rect 348050 563048 348056 563060
rect 348108 563048 348114 563100
rect 364429 563091 364487 563097
rect 364429 563057 364441 563091
rect 364475 563088 364487 563091
rect 364610 563088 364616 563100
rect 364475 563060 364616 563088
rect 364475 563057 364487 563060
rect 364429 563051 364487 563057
rect 364610 563048 364616 563060
rect 364668 563048 364674 563100
rect 7926 562912 7932 562964
rect 7984 562952 7990 562964
rect 8110 562952 8116 562964
rect 7984 562924 8116 562952
rect 7984 562912 7990 562924
rect 8110 562912 8116 562924
rect 8168 562912 8174 562964
rect 72620 562952 72648 563048
rect 72694 562952 72700 562964
rect 72620 562924 72700 562952
rect 72694 562912 72700 562924
rect 72752 562912 72758 562964
rect 137572 562952 137600 563048
rect 137646 562952 137652 562964
rect 137572 562924 137652 562952
rect 137646 562912 137652 562924
rect 137704 562912 137710 562964
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 412744 563032 412772 563116
rect 429304 563032 429332 563116
rect 477589 563091 477647 563097
rect 477589 563057 477601 563091
rect 477635 563088 477647 563091
rect 477770 563088 477776 563100
rect 477635 563060 477776 563088
rect 477635 563057 477647 563060
rect 477589 563051 477647 563057
rect 477770 563048 477776 563060
rect 477828 563048 477834 563100
rect 494149 563091 494207 563097
rect 494149 563057 494161 563091
rect 494195 563088 494207 563091
rect 494330 563088 494336 563100
rect 494195 563060 494336 563088
rect 494195 563057 494207 563060
rect 494149 563051 494207 563057
rect 494330 563048 494336 563060
rect 494388 563048 494394 563100
rect 542464 563032 542492 563116
rect 559024 563032 559052 563116
rect 412726 562980 412732 563032
rect 412784 562980 412790 563032
rect 429286 562980 429292 563032
rect 429344 562980 429350 563032
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 283926 562912 283932 562964
rect 283984 562952 283990 562964
rect 284110 562952 284116 562964
rect 283984 562924 284116 562952
rect 283984 562912 283990 562924
rect 284110 562912 284116 562924
rect 284168 562912 284174 562964
rect 72694 560232 72700 560244
rect 72655 560204 72700 560232
rect 72694 560192 72700 560204
rect 72752 560192 72758 560244
rect 137646 560232 137652 560244
rect 137607 560204 137652 560232
rect 137646 560192 137652 560204
rect 137704 560192 137710 560244
rect 218974 560232 218980 560244
rect 218935 560204 218980 560232
rect 218974 560192 218980 560204
rect 219032 560192 219038 560244
rect 412726 560232 412732 560244
rect 412687 560204 412732 560232
rect 412726 560192 412732 560204
rect 412784 560192 412790 560244
rect 429286 560232 429292 560244
rect 429247 560204 429292 560232
rect 429286 560192 429292 560204
rect 429344 560192 429350 560244
rect 542446 560232 542452 560244
rect 542407 560204 542452 560232
rect 542446 560192 542452 560204
rect 542504 560192 542510 560244
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 483658 556180 483664 556232
rect 483716 556220 483722 556232
rect 580166 556220 580172 556232
rect 483716 556192 580172 556220
rect 483716 556180 483722 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 72697 550647 72755 550653
rect 72697 550613 72709 550647
rect 72743 550644 72755 550647
rect 72878 550644 72884 550656
rect 72743 550616 72884 550644
rect 72743 550613 72755 550616
rect 72697 550607 72755 550613
rect 72878 550604 72884 550616
rect 72936 550604 72942 550656
rect 137649 550647 137707 550653
rect 137649 550613 137661 550647
rect 137695 550644 137707 550647
rect 137830 550644 137836 550656
rect 137695 550616 137836 550644
rect 137695 550613 137707 550616
rect 137649 550607 137707 550613
rect 137830 550604 137836 550616
rect 137888 550604 137894 550656
rect 218977 550647 219035 550653
rect 218977 550613 218989 550647
rect 219023 550644 219035 550647
rect 219158 550644 219164 550656
rect 219023 550616 219164 550644
rect 219023 550613 219035 550616
rect 218977 550607 219035 550613
rect 219158 550604 219164 550616
rect 219216 550604 219222 550656
rect 347866 550604 347872 550656
rect 347924 550644 347930 550656
rect 348142 550644 348148 550656
rect 347924 550616 348148 550644
rect 347924 550604 347930 550616
rect 348142 550604 348148 550616
rect 348200 550604 348206 550656
rect 364426 550604 364432 550656
rect 364484 550644 364490 550656
rect 364702 550644 364708 550656
rect 364484 550616 364708 550644
rect 364484 550604 364490 550616
rect 364702 550604 364708 550616
rect 364760 550604 364766 550656
rect 412729 550647 412787 550653
rect 412729 550613 412741 550647
rect 412775 550644 412787 550647
rect 412910 550644 412916 550656
rect 412775 550616 412916 550644
rect 412775 550613 412787 550616
rect 412729 550607 412787 550613
rect 412910 550604 412916 550616
rect 412968 550604 412974 550656
rect 429289 550647 429347 550653
rect 429289 550613 429301 550647
rect 429335 550644 429347 550647
rect 429470 550644 429476 550656
rect 429335 550616 429476 550644
rect 429335 550613 429347 550616
rect 429289 550607 429347 550613
rect 429470 550604 429476 550616
rect 429528 550604 429534 550656
rect 477586 550604 477592 550656
rect 477644 550644 477650 550656
rect 477862 550644 477868 550656
rect 477644 550616 477868 550644
rect 477644 550604 477650 550616
rect 477862 550604 477868 550616
rect 477920 550604 477926 550656
rect 494146 550604 494152 550656
rect 494204 550644 494210 550656
rect 494422 550644 494428 550656
rect 494204 550616 494428 550644
rect 494204 550604 494210 550616
rect 494422 550604 494428 550616
rect 494480 550604 494486 550656
rect 542449 550647 542507 550653
rect 542449 550613 542461 550647
rect 542495 550644 542507 550647
rect 542630 550644 542636 550656
rect 542495 550616 542636 550644
rect 542495 550613 542507 550616
rect 542449 550607 542507 550613
rect 542630 550604 542636 550616
rect 542688 550604 542694 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559190 550644 559196 550656
rect 559055 550616 559196 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559190 550604 559196 550616
rect 559248 550604 559254 550656
rect 8018 550576 8024 550588
rect 7979 550548 8024 550576
rect 8018 550536 8024 550548
rect 8076 550536 8082 550588
rect 154298 550576 154304 550588
rect 154259 550548 154304 550576
rect 154298 550536 154304 550548
rect 154356 550536 154362 550588
rect 284018 550576 284024 550588
rect 283979 550548 284024 550576
rect 284018 550536 284024 550548
rect 284076 550536 284082 550588
rect 475378 545096 475384 545148
rect 475436 545136 475442 545148
rect 579890 545136 579896 545148
rect 475436 545108 579896 545136
rect 475436 545096 475442 545108
rect 579890 545096 579896 545108
rect 579948 545096 579954 545148
rect 348142 543844 348148 543856
rect 348068 543816 348148 543844
rect 8021 543779 8079 543785
rect 8021 543745 8033 543779
rect 8067 543776 8079 543779
rect 8202 543776 8208 543788
rect 8067 543748 8208 543776
rect 8067 543745 8079 543748
rect 8021 543739 8079 543745
rect 8202 543736 8208 543748
rect 8260 543736 8266 543788
rect 154301 543779 154359 543785
rect 154301 543745 154313 543779
rect 154347 543776 154359 543779
rect 154482 543776 154488 543788
rect 154347 543748 154488 543776
rect 154347 543745 154359 543748
rect 154301 543739 154359 543745
rect 154482 543736 154488 543748
rect 154540 543736 154546 543788
rect 284021 543779 284079 543785
rect 284021 543745 284033 543779
rect 284067 543776 284079 543779
rect 284202 543776 284208 543788
rect 284067 543748 284208 543776
rect 284067 543745 284079 543748
rect 284021 543739 284079 543745
rect 284202 543736 284208 543748
rect 284260 543736 284266 543788
rect 348068 543720 348096 543816
rect 348142 543804 348148 543816
rect 348200 543804 348206 543856
rect 364702 543844 364708 543856
rect 364628 543816 364708 543844
rect 364628 543720 364656 543816
rect 364702 543804 364708 543816
rect 364760 543804 364766 543856
rect 477862 543844 477868 543856
rect 477788 543816 477868 543844
rect 477788 543720 477816 543816
rect 477862 543804 477868 543816
rect 477920 543804 477926 543856
rect 494422 543844 494428 543856
rect 494348 543816 494428 543844
rect 494348 543720 494376 543816
rect 494422 543804 494428 543816
rect 494480 543804 494486 543856
rect 348050 543668 348056 543720
rect 348108 543668 348114 543720
rect 364610 543668 364616 543720
rect 364668 543668 364674 543720
rect 477770 543668 477776 543720
rect 477828 543668 477834 543720
rect 494330 543668 494336 543720
rect 494388 543668 494394 543720
rect 72694 543600 72700 543652
rect 72752 543640 72758 543652
rect 72878 543640 72884 543652
rect 72752 543612 72884 543640
rect 72752 543600 72758 543612
rect 72878 543600 72884 543612
rect 72936 543600 72942 543652
rect 137646 543600 137652 543652
rect 137704 543640 137710 543652
rect 137830 543640 137836 543652
rect 137704 543612 137836 543640
rect 137704 543600 137710 543612
rect 137830 543600 137836 543612
rect 137888 543600 137894 543652
rect 218974 543600 218980 543652
rect 219032 543640 219038 543652
rect 219158 543640 219164 543652
rect 219032 543612 219164 543640
rect 219032 543600 219038 543612
rect 219158 543600 219164 543612
rect 219216 543600 219222 543652
rect 412726 543600 412732 543652
rect 412784 543640 412790 543652
rect 412910 543640 412916 543652
rect 412784 543612 412916 543640
rect 412784 543600 412790 543612
rect 412910 543600 412916 543612
rect 412968 543600 412974 543652
rect 429286 543600 429292 543652
rect 429344 543640 429350 543652
rect 429470 543640 429476 543652
rect 429344 543612 429476 543640
rect 429344 543600 429350 543612
rect 429470 543600 429476 543612
rect 429528 543600 429534 543652
rect 542446 543600 542452 543652
rect 542504 543640 542510 543652
rect 542630 543640 542636 543652
rect 542504 543612 542636 543640
rect 542504 543600 542510 543612
rect 542630 543600 542636 543612
rect 542688 543600 542694 543652
rect 559006 543600 559012 543652
rect 559064 543640 559070 543652
rect 559190 543640 559196 543652
rect 559064 543612 559196 543640
rect 559064 543600 559070 543612
rect 559190 543600 559196 543612
rect 559248 543600 559254 543652
rect 3694 538228 3700 538280
rect 3752 538268 3758 538280
rect 15838 538268 15844 538280
rect 3752 538240 15844 538268
rect 3752 538228 3758 538240
rect 15838 538228 15844 538240
rect 15896 538228 15902 538280
rect 72694 534012 72700 534064
rect 72752 534052 72758 534064
rect 72878 534052 72884 534064
rect 72752 534024 72884 534052
rect 72752 534012 72758 534024
rect 72878 534012 72884 534024
rect 72936 534012 72942 534064
rect 137646 534012 137652 534064
rect 137704 534052 137710 534064
rect 137830 534052 137836 534064
rect 137704 534024 137836 534052
rect 137704 534012 137710 534024
rect 137830 534012 137836 534024
rect 137888 534012 137894 534064
rect 218974 534012 218980 534064
rect 219032 534052 219038 534064
rect 219158 534052 219164 534064
rect 219032 534024 219164 534052
rect 219032 534012 219038 534024
rect 219158 534012 219164 534024
rect 219216 534012 219222 534064
rect 485038 532720 485044 532772
rect 485096 532760 485102 532772
rect 580166 532760 580172 532772
rect 485096 532732 580172 532760
rect 485096 532720 485102 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 7926 531292 7932 531344
rect 7984 531332 7990 531344
rect 8018 531332 8024 531344
rect 7984 531304 8024 531332
rect 7984 531292 7990 531304
rect 8018 531292 8024 531304
rect 8076 531292 8082 531344
rect 154206 531292 154212 531344
rect 154264 531332 154270 531344
rect 154298 531332 154304 531344
rect 154264 531304 154304 531332
rect 154264 531292 154270 531304
rect 154298 531292 154304 531304
rect 154356 531292 154362 531344
rect 347866 531292 347872 531344
rect 347924 531332 347930 531344
rect 348142 531332 348148 531344
rect 347924 531304 348148 531332
rect 347924 531292 347930 531304
rect 348142 531292 348148 531304
rect 348200 531292 348206 531344
rect 364426 531292 364432 531344
rect 364484 531332 364490 531344
rect 364702 531332 364708 531344
rect 364484 531304 364708 531332
rect 364484 531292 364490 531304
rect 364702 531292 364708 531304
rect 364760 531292 364766 531344
rect 477586 531292 477592 531344
rect 477644 531332 477650 531344
rect 477862 531332 477868 531344
rect 477644 531304 477868 531332
rect 477644 531292 477650 531304
rect 477862 531292 477868 531304
rect 477920 531292 477926 531344
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 72786 524464 72792 524476
rect 72747 524436 72792 524464
rect 72786 524424 72792 524436
rect 72844 524424 72850 524476
rect 137738 524464 137744 524476
rect 137699 524436 137744 524464
rect 137738 524424 137744 524436
rect 137796 524424 137802 524476
rect 154298 524424 154304 524476
rect 154356 524424 154362 524476
rect 219066 524464 219072 524476
rect 219027 524436 219072 524464
rect 219066 524424 219072 524436
rect 219124 524424 219130 524476
rect 8110 524288 8116 524340
rect 8168 524328 8174 524340
rect 8294 524328 8300 524340
rect 8168 524300 8300 524328
rect 8168 524288 8174 524300
rect 8294 524288 8300 524300
rect 8352 524288 8358 524340
rect 154316 524328 154344 524424
rect 154390 524328 154396 524340
rect 154316 524300 154396 524328
rect 154390 524288 154396 524300
rect 154448 524288 154454 524340
rect 284110 524288 284116 524340
rect 284168 524328 284174 524340
rect 284294 524328 284300 524340
rect 284168 524300 284300 524328
rect 284168 524288 284174 524300
rect 284294 524288 284300 524300
rect 284352 524288 284358 524340
rect 72786 521676 72792 521688
rect 72747 521648 72792 521676
rect 72786 521636 72792 521648
rect 72844 521636 72850 521688
rect 137738 521676 137744 521688
rect 137699 521648 137744 521676
rect 137738 521636 137744 521648
rect 137796 521636 137802 521688
rect 219066 521676 219072 521688
rect 219027 521648 219072 521676
rect 219066 521636 219072 521648
rect 219124 521636 219130 521688
rect 347958 521636 347964 521688
rect 348016 521676 348022 521688
rect 348142 521676 348148 521688
rect 348016 521648 348148 521676
rect 348016 521636 348022 521648
rect 348142 521636 348148 521648
rect 348200 521636 348206 521688
rect 364518 521636 364524 521688
rect 364576 521676 364582 521688
rect 364702 521676 364708 521688
rect 364576 521648 364708 521676
rect 364576 521636 364582 521648
rect 364702 521636 364708 521648
rect 364760 521636 364766 521688
rect 477678 521636 477684 521688
rect 477736 521676 477742 521688
rect 477862 521676 477868 521688
rect 477736 521648 477868 521676
rect 477736 521636 477742 521648
rect 477862 521636 477868 521648
rect 477920 521636 477926 521688
rect 494238 521636 494244 521688
rect 494296 521676 494302 521688
rect 494422 521676 494428 521688
rect 494296 521648 494428 521676
rect 494296 521636 494302 521648
rect 494422 521636 494428 521648
rect 494480 521636 494486 521688
rect 284110 516060 284116 516112
rect 284168 516100 284174 516112
rect 291102 516100 291108 516112
rect 284168 516072 291108 516100
rect 284168 516060 284174 516072
rect 291102 516060 291108 516072
rect 291160 516060 291166 516112
rect 106182 515720 106188 515772
rect 106240 515760 106246 515772
rect 196802 515760 196808 515772
rect 106240 515732 196808 515760
rect 106240 515720 106246 515732
rect 196802 515720 196808 515732
rect 196860 515720 196866 515772
rect 385494 515720 385500 515772
rect 385552 515760 385558 515772
rect 462314 515760 462320 515772
rect 385552 515732 462320 515760
rect 385552 515720 385558 515732
rect 462314 515720 462320 515732
rect 462372 515720 462378 515772
rect 89622 515652 89628 515704
rect 89680 515692 89686 515704
rect 185026 515692 185032 515704
rect 89680 515664 185032 515692
rect 89680 515652 89686 515664
rect 185026 515652 185032 515664
rect 185084 515652 185090 515704
rect 397270 515652 397276 515704
rect 397328 515692 397334 515704
rect 477678 515692 477684 515704
rect 397328 515664 477684 515692
rect 397328 515652 397334 515664
rect 477678 515652 477684 515664
rect 477736 515652 477742 515704
rect 72786 515584 72792 515636
rect 72844 515624 72850 515636
rect 173250 515624 173256 515636
rect 72844 515596 173256 515624
rect 72844 515584 72850 515596
rect 173250 515584 173256 515596
rect 173308 515584 173314 515636
rect 202782 515584 202788 515636
rect 202840 515624 202846 515636
rect 243998 515624 244004 515636
rect 202840 515596 244004 515624
rect 202840 515584 202846 515596
rect 243998 515584 244004 515596
rect 244056 515584 244062 515636
rect 409046 515584 409052 515636
rect 409104 515624 409110 515636
rect 494238 515624 494244 515636
rect 409104 515596 494244 515624
rect 409104 515584 409110 515596
rect 494238 515584 494244 515596
rect 494296 515584 494302 515636
rect 41322 515516 41328 515568
rect 41380 515556 41386 515568
rect 161474 515556 161480 515568
rect 41380 515528 161480 515556
rect 41380 515516 41386 515528
rect 161474 515516 161480 515528
rect 161532 515516 161538 515568
rect 171042 515516 171048 515568
rect 171100 515556 171106 515568
rect 232222 515556 232228 515568
rect 171100 515528 232228 515556
rect 171100 515516 171106 515528
rect 232222 515516 232228 515528
rect 232280 515516 232286 515568
rect 350074 515516 350080 515568
rect 350132 515556 350138 515568
rect 397454 515556 397460 515568
rect 350132 515528 397460 515556
rect 350132 515516 350138 515528
rect 397454 515516 397460 515528
rect 397512 515516 397518 515568
rect 420822 515516 420828 515568
rect 420880 515556 420886 515568
rect 527174 515556 527180 515568
rect 420880 515528 527180 515556
rect 420880 515516 420886 515528
rect 527174 515516 527180 515528
rect 527232 515516 527238 515568
rect 24762 515448 24768 515500
rect 24820 515488 24826 515500
rect 149698 515488 149704 515500
rect 24820 515460 149704 515488
rect 24820 515448 24826 515460
rect 149698 515448 149704 515460
rect 149756 515448 149762 515500
rect 154390 515448 154396 515500
rect 154448 515488 154454 515500
rect 220446 515488 220452 515500
rect 154448 515460 220452 515488
rect 154448 515448 154454 515460
rect 220446 515448 220452 515460
rect 220504 515448 220510 515500
rect 235902 515448 235908 515500
rect 235960 515488 235966 515500
rect 267550 515488 267556 515500
rect 235960 515460 267556 515488
rect 235960 515448 235966 515460
rect 267550 515448 267556 515460
rect 267608 515448 267614 515500
rect 326522 515448 326528 515500
rect 326580 515488 326586 515500
rect 347958 515488 347964 515500
rect 326580 515460 347964 515488
rect 326580 515448 326586 515460
rect 347958 515448 347964 515460
rect 348016 515448 348022 515500
rect 361850 515448 361856 515500
rect 361908 515488 361914 515500
rect 412910 515488 412916 515500
rect 361908 515460 412916 515488
rect 361908 515448 361914 515460
rect 412910 515448 412916 515460
rect 412968 515448 412974 515500
rect 432598 515448 432604 515500
rect 432656 515488 432662 515500
rect 542630 515488 542636 515500
rect 432656 515460 542636 515488
rect 432656 515448 432662 515460
rect 542630 515448 542636 515460
rect 542688 515448 542694 515500
rect 8110 515380 8116 515432
rect 8168 515420 8174 515432
rect 137922 515420 137928 515432
rect 8168 515392 137928 515420
rect 8168 515380 8174 515392
rect 137922 515380 137928 515392
rect 137980 515380 137986 515432
rect 138014 515380 138020 515432
rect 138072 515420 138078 515432
rect 208578 515420 208584 515432
rect 138072 515392 208584 515420
rect 138072 515380 138078 515392
rect 208578 515380 208584 515392
rect 208636 515380 208642 515432
rect 219066 515380 219072 515432
rect 219124 515420 219130 515432
rect 255774 515420 255780 515432
rect 219124 515392 255780 515420
rect 219124 515380 219130 515392
rect 255774 515380 255780 515392
rect 255832 515380 255838 515432
rect 267642 515380 267648 515432
rect 267700 515420 267706 515432
rect 279326 515420 279332 515432
rect 267700 515392 279332 515420
rect 267700 515380 267706 515392
rect 279326 515380 279332 515392
rect 279384 515380 279390 515432
rect 314746 515380 314752 515432
rect 314804 515420 314810 515432
rect 331214 515420 331220 515432
rect 314804 515392 331220 515420
rect 314804 515380 314810 515392
rect 331214 515380 331220 515392
rect 331272 515380 331278 515432
rect 338298 515380 338304 515432
rect 338356 515420 338362 515432
rect 364518 515420 364524 515432
rect 338356 515392 364524 515420
rect 338356 515380 338362 515392
rect 364518 515380 364524 515392
rect 364576 515380 364582 515432
rect 373626 515380 373632 515432
rect 373684 515420 373690 515432
rect 429470 515420 429476 515432
rect 373684 515392 429476 515420
rect 373684 515380 373690 515392
rect 429470 515380 429476 515392
rect 429528 515380 429534 515432
rect 444374 515380 444380 515432
rect 444432 515420 444438 515432
rect 559190 515420 559196 515432
rect 444432 515392 559196 515420
rect 444432 515380 444438 515392
rect 559190 515380 559196 515392
rect 559248 515380 559254 515432
rect 300762 514836 300768 514888
rect 300820 514876 300826 514888
rect 302970 514876 302976 514888
rect 300820 514848 302976 514876
rect 300820 514836 300826 514848
rect 302970 514836 302976 514848
rect 303028 514836 303034 514888
rect 2866 509260 2872 509312
rect 2924 509300 2930 509312
rect 13078 509300 13084 509312
rect 2924 509272 13084 509300
rect 2924 509260 2930 509272
rect 13078 509260 13084 509272
rect 13136 509260 13142 509312
rect 462958 509260 462964 509312
rect 463016 509300 463022 509312
rect 580166 509300 580172 509312
rect 463016 509272 580172 509300
rect 463016 509260 463022 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 8938 509192 8944 509244
rect 8996 509232 9002 509244
rect 128354 509232 128360 509244
rect 8996 509204 128360 509232
rect 8996 509192 9002 509204
rect 128354 509192 128360 509204
rect 128412 509192 128418 509244
rect 453206 509192 453212 509244
rect 453264 509232 453270 509244
rect 472618 509232 472624 509244
rect 453264 509204 472624 509232
rect 453264 509192 453270 509204
rect 472618 509192 472624 509204
rect 472676 509192 472682 509244
rect 17218 502256 17224 502308
rect 17276 502296 17282 502308
rect 128354 502296 128360 502308
rect 17276 502268 128360 502296
rect 17276 502256 17282 502268
rect 128354 502256 128360 502268
rect 128412 502256 128418 502308
rect 453390 502256 453396 502308
rect 453448 502296 453454 502308
rect 580258 502296 580264 502308
rect 453448 502268 580264 502296
rect 453448 502256 453454 502268
rect 580258 502256 580264 502268
rect 580316 502256 580322 502308
rect 460198 498176 460204 498228
rect 460256 498216 460262 498228
rect 580166 498216 580172 498228
rect 460256 498188 580172 498216
rect 460256 498176 460262 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 453942 495388 453948 495440
rect 454000 495428 454006 495440
rect 490558 495428 490564 495440
rect 454000 495400 490564 495428
rect 454000 495388 454006 495400
rect 490558 495388 490564 495400
rect 490616 495388 490622 495440
rect 14458 493960 14464 494012
rect 14516 494000 14522 494012
rect 128354 494000 128360 494012
rect 14516 493972 128360 494000
rect 14516 493960 14522 493972
rect 128354 493960 128360 493972
rect 128412 493960 128418 494012
rect 453758 488452 453764 488504
rect 453816 488492 453822 488504
rect 471238 488492 471244 488504
rect 453816 488464 471244 488492
rect 453816 488452 453822 488464
rect 471238 488452 471244 488464
rect 471296 488452 471302 488504
rect 456058 485800 456064 485852
rect 456116 485840 456122 485852
rect 580166 485840 580172 485852
rect 456116 485812 580172 485840
rect 456116 485800 456122 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 10318 485732 10324 485784
rect 10376 485772 10382 485784
rect 128354 485772 128360 485784
rect 10376 485744 128360 485772
rect 10376 485732 10382 485744
rect 128354 485732 128360 485744
rect 128412 485732 128418 485784
rect 453758 481584 453764 481636
rect 453816 481624 453822 481636
rect 580350 481624 580356 481636
rect 453816 481596 580356 481624
rect 453816 481584 453822 481596
rect 580350 481584 580356 481596
rect 580408 481584 580414 481636
rect 3326 480224 3332 480276
rect 3384 480264 3390 480276
rect 8938 480264 8944 480276
rect 3384 480236 8944 480264
rect 3384 480224 3390 480236
rect 8938 480224 8944 480236
rect 8996 480224 9002 480276
rect 19978 478796 19984 478848
rect 20036 478836 20042 478848
rect 128354 478836 128360 478848
rect 20036 478808 128360 478836
rect 20036 478796 20042 478808
rect 128354 478796 128360 478808
rect 128412 478796 128418 478848
rect 453942 473288 453948 473340
rect 454000 473328 454006 473340
rect 479518 473328 479524 473340
rect 454000 473300 479524 473328
rect 454000 473288 454006 473300
rect 479518 473288 479524 473300
rect 479576 473288 479582 473340
rect 452746 466352 452752 466404
rect 452804 466392 452810 466404
rect 467098 466392 467104 466404
rect 452804 466364 467104 466392
rect 452804 466352 452810 466364
rect 467098 466352 467104 466364
rect 467156 466352 467162 466404
rect 11698 463632 11704 463684
rect 11756 463672 11762 463684
rect 128354 463672 128360 463684
rect 11756 463644 128360 463672
rect 11756 463632 11762 463644
rect 128354 463632 128360 463644
rect 128412 463632 128418 463684
rect 454678 462340 454684 462392
rect 454736 462380 454742 462392
rect 580166 462380 580172 462392
rect 454736 462352 580172 462380
rect 454736 462340 454742 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 453390 459484 453396 459536
rect 453448 459524 453454 459536
rect 476758 459524 476764 459536
rect 453448 459496 476764 459524
rect 453448 459484 453454 459496
rect 476758 459484 476764 459496
rect 476816 459484 476822 459536
rect 3418 455336 3424 455388
rect 3476 455376 3482 455388
rect 128354 455376 128360 455388
rect 3476 455348 128360 455376
rect 3476 455336 3482 455348
rect 128354 455336 128360 455348
rect 128412 455336 128418 455388
rect 453942 452548 453948 452600
rect 454000 452588 454006 452600
rect 489178 452588 489184 452600
rect 454000 452560 489184 452588
rect 454000 452548 454006 452560
rect 489178 452548 489184 452560
rect 489236 452548 489242 452600
rect 3142 451256 3148 451308
rect 3200 451296 3206 451308
rect 58618 451296 58624 451308
rect 3200 451268 58624 451296
rect 3200 451256 3206 451268
rect 58618 451256 58624 451268
rect 58676 451256 58682 451308
rect 15838 448468 15844 448520
rect 15896 448508 15902 448520
rect 128354 448508 128360 448520
rect 15896 448480 128360 448508
rect 15896 448468 15902 448480
rect 128354 448468 128360 448480
rect 128412 448468 128418 448520
rect 453666 445680 453672 445732
rect 453724 445720 453730 445732
rect 483658 445720 483664 445732
rect 453724 445692 483664 445720
rect 453724 445680 453730 445692
rect 483658 445680 483664 445692
rect 483716 445680 483722 445732
rect 13078 440172 13084 440224
rect 13136 440212 13142 440224
rect 128354 440212 128360 440224
rect 13136 440184 128360 440212
rect 13136 440172 13142 440184
rect 128354 440172 128360 440184
rect 128412 440172 128418 440224
rect 453298 438880 453304 438932
rect 453356 438920 453362 438932
rect 579890 438920 579896 438932
rect 453356 438892 579896 438920
rect 453356 438880 453362 438892
rect 579890 438880 579896 438892
rect 579948 438880 579954 438932
rect 453758 438812 453764 438864
rect 453816 438852 453822 438864
rect 475378 438852 475384 438864
rect 453816 438824 475384 438852
rect 453816 438812 453822 438824
rect 475378 438812 475384 438824
rect 475436 438812 475442 438864
rect 3510 433236 3516 433288
rect 3568 433276 3574 433288
rect 128354 433276 128360 433288
rect 3568 433248 128360 433276
rect 3568 433236 3574 433248
rect 128354 433236 128360 433248
rect 128412 433236 128418 433288
rect 453942 430516 453948 430568
rect 454000 430556 454006 430568
rect 485038 430556 485044 430568
rect 454000 430528 485044 430556
rect 454000 430516 454006 430528
rect 485038 430516 485044 430528
rect 485096 430516 485102 430568
rect 8938 425008 8944 425060
rect 8996 425048 9002 425060
rect 128354 425048 128360 425060
rect 8996 425020 128360 425048
rect 8996 425008 9002 425020
rect 128354 425008 128360 425020
rect 128412 425008 128418 425060
rect 453942 423580 453948 423632
rect 454000 423620 454006 423632
rect 462958 423620 462964 423632
rect 454000 423592 462964 423620
rect 454000 423580 454006 423592
rect 462958 423580 462964 423592
rect 463016 423580 463022 423632
rect 58618 418072 58624 418124
rect 58676 418112 58682 418124
rect 128354 418112 128360 418124
rect 58676 418084 128360 418112
rect 58676 418072 58682 418084
rect 128354 418072 128360 418084
rect 128412 418072 128418 418124
rect 453942 416372 453948 416424
rect 454000 416412 454006 416424
rect 460198 416412 460204 416424
rect 454000 416384 460204 416412
rect 454000 416372 454006 416384
rect 460198 416372 460204 416384
rect 460256 416372 460262 416424
rect 542998 414672 543004 414724
rect 543056 414712 543062 414724
rect 580166 414712 580172 414724
rect 543056 414684 580172 414712
rect 543056 414672 543062 414684
rect 580166 414672 580172 414684
rect 580224 414672 580230 414724
rect 3418 409776 3424 409828
rect 3476 409816 3482 409828
rect 128354 409816 128360 409828
rect 3476 409788 128360 409816
rect 3476 409776 3482 409788
rect 128354 409776 128360 409788
rect 128412 409776 128418 409828
rect 453390 409368 453396 409420
rect 453448 409408 453454 409420
rect 456058 409408 456064 409420
rect 453448 409380 456064 409408
rect 453448 409368 453454 409380
rect 456058 409368 456064 409380
rect 456116 409368 456122 409420
rect 3510 402908 3516 402960
rect 3568 402948 3574 402960
rect 128354 402948 128360 402960
rect 3568 402920 128360 402948
rect 3568 402908 3574 402920
rect 128354 402908 128360 402920
rect 128412 402908 128418 402960
rect 452838 402500 452844 402552
rect 452896 402540 452902 402552
rect 454678 402540 454684 402552
rect 452896 402512 454684 402540
rect 452896 402500 452902 402512
rect 454678 402500 454684 402512
rect 454736 402500 454742 402552
rect 453758 395972 453764 396024
rect 453816 396012 453822 396024
rect 580258 396012 580264 396024
rect 453816 395984 580264 396012
rect 453816 395972 453822 395984
rect 580258 395972 580264 395984
rect 580316 395972 580322 396024
rect 3418 394612 3424 394664
rect 3476 394652 3482 394664
rect 128354 394652 128360 394664
rect 3476 394624 128360 394652
rect 3476 394612 3482 394624
rect 128354 394612 128360 394624
rect 128412 394612 128418 394664
rect 454678 391960 454684 392012
rect 454736 392000 454742 392012
rect 580166 392000 580172 392012
rect 454736 391972 580172 392000
rect 454736 391960 454742 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 128998 380848 129004 380860
rect 3292 380820 129004 380848
rect 3292 380808 3298 380820
rect 128998 380808 129004 380820
rect 129056 380808 129062 380860
rect 453942 380808 453948 380860
rect 454000 380848 454006 380860
rect 542998 380848 543004 380860
rect 454000 380820 543004 380848
rect 454000 380808 454006 380820
rect 542998 380808 543004 380820
rect 543056 380808 543062 380860
rect 453390 373940 453396 373992
rect 453448 373980 453454 373992
rect 580350 373980 580356 373992
rect 453448 373952 580356 373980
rect 453448 373940 453454 373952
rect 580350 373940 580356 373952
rect 580408 373940 580414 373992
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 128998 367044 129004 367056
rect 3200 367016 129004 367044
rect 3200 367004 3206 367016
rect 128998 367004 129004 367016
rect 129056 367004 129062 367056
rect 452654 367004 452660 367056
rect 452712 367044 452718 367056
rect 454678 367044 454684 367056
rect 452712 367016 454684 367044
rect 452712 367004 452718 367016
rect 454678 367004 454684 367016
rect 454736 367004 454742 367056
rect 453942 360136 453948 360188
rect 454000 360176 454006 360188
rect 580258 360176 580264 360188
rect 454000 360148 580264 360176
rect 454000 360136 454006 360148
rect 580258 360136 580264 360148
rect 580316 360136 580322 360188
rect 453758 353200 453764 353252
rect 453816 353240 453822 353252
rect 580258 353240 580264 353252
rect 453816 353212 580264 353240
rect 453816 353200 453822 353212
rect 580258 353200 580264 353212
rect 580316 353200 580322 353252
rect 8938 347760 8944 347812
rect 8996 347800 9002 347812
rect 128354 347800 128360 347812
rect 8996 347772 128360 347800
rect 8996 347760 9002 347772
rect 128354 347760 128360 347772
rect 128412 347760 128418 347812
rect 453942 345652 453948 345704
rect 454000 345692 454006 345704
rect 580166 345692 580172 345704
rect 454000 345664 580172 345692
rect 454000 345652 454006 345664
rect 580166 345652 580172 345664
rect 580224 345652 580230 345704
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 129274 338076 129280 338088
rect 3476 338048 129280 338076
rect 3476 338036 3482 338048
rect 129274 338036 129280 338048
rect 129332 338036 129338 338088
rect 13078 332596 13084 332648
rect 13136 332636 13142 332648
rect 128354 332636 128360 332648
rect 13136 332608 128360 332636
rect 13136 332596 13142 332608
rect 128354 332596 128360 332608
rect 128412 332596 128418 332648
rect 11698 324300 11704 324352
rect 11756 324340 11762 324352
rect 128354 324340 128360 324352
rect 11756 324312 128360 324340
rect 11756 324300 11762 324312
rect 128354 324300 128360 324312
rect 128412 324300 128418 324352
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 128998 324272 129004 324284
rect 3292 324244 129004 324272
rect 3292 324232 3298 324244
rect 128998 324232 129004 324244
rect 129056 324232 129062 324284
rect 453482 322872 453488 322924
rect 453540 322912 453546 322924
rect 580166 322912 580172 322924
rect 453540 322884 580172 322912
rect 453540 322872 453546 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 453390 311788 453396 311840
rect 453448 311828 453454 311840
rect 580166 311828 580172 311840
rect 453448 311800 580172 311828
rect 453448 311788 453454 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 15838 309136 15844 309188
rect 15896 309176 15902 309188
rect 128354 309176 128360 309188
rect 15896 309148 128360 309176
rect 15896 309136 15902 309148
rect 128354 309136 128360 309148
rect 128412 309136 128418 309188
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 129182 309108 129188 309120
rect 3384 309080 129188 309108
rect 3384 309068 3390 309080
rect 129182 309068 129188 309080
rect 129240 309068 129246 309120
rect 452930 302336 452936 302388
rect 452988 302376 452994 302388
rect 454678 302376 454684 302388
rect 452988 302348 454684 302376
rect 452988 302336 452994 302348
rect 454678 302336 454684 302348
rect 454736 302336 454742 302388
rect 10318 302200 10324 302252
rect 10376 302240 10382 302252
rect 128354 302240 128360 302252
rect 10376 302212 128360 302240
rect 10376 302200 10382 302212
rect 128354 302200 128360 302212
rect 128412 302200 128418 302252
rect 453298 299412 453304 299464
rect 453356 299452 453362 299464
rect 579798 299452 579804 299464
rect 453356 299424 579804 299452
rect 453356 299412 453362 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 3510 294856 3516 294908
rect 3568 294896 3574 294908
rect 8938 294896 8944 294908
rect 3568 294868 8944 294896
rect 3568 294856 3574 294868
rect 8938 294856 8944 294868
rect 8996 294856 9002 294908
rect 17218 287036 17224 287088
rect 17276 287076 17282 287088
rect 128354 287076 128360 287088
rect 17276 287048 128360 287076
rect 17276 287036 17282 287048
rect 128354 287036 128360 287048
rect 128412 287036 128418 287088
rect 453022 280168 453028 280220
rect 453080 280208 453086 280220
rect 456058 280208 456064 280220
rect 453080 280180 456064 280208
rect 453080 280168 453086 280180
rect 456058 280168 456064 280180
rect 456116 280168 456122 280220
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 129090 280140 129096 280152
rect 3476 280112 129096 280140
rect 3476 280100 3482 280112
rect 129090 280100 129096 280112
rect 129148 280100 129154 280152
rect 126238 278740 126244 278792
rect 126296 278780 126302 278792
rect 129090 278780 129096 278792
rect 126296 278752 129096 278780
rect 126296 278740 126302 278752
rect 129090 278740 129096 278752
rect 129148 278740 129154 278792
rect 453574 275952 453580 276004
rect 453632 275992 453638 276004
rect 580166 275992 580172 276004
rect 453632 275964 580172 275992
rect 453632 275952 453638 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3142 266296 3148 266348
rect 3200 266336 3206 266348
rect 13078 266336 13084 266348
rect 3200 266308 13084 266336
rect 3200 266296 3206 266308
rect 13078 266296 13084 266308
rect 13136 266296 13142 266348
rect 453482 264868 453488 264920
rect 453540 264908 453546 264920
rect 580166 264908 580172 264920
rect 453540 264880 580172 264908
rect 453540 264868 453546 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 13078 263576 13084 263628
rect 13136 263616 13142 263628
rect 128354 263616 128360 263628
rect 13136 263588 128360 263616
rect 13136 263576 13142 263588
rect 128354 263576 128360 263588
rect 128412 263576 128418 263628
rect 453942 259428 453948 259480
rect 454000 259468 454006 259480
rect 471238 259468 471244 259480
rect 454000 259440 471244 259468
rect 454000 259428 454006 259440
rect 471238 259428 471244 259440
rect 471296 259428 471302 259480
rect 14458 256708 14464 256760
rect 14516 256748 14522 256760
rect 128354 256748 128360 256760
rect 14516 256720 128360 256748
rect 14516 256708 14522 256720
rect 128354 256708 128360 256720
rect 128412 256708 128418 256760
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 11698 252532 11704 252544
rect 3476 252504 11704 252532
rect 3476 252492 3482 252504
rect 11698 252492 11704 252504
rect 11756 252492 11762 252544
rect 454678 252492 454684 252544
rect 454736 252532 454742 252544
rect 579798 252532 579804 252544
rect 454736 252504 579804 252532
rect 454736 252492 454742 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 452838 250452 452844 250504
rect 452896 250492 452902 250504
rect 479518 250492 479524 250504
rect 452896 250464 479524 250492
rect 452896 250452 452902 250464
rect 479518 250452 479524 250464
rect 479576 250452 479582 250504
rect 19978 241476 19984 241528
rect 20036 241516 20042 241528
rect 128354 241516 128360 241528
rect 20036 241488 128360 241516
rect 20036 241476 20042 241488
rect 128354 241476 128360 241488
rect 128412 241476 128418 241528
rect 453942 237396 453948 237448
rect 454000 237436 454006 237448
rect 469858 237436 469864 237448
rect 454000 237408 469864 237436
rect 454000 237396 454006 237408
rect 469858 237396 469864 237408
rect 469916 237396 469922 237448
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 128998 237368 129004 237380
rect 3476 237340 129004 237368
rect 3476 237328 3482 237340
rect 128998 237328 129004 237340
rect 129056 237328 129062 237380
rect 8938 233248 8944 233300
rect 8996 233288 9002 233300
rect 128354 233288 128360 233300
rect 8996 233260 128360 233288
rect 8996 233248 9002 233260
rect 128354 233248 128360 233260
rect 128412 233248 128418 233300
rect 453114 230460 453120 230512
rect 453172 230500 453178 230512
rect 472618 230500 472624 230512
rect 453172 230472 472624 230500
rect 453172 230460 453178 230472
rect 472618 230460 472624 230472
rect 472676 230460 472682 230512
rect 453390 229032 453396 229084
rect 453448 229072 453454 229084
rect 580166 229072 580172 229084
rect 453448 229044 580172 229072
rect 453448 229032 453454 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 15838 223564 15844 223576
rect 3200 223536 15844 223564
rect 3200 223524 3206 223536
rect 15838 223524 15844 223536
rect 15896 223524 15902 223576
rect 15838 218016 15844 218068
rect 15896 218056 15902 218068
rect 128354 218056 128360 218068
rect 15896 218028 128360 218056
rect 15896 218016 15902 218028
rect 128354 218016 128360 218028
rect 128412 218016 128418 218068
rect 453298 217948 453304 218000
rect 453356 217988 453362 218000
rect 580166 217988 580172 218000
rect 453356 217960 580172 217988
rect 453356 217948 453362 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 452930 216792 452936 216844
rect 452988 216832 452994 216844
rect 454678 216832 454684 216844
rect 452988 216804 454684 216832
rect 452988 216792 452994 216804
rect 454678 216792 454684 216804
rect 454736 216792 454742 216844
rect 11698 211148 11704 211200
rect 11756 211188 11762 211200
rect 128354 211188 128360 211200
rect 11756 211160 128360 211188
rect 11756 211148 11762 211160
rect 128354 211148 128360 211160
rect 128412 211148 128418 211200
rect 453942 209788 453948 209840
rect 454000 209828 454006 209840
rect 478138 209828 478144 209840
rect 454000 209800 478144 209828
rect 454000 209788 454006 209800
rect 478138 209788 478144 209800
rect 478196 209788 478202 209840
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 10318 208332 10324 208344
rect 3476 208304 10324 208332
rect 3476 208292 3482 208304
rect 10318 208292 10324 208304
rect 10376 208292 10382 208344
rect 456058 205572 456064 205624
rect 456116 205612 456122 205624
rect 579798 205612 579804 205624
rect 456116 205584 579804 205612
rect 456116 205572 456122 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 10318 194556 10324 194608
rect 10376 194596 10382 194608
rect 128630 194596 128636 194608
rect 10376 194568 128636 194596
rect 10376 194556 10382 194568
rect 128630 194556 128636 194568
rect 128688 194556 128694 194608
rect 453942 194556 453948 194608
rect 454000 194596 454006 194608
rect 483658 194596 483664 194608
rect 454000 194568 483664 194596
rect 454000 194556 454006 194568
rect 483658 194556 483664 194568
rect 483716 194556 483722 194608
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 129366 194528 129372 194540
rect 3200 194500 129372 194528
rect 3200 194488 3206 194500
rect 129366 194488 129372 194500
rect 129424 194488 129430 194540
rect 295610 190340 295616 190392
rect 295668 190380 295674 190392
rect 296530 190380 296536 190392
rect 295668 190352 296536 190380
rect 295668 190340 295674 190352
rect 296530 190340 296536 190352
rect 296588 190340 296594 190392
rect 303890 190340 303896 190392
rect 303948 190380 303954 190392
rect 304810 190380 304816 190392
rect 303948 190352 304816 190380
rect 303948 190340 303954 190352
rect 304810 190340 304816 190352
rect 304868 190340 304874 190392
rect 439130 190340 439136 190392
rect 439188 190380 439194 190392
rect 440050 190380 440056 190392
rect 439188 190352 440056 190380
rect 439188 190340 439194 190352
rect 440050 190340 440056 190352
rect 440108 190340 440114 190392
rect 168650 190272 168656 190324
rect 168708 190312 168714 190324
rect 169570 190312 169576 190324
rect 168708 190284 169576 190312
rect 168708 190272 168714 190284
rect 169570 190272 169576 190284
rect 169628 190272 169634 190324
rect 320358 190272 320364 190324
rect 320416 190312 320422 190324
rect 321370 190312 321376 190324
rect 320416 190284 321376 190312
rect 320416 190272 320422 190284
rect 321370 190272 321376 190284
rect 321428 190272 321434 190324
rect 328638 190272 328644 190324
rect 328696 190312 328702 190324
rect 329650 190312 329656 190324
rect 328696 190284 329656 190312
rect 328696 190272 328702 190284
rect 329650 190272 329656 190284
rect 329708 190272 329714 190324
rect 219802 190204 219808 190256
rect 219860 190244 219866 190256
rect 220630 190244 220636 190256
rect 219860 190216 220636 190244
rect 219860 190204 219866 190216
rect 220630 190204 220636 190216
rect 220688 190204 220694 190256
rect 332778 190204 332784 190256
rect 332836 190244 332842 190256
rect 333882 190244 333888 190256
rect 332836 190216 333888 190244
rect 332836 190204 332842 190216
rect 333882 190204 333888 190216
rect 333940 190204 333946 190256
rect 355042 190204 355048 190256
rect 355100 190244 355106 190256
rect 355870 190244 355876 190256
rect 355100 190216 355876 190244
rect 355100 190204 355106 190216
rect 355870 190204 355876 190216
rect 355928 190204 355934 190256
rect 443270 190204 443276 190256
rect 443328 190244 443334 190256
rect 444190 190244 444196 190256
rect 443328 190216 444196 190244
rect 443328 190204 443334 190216
rect 444190 190204 444196 190216
rect 444248 190204 444254 190256
rect 201586 190136 201592 190188
rect 201644 190176 201650 190188
rect 202690 190176 202696 190188
rect 201644 190148 202696 190176
rect 201644 190136 201650 190148
rect 202690 190136 202696 190148
rect 202748 190136 202754 190188
rect 281626 190136 281632 190188
rect 281684 190176 281690 190188
rect 282730 190176 282736 190188
rect 281684 190148 282736 190176
rect 281684 190136 281690 190148
rect 282730 190136 282736 190148
rect 282788 190136 282794 190188
rect 408586 190136 408592 190188
rect 408644 190176 408650 190188
rect 409690 190176 409696 190188
rect 408644 190148 409696 190176
rect 408644 190136 408650 190148
rect 409690 190136 409696 190148
rect 409748 190136 409754 190188
rect 416866 190136 416872 190188
rect 416924 190176 416930 190188
rect 417970 190176 417976 190188
rect 416924 190148 417976 190176
rect 416924 190136 416930 190148
rect 417970 190136 417976 190148
rect 418028 190136 418034 190188
rect 154666 190068 154672 190120
rect 154724 190108 154730 190120
rect 155770 190108 155776 190120
rect 154724 190080 155776 190108
rect 154724 190068 154730 190080
rect 155770 190068 155776 190080
rect 155828 190068 155834 190120
rect 244550 190068 244556 190120
rect 244608 190108 244614 190120
rect 245470 190108 245476 190120
rect 244608 190080 245476 190108
rect 244608 190068 244614 190080
rect 245470 190068 245476 190080
rect 245528 190068 245534 190120
rect 253566 190068 253572 190120
rect 253624 190108 253630 190120
rect 257338 190108 257344 190120
rect 253624 190080 257344 190108
rect 253624 190068 253630 190080
rect 257338 190068 257344 190080
rect 257396 190068 257402 190120
rect 316218 190068 316224 190120
rect 316276 190108 316282 190120
rect 317230 190108 317236 190120
rect 316276 190080 317236 190108
rect 316276 190068 316282 190080
rect 317230 190068 317236 190080
rect 317288 190068 317294 190120
rect 353386 190068 353392 190120
rect 353444 190108 353450 190120
rect 354490 190108 354496 190120
rect 353444 190080 354496 190108
rect 353444 190068 353450 190080
rect 354490 190068 354496 190080
rect 354548 190068 354554 190120
rect 379790 190068 379796 190120
rect 379848 190108 379854 190120
rect 380710 190108 380716 190120
rect 379848 190080 380716 190108
rect 379848 190068 379854 190080
rect 380710 190068 380716 190080
rect 380768 190068 380774 190120
rect 441614 190068 441620 190120
rect 441672 190108 441678 190120
rect 442810 190108 442816 190120
rect 441672 190080 442816 190108
rect 441672 190068 441678 190080
rect 442810 190068 442816 190080
rect 442868 190068 442874 190120
rect 361574 190000 361580 190052
rect 361632 190040 361638 190052
rect 362770 190040 362776 190052
rect 361632 190012 362776 190040
rect 361632 190000 361638 190012
rect 362770 190000 362776 190012
rect 362828 190000 362834 190052
rect 369854 190000 369860 190052
rect 369912 190040 369918 190052
rect 371050 190040 371056 190052
rect 369912 190012 371056 190040
rect 369912 190000 369918 190012
rect 371050 190000 371056 190012
rect 371108 190000 371114 190052
rect 433334 190000 433340 190052
rect 433392 190040 433398 190052
rect 434530 190040 434536 190052
rect 433392 190012 434536 190040
rect 433392 190000 433398 190012
rect 434530 190000 434536 190012
rect 434588 190000 434594 190052
rect 237926 189932 237932 189984
rect 237984 189972 237990 189984
rect 238662 189972 238668 189984
rect 237984 189944 238668 189972
rect 237984 189932 237990 189944
rect 238662 189932 238668 189944
rect 238720 189932 238726 189984
rect 269206 189932 269212 189984
rect 269264 189972 269270 189984
rect 270310 189972 270316 189984
rect 269264 189944 270316 189972
rect 269264 189932 269270 189944
rect 270310 189932 270316 189944
rect 270368 189932 270374 189984
rect 270862 189932 270868 189984
rect 270920 189972 270926 189984
rect 271966 189972 271972 189984
rect 270920 189944 271972 189972
rect 270920 189932 270926 189944
rect 271966 189932 271972 189944
rect 272024 189932 272030 189984
rect 340966 189932 340972 189984
rect 341024 189972 341030 189984
rect 342070 189972 342076 189984
rect 341024 189944 342076 189972
rect 341024 189932 341030 189944
rect 342070 189932 342076 189944
rect 342128 189932 342134 189984
rect 373166 189932 373172 189984
rect 373224 189972 373230 189984
rect 373902 189972 373908 189984
rect 373224 189944 373908 189972
rect 373224 189932 373230 189944
rect 373902 189932 373908 189944
rect 373960 189932 373966 189984
rect 421006 189932 421012 189984
rect 421064 189972 421070 189984
rect 422110 189972 422116 189984
rect 421064 189944 422116 189972
rect 421064 189932 421070 189944
rect 422110 189932 422116 189944
rect 422168 189932 422174 189984
rect 158714 189796 158720 189848
rect 158772 189836 158778 189848
rect 159910 189836 159916 189848
rect 158772 189808 159916 189836
rect 158772 189796 158778 189808
rect 159910 189796 159916 189808
rect 159968 189796 159974 189848
rect 176102 189796 176108 189848
rect 176160 189836 176166 189848
rect 184198 189836 184204 189848
rect 176160 189808 184204 189836
rect 176160 189796 176166 189808
rect 184198 189796 184204 189808
rect 184256 189796 184262 189848
rect 240410 189796 240416 189848
rect 240468 189836 240474 189848
rect 255958 189836 255964 189848
rect 240468 189808 255964 189836
rect 240468 189796 240474 189808
rect 255958 189796 255964 189808
rect 256016 189796 256022 189848
rect 257706 189796 257712 189848
rect 257764 189836 257770 189848
rect 301498 189836 301504 189848
rect 257764 189808 301504 189836
rect 257764 189796 257770 189808
rect 301498 189796 301504 189808
rect 301556 189796 301562 189848
rect 448238 189796 448244 189848
rect 448296 189836 448302 189848
rect 456058 189836 456064 189848
rect 448296 189808 456064 189836
rect 448296 189796 448302 189808
rect 456058 189796 456064 189808
rect 456116 189796 456122 189848
rect 180978 189728 180984 189780
rect 181036 189768 181042 189780
rect 192478 189768 192484 189780
rect 181036 189740 192484 189768
rect 181036 189728 181042 189740
rect 192478 189728 192484 189740
rect 192536 189728 192542 189780
rect 195882 189728 195888 189780
rect 195940 189768 195946 189780
rect 213178 189768 213184 189780
rect 195940 189740 213184 189768
rect 195940 189728 195946 189740
rect 213178 189728 213184 189740
rect 213236 189728 213242 189780
rect 223114 189728 223120 189780
rect 223172 189768 223178 189780
rect 242158 189768 242164 189780
rect 223172 189740 242164 189768
rect 223172 189728 223178 189740
rect 242158 189728 242164 189740
rect 242216 189728 242222 189780
rect 274174 189728 274180 189780
rect 274232 189768 274238 189780
rect 280798 189768 280804 189780
rect 274232 189740 280804 189768
rect 274232 189728 274238 189740
rect 280798 189728 280804 189740
rect 280856 189728 280862 189780
rect 294782 189728 294788 189780
rect 294840 189768 294846 189780
rect 352558 189768 352564 189780
rect 294840 189740 352564 189768
rect 294840 189728 294846 189740
rect 352558 189728 352564 189740
rect 352616 189728 352622 189780
rect 359182 189728 359188 189780
rect 359240 189768 359246 189780
rect 381538 189768 381544 189780
rect 359240 189740 381544 189768
rect 359240 189728 359246 189740
rect 381538 189728 381544 189740
rect 381596 189728 381602 189780
rect 383838 189728 383844 189780
rect 383896 189768 383902 189780
rect 485774 189768 485780 189780
rect 383896 189740 485780 189768
rect 383896 189728 383902 189740
rect 485774 189728 485780 189740
rect 485832 189728 485838 189780
rect 229646 189660 229652 189712
rect 229704 189700 229710 189712
rect 230382 189700 230388 189712
rect 229704 189672 230388 189700
rect 229704 189660 229710 189672
rect 230382 189660 230388 189672
rect 230440 189660 230446 189712
rect 309686 189660 309692 189712
rect 309744 189700 309750 189712
rect 310422 189700 310428 189712
rect 309744 189672 310428 189700
rect 309744 189660 309750 189672
rect 310422 189660 310428 189672
rect 310480 189660 310486 189712
rect 334434 189660 334440 189712
rect 334492 189700 334498 189712
rect 335262 189700 335268 189712
rect 334492 189672 335268 189700
rect 334492 189660 334498 189672
rect 335262 189660 335268 189672
rect 335320 189660 335326 189712
rect 364886 189660 364892 189712
rect 364944 189700 364950 189712
rect 365622 189700 365628 189712
rect 364944 189672 365628 189700
rect 364944 189660 364950 189672
rect 365622 189660 365628 189672
rect 365680 189660 365686 189712
rect 428366 189660 428372 189712
rect 428424 189700 428430 189712
rect 429102 189700 429108 189712
rect 428424 189672 429108 189700
rect 428424 189660 428430 189672
rect 429102 189660 429108 189672
rect 429160 189660 429166 189712
rect 234614 189524 234620 189576
rect 234672 189564 234678 189576
rect 235810 189564 235816 189576
rect 234672 189536 235816 189564
rect 234672 189524 234678 189536
rect 235810 189524 235816 189536
rect 235868 189524 235874 189576
rect 397914 189524 397920 189576
rect 397972 189564 397978 189576
rect 398742 189564 398748 189576
rect 397972 189536 398748 189564
rect 397972 189524 397978 189536
rect 398742 189524 398748 189536
rect 398800 189524 398806 189576
rect 449894 189524 449900 189576
rect 449952 189564 449958 189576
rect 451182 189564 451188 189576
rect 449952 189536 451188 189564
rect 449952 189524 449958 189536
rect 451182 189524 451188 189536
rect 451240 189524 451246 189576
rect 222286 189456 222292 189508
rect 222344 189496 222350 189508
rect 223482 189496 223488 189508
rect 222344 189468 223488 189496
rect 222344 189456 222350 189468
rect 223482 189456 223488 189468
rect 223540 189456 223546 189508
rect 250254 189456 250260 189508
rect 250312 189496 250318 189508
rect 251082 189496 251088 189508
rect 250312 189468 251088 189496
rect 250312 189456 250318 189468
rect 251082 189456 251088 189468
rect 251140 189456 251146 189508
rect 285766 189456 285772 189508
rect 285824 189496 285830 189508
rect 286962 189496 286968 189508
rect 285824 189468 286968 189496
rect 285824 189456 285830 189468
rect 286962 189456 286968 189468
rect 287020 189456 287026 189508
rect 322014 189456 322020 189508
rect 322072 189496 322078 189508
rect 322842 189496 322848 189508
rect 322072 189468 322848 189496
rect 322072 189456 322078 189468
rect 322842 189456 322848 189468
rect 322900 189456 322906 189508
rect 330294 189456 330300 189508
rect 330352 189496 330358 189508
rect 331122 189496 331128 189508
rect 330352 189468 331128 189496
rect 330352 189456 330358 189468
rect 331122 189456 331128 189468
rect 331180 189456 331186 189508
rect 387978 189456 387984 189508
rect 388036 189496 388042 189508
rect 389082 189496 389088 189508
rect 388036 189468 389088 189496
rect 388036 189456 388042 189468
rect 389082 189456 389088 189468
rect 389140 189456 389146 189508
rect 175274 189388 175280 189440
rect 175332 189428 175338 189440
rect 176562 189428 176568 189440
rect 175332 189400 176568 189428
rect 175332 189388 175338 189400
rect 176562 189388 176568 189400
rect 176620 189388 176626 189440
rect 182634 189388 182640 189440
rect 182692 189428 182698 189440
rect 183462 189428 183468 189440
rect 182692 189400 183468 189428
rect 182692 189388 182698 189400
rect 183462 189388 183468 189400
rect 183520 189388 183526 189440
rect 203242 189388 203248 189440
rect 203300 189428 203306 189440
rect 204162 189428 204168 189440
rect 203300 189400 204168 189428
rect 203300 189388 203306 189400
rect 204162 189388 204168 189400
rect 204220 189388 204226 189440
rect 275002 189388 275008 189440
rect 275060 189428 275066 189440
rect 275922 189428 275928 189440
rect 275060 189400 275928 189428
rect 275060 189388 275066 189400
rect 275922 189388 275928 189400
rect 275980 189388 275986 189440
rect 293954 189388 293960 189440
rect 294012 189428 294018 189440
rect 295242 189428 295248 189440
rect 294012 189400 295248 189428
rect 294012 189388 294018 189400
rect 295242 189388 295248 189400
rect 295300 189388 295306 189440
rect 317874 189388 317880 189440
rect 317932 189428 317938 189440
rect 318702 189428 318708 189440
rect 317932 189400 318708 189428
rect 317932 189388 317938 189400
rect 318702 189388 318708 189400
rect 318760 189388 318766 189440
rect 346762 189388 346768 189440
rect 346820 189428 346826 189440
rect 347682 189428 347688 189440
rect 346820 189400 347688 189428
rect 346820 189388 346826 189400
rect 347682 189388 347688 189400
rect 347740 189388 347746 189440
rect 410242 189388 410248 189440
rect 410300 189428 410306 189440
rect 411162 189428 411168 189440
rect 410300 189400 411168 189428
rect 410300 189388 410306 189400
rect 411162 189388 411168 189400
rect 411220 189388 411226 189440
rect 447410 189388 447416 189440
rect 447468 189428 447474 189440
rect 448422 189428 448428 189440
rect 447468 189400 448428 189428
rect 447468 189388 447474 189400
rect 448422 189388 448428 189400
rect 448480 189388 448486 189440
rect 156230 189320 156236 189372
rect 156288 189360 156294 189372
rect 157242 189360 157248 189372
rect 156288 189332 157248 189360
rect 156288 189320 156294 189332
rect 157242 189320 157248 189332
rect 157300 189320 157306 189372
rect 164510 189320 164516 189372
rect 164568 189360 164574 189372
rect 165522 189360 165528 189372
rect 164568 189332 165528 189360
rect 164568 189320 164574 189332
rect 165522 189320 165528 189332
rect 165580 189320 165586 189372
rect 172790 189320 172796 189372
rect 172848 189360 172854 189372
rect 173802 189360 173808 189372
rect 172848 189332 173808 189360
rect 172848 189320 172854 189332
rect 173802 189320 173808 189332
rect 173860 189320 173866 189372
rect 197538 189320 197544 189372
rect 197596 189360 197602 189372
rect 198642 189360 198648 189372
rect 197596 189332 198648 189360
rect 197596 189320 197602 189332
rect 198642 189320 198648 189332
rect 198700 189320 198706 189372
rect 214006 189320 214012 189372
rect 214064 189360 214070 189372
rect 215202 189360 215208 189372
rect 214064 189332 215208 189360
rect 214064 189320 214070 189332
rect 215202 189320 215208 189332
rect 215260 189320 215266 189372
rect 236270 189320 236276 189372
rect 236328 189360 236334 189372
rect 237282 189360 237288 189372
rect 236328 189332 237288 189360
rect 236328 189320 236334 189332
rect 237282 189320 237288 189332
rect 237340 189320 237346 189372
rect 261018 189320 261024 189372
rect 261076 189360 261082 189372
rect 262122 189360 262128 189372
rect 261076 189332 262128 189360
rect 261076 189320 261082 189332
rect 262122 189320 262128 189332
rect 262180 189320 262186 189372
rect 277486 189320 277492 189372
rect 277544 189360 277550 189372
rect 278682 189360 278688 189372
rect 277544 189332 278688 189360
rect 277544 189320 277550 189332
rect 278682 189320 278688 189332
rect 278740 189320 278746 189372
rect 299750 189320 299756 189372
rect 299808 189360 299814 189372
rect 300762 189360 300768 189372
rect 299808 189332 300768 189360
rect 299808 189320 299814 189332
rect 300762 189320 300768 189332
rect 300820 189320 300826 189372
rect 349246 189320 349252 189372
rect 349304 189360 349310 189372
rect 350442 189360 350448 189372
rect 349304 189332 350448 189360
rect 349304 189320 349310 189332
rect 350442 189320 350448 189332
rect 350500 189320 350506 189372
rect 371510 189320 371516 189372
rect 371568 189360 371574 189372
rect 372522 189360 372528 189372
rect 371568 189332 372528 189360
rect 371568 189320 371574 189332
rect 372522 189320 372528 189332
rect 372580 189320 372586 189372
rect 412726 189320 412732 189372
rect 412784 189360 412790 189372
rect 413922 189360 413928 189372
rect 412784 189332 413928 189360
rect 412784 189320 412790 189332
rect 413922 189320 413928 189332
rect 413980 189320 413986 189372
rect 434990 189320 434996 189372
rect 435048 189360 435054 189372
rect 436002 189360 436008 189372
rect 435048 189332 436008 189360
rect 435048 189320 435054 189332
rect 436002 189320 436008 189332
rect 436060 189320 436066 189372
rect 185118 189252 185124 189304
rect 185176 189292 185182 189304
rect 186222 189292 186228 189304
rect 185176 189264 186228 189292
rect 185176 189252 185182 189264
rect 186222 189252 186228 189264
rect 186280 189252 186286 189304
rect 193398 189252 193404 189304
rect 193456 189292 193462 189304
rect 194502 189292 194508 189304
rect 193456 189264 194508 189292
rect 193456 189252 193462 189264
rect 194502 189252 194508 189264
rect 194560 189252 194566 189304
rect 205726 189252 205732 189304
rect 205784 189292 205790 189304
rect 206922 189292 206928 189304
rect 205784 189264 206928 189292
rect 205784 189252 205790 189264
rect 206922 189252 206928 189264
rect 206980 189252 206986 189304
rect 209866 189252 209872 189304
rect 209924 189292 209930 189304
rect 211062 189292 211068 189304
rect 209924 189264 211068 189292
rect 209924 189252 209930 189264
rect 211062 189252 211068 189264
rect 211120 189252 211126 189304
rect 223850 189252 223856 189304
rect 223908 189292 223914 189304
rect 224862 189292 224868 189304
rect 223908 189264 224868 189292
rect 223908 189252 223914 189264
rect 224862 189252 224868 189264
rect 224920 189252 224926 189304
rect 230474 189252 230480 189304
rect 230532 189292 230538 189304
rect 231762 189292 231768 189304
rect 230532 189264 231768 189292
rect 230532 189252 230538 189264
rect 231762 189252 231768 189264
rect 231820 189252 231826 189304
rect 238754 189252 238760 189304
rect 238812 189292 238818 189304
rect 240042 189292 240048 189304
rect 238812 189264 240048 189292
rect 238812 189252 238818 189264
rect 240042 189252 240048 189264
rect 240100 189252 240106 189304
rect 248598 189252 248604 189304
rect 248656 189292 248662 189304
rect 249702 189292 249708 189304
rect 248656 189264 249708 189292
rect 248656 189252 248662 189264
rect 249702 189252 249708 189264
rect 249760 189252 249766 189304
rect 265158 189252 265164 189304
rect 265216 189292 265222 189304
rect 266262 189292 266268 189304
rect 265216 189264 266268 189292
rect 265216 189252 265222 189264
rect 266262 189252 266268 189264
rect 266320 189252 266326 189304
rect 302234 189252 302240 189304
rect 302292 189292 302298 189304
rect 303522 189292 303528 189304
rect 302292 189264 303528 189292
rect 302292 189252 302298 189264
rect 303522 189252 303528 189264
rect 303580 189252 303586 189304
rect 306374 189252 306380 189304
rect 306432 189292 306438 189304
rect 307662 189292 307668 189304
rect 306432 189264 307668 189292
rect 306432 189252 306438 189264
rect 307662 189252 307668 189264
rect 307720 189252 307726 189304
rect 310514 189252 310520 189304
rect 310572 189292 310578 189304
rect 311802 189292 311808 189304
rect 310572 189264 311808 189292
rect 310572 189252 310578 189264
rect 311802 189252 311808 189264
rect 311860 189252 311866 189304
rect 312170 189252 312176 189304
rect 312228 189292 312234 189304
rect 313182 189292 313188 189304
rect 312228 189264 313188 189292
rect 312228 189252 312234 189264
rect 313182 189252 313188 189264
rect 313240 189252 313246 189304
rect 336918 189252 336924 189304
rect 336976 189292 336982 189304
rect 338022 189292 338028 189304
rect 336976 189264 338028 189292
rect 336976 189252 336982 189264
rect 338022 189252 338028 189264
rect 338080 189252 338086 189304
rect 345106 189252 345112 189304
rect 345164 189292 345170 189304
rect 346302 189292 346308 189304
rect 345164 189264 346308 189292
rect 345164 189252 345170 189264
rect 346302 189252 346308 189264
rect 346360 189252 346366 189304
rect 365714 189252 365720 189304
rect 365772 189292 365778 189304
rect 367002 189292 367008 189304
rect 365772 189264 367008 189292
rect 365772 189252 365778 189264
rect 367002 189252 367008 189264
rect 367060 189252 367066 189304
rect 373994 189252 374000 189304
rect 374052 189292 374058 189304
rect 375282 189292 375288 189304
rect 374052 189264 375288 189292
rect 374052 189252 374058 189264
rect 375282 189252 375288 189264
rect 375340 189252 375346 189304
rect 375650 189252 375656 189304
rect 375708 189292 375714 189304
rect 376662 189292 376668 189304
rect 375708 189264 376668 189292
rect 375708 189252 375714 189264
rect 376662 189252 376668 189264
rect 376720 189252 376726 189304
rect 378134 189252 378140 189304
rect 378192 189292 378198 189304
rect 379422 189292 379428 189304
rect 378192 189264 379428 189292
rect 378192 189252 378198 189264
rect 379422 189252 379428 189264
rect 379480 189252 379486 189304
rect 400398 189252 400404 189304
rect 400456 189292 400462 189304
rect 401502 189292 401508 189304
rect 400456 189264 401508 189292
rect 400456 189252 400462 189264
rect 401502 189252 401508 189264
rect 401560 189252 401566 189304
rect 437474 189252 437480 189304
rect 437532 189292 437538 189304
rect 438762 189292 438768 189304
rect 437532 189264 438768 189292
rect 437532 189252 437538 189264
rect 438762 189252 438768 189264
rect 438820 189252 438826 189304
rect 160370 189116 160376 189168
rect 160428 189156 160434 189168
rect 161382 189156 161388 189168
rect 160428 189128 161388 189156
rect 160428 189116 160434 189128
rect 161382 189116 161388 189128
rect 161440 189116 161446 189168
rect 213546 189116 213552 189168
rect 213604 189156 213610 189168
rect 221274 189156 221280 189168
rect 213604 189128 221280 189156
rect 213604 189116 213610 189128
rect 221274 189116 221280 189128
rect 221332 189116 221338 189168
rect 283282 189116 283288 189168
rect 283340 189156 283346 189168
rect 284110 189156 284116 189168
rect 283340 189128 284116 189156
rect 283340 189116 283346 189128
rect 284110 189116 284116 189128
rect 284168 189116 284174 189168
rect 307202 189116 307208 189168
rect 307260 189156 307266 189168
rect 309778 189156 309784 189168
rect 307260 189128 309784 189156
rect 307260 189116 307266 189128
rect 309778 189116 309784 189128
rect 309836 189116 309842 189168
rect 378962 189116 378968 189168
rect 379020 189156 379026 189168
rect 384298 189156 384304 189168
rect 379020 189128 384304 189156
rect 379020 189116 379026 189128
rect 384298 189116 384304 189128
rect 384356 189116 384362 189168
rect 418522 189116 418528 189168
rect 418580 189156 418586 189168
rect 419350 189156 419356 189168
rect 418580 189128 419356 189156
rect 418580 189116 418586 189128
rect 419350 189116 419356 189128
rect 419408 189116 419414 189168
rect 445754 189116 445760 189168
rect 445812 189156 445818 189168
rect 451918 189156 451924 189168
rect 445812 189128 451924 189156
rect 445812 189116 445818 189128
rect 451918 189116 451924 189128
rect 451976 189116 451982 189168
rect 157886 189048 157892 189100
rect 157944 189088 157950 189100
rect 158622 189088 158628 189100
rect 157944 189060 158628 189088
rect 157944 189048 157950 189060
rect 158622 189048 158628 189060
rect 158680 189048 158686 189100
rect 162854 189048 162860 189100
rect 162912 189088 162918 189100
rect 164142 189088 164148 189100
rect 162912 189060 164148 189088
rect 162912 189048 162918 189060
rect 164142 189048 164148 189060
rect 164200 189048 164206 189100
rect 166166 189048 166172 189100
rect 166224 189088 166230 189100
rect 166902 189088 166908 189100
rect 166224 189060 166908 189088
rect 166224 189048 166230 189060
rect 166902 189048 166908 189060
rect 166960 189048 166966 189100
rect 166994 189048 167000 189100
rect 167052 189088 167058 189100
rect 168190 189088 168196 189100
rect 167052 189060 168196 189088
rect 167052 189048 167058 189060
rect 168190 189048 168196 189060
rect 168248 189048 168254 189100
rect 171134 189048 171140 189100
rect 171192 189088 171198 189100
rect 172330 189088 172336 189100
rect 171192 189060 172336 189088
rect 171192 189048 171198 189060
rect 172330 189048 172336 189060
rect 172388 189048 172394 189100
rect 174446 189048 174452 189100
rect 174504 189088 174510 189100
rect 175182 189088 175188 189100
rect 174504 189060 175188 189088
rect 174504 189048 174510 189060
rect 175182 189048 175188 189060
rect 175240 189048 175246 189100
rect 176930 189048 176936 189100
rect 176988 189088 176994 189100
rect 177850 189088 177856 189100
rect 176988 189060 177856 189088
rect 176988 189048 176994 189060
rect 177850 189048 177856 189060
rect 177908 189048 177914 189100
rect 178494 189048 178500 189100
rect 178552 189088 178558 189100
rect 179230 189088 179236 189100
rect 178552 189060 179236 189088
rect 178552 189048 178558 189060
rect 179230 189048 179236 189060
rect 179288 189048 179294 189100
rect 186774 189048 186780 189100
rect 186832 189088 186838 189100
rect 187510 189088 187516 189100
rect 186832 189060 187516 189088
rect 186832 189048 186838 189060
rect 187510 189048 187516 189060
rect 187568 189048 187574 189100
rect 189258 189048 189264 189100
rect 189316 189088 189322 189100
rect 190270 189088 190276 189100
rect 189316 189060 190276 189088
rect 189316 189048 189322 189060
rect 190270 189048 190276 189060
rect 190328 189048 190334 189100
rect 190914 189048 190920 189100
rect 190972 189088 190978 189100
rect 191742 189088 191748 189100
rect 190972 189060 191748 189088
rect 190972 189048 190978 189060
rect 191742 189048 191748 189060
rect 191800 189048 191806 189100
rect 195054 189048 195060 189100
rect 195112 189088 195118 189100
rect 195882 189088 195888 189100
rect 195112 189060 195888 189088
rect 195112 189048 195118 189060
rect 195882 189048 195888 189060
rect 195940 189048 195946 189100
rect 199194 189048 199200 189100
rect 199252 189088 199258 189100
rect 200758 189088 200764 189100
rect 199252 189060 200764 189088
rect 199252 189048 199258 189060
rect 200758 189048 200764 189060
rect 200816 189048 200822 189100
rect 207382 189048 207388 189100
rect 207440 189088 207446 189100
rect 208302 189088 208308 189100
rect 207440 189060 208308 189088
rect 207440 189048 207446 189060
rect 208302 189048 208308 189060
rect 208360 189048 208366 189100
rect 211522 189048 211528 189100
rect 211580 189088 211586 189100
rect 212350 189088 212356 189100
rect 211580 189060 212356 189088
rect 211580 189048 211586 189060
rect 212350 189048 212356 189060
rect 212408 189048 212414 189100
rect 215662 189048 215668 189100
rect 215720 189088 215726 189100
rect 216582 189088 216588 189100
rect 215720 189060 216588 189088
rect 215720 189048 215726 189060
rect 216582 189048 216588 189060
rect 216640 189048 216646 189100
rect 218146 189048 218152 189100
rect 218204 189088 218210 189100
rect 219342 189088 219348 189100
rect 218204 189060 219348 189088
rect 218204 189048 218210 189060
rect 219342 189048 219348 189060
rect 219400 189048 219406 189100
rect 221458 189048 221464 189100
rect 221516 189088 221522 189100
rect 222838 189088 222844 189100
rect 221516 189060 222844 189088
rect 221516 189048 221522 189060
rect 222838 189048 222844 189060
rect 222896 189048 222902 189100
rect 226334 189048 226340 189100
rect 226392 189088 226398 189100
rect 227622 189088 227628 189100
rect 226392 189060 227628 189088
rect 226392 189048 226398 189060
rect 227622 189048 227628 189060
rect 227680 189048 227686 189100
rect 227990 189048 227996 189100
rect 228048 189088 228054 189100
rect 229002 189088 229008 189100
rect 228048 189060 229008 189088
rect 228048 189048 228054 189060
rect 229002 189048 229008 189060
rect 229060 189048 229066 189100
rect 232130 189048 232136 189100
rect 232188 189088 232194 189100
rect 233050 189088 233056 189100
rect 232188 189060 233056 189088
rect 232188 189048 232194 189060
rect 233050 189048 233056 189060
rect 233108 189048 233114 189100
rect 242894 189048 242900 189100
rect 242952 189088 242958 189100
rect 244182 189088 244188 189100
rect 242952 189060 244188 189088
rect 242952 189048 242958 189060
rect 244182 189048 244188 189060
rect 244240 189048 244246 189100
rect 246114 189048 246120 189100
rect 246172 189088 246178 189100
rect 246942 189088 246948 189100
rect 246172 189060 246948 189088
rect 246172 189048 246178 189060
rect 246942 189048 246948 189060
rect 247000 189048 247006 189100
rect 256878 189048 256884 189100
rect 256936 189088 256942 189100
rect 257982 189088 257988 189100
rect 256936 189060 257988 189088
rect 256936 189048 256942 189060
rect 257982 189048 257988 189060
rect 258040 189048 258046 189100
rect 258534 189048 258540 189100
rect 258592 189088 258598 189100
rect 259270 189088 259276 189100
rect 258592 189060 259276 189088
rect 258592 189048 258598 189060
rect 259270 189048 259276 189060
rect 259328 189048 259334 189100
rect 262674 189048 262680 189100
rect 262732 189088 262738 189100
rect 263502 189088 263508 189100
rect 262732 189060 263508 189088
rect 262732 189048 262738 189060
rect 263502 189048 263508 189060
rect 263560 189048 263566 189100
rect 266814 189048 266820 189100
rect 266872 189088 266878 189100
rect 267550 189088 267556 189100
rect 266872 189060 267556 189088
rect 266872 189048 266878 189060
rect 267550 189048 267556 189060
rect 267608 189048 267614 189100
rect 273346 189048 273352 189100
rect 273404 189088 273410 189100
rect 274542 189088 274548 189100
rect 273404 189060 274548 189088
rect 273404 189048 273410 189060
rect 274542 189048 274548 189060
rect 274600 189048 274606 189100
rect 279142 189048 279148 189100
rect 279200 189088 279206 189100
rect 279970 189088 279976 189100
rect 279200 189060 279976 189088
rect 279200 189048 279206 189060
rect 279970 189048 279976 189060
rect 280028 189048 280034 189100
rect 287422 189048 287428 189100
rect 287480 189088 287486 189100
rect 288342 189088 288348 189100
rect 287480 189060 288348 189088
rect 287480 189048 287486 189060
rect 288342 189048 288348 189060
rect 288400 189048 288406 189100
rect 289906 189048 289912 189100
rect 289964 189088 289970 189100
rect 291102 189088 291108 189100
rect 289964 189060 291108 189088
rect 289964 189048 289970 189060
rect 291102 189048 291108 189060
rect 291160 189048 291166 189100
rect 291562 189048 291568 189100
rect 291620 189088 291626 189100
rect 292390 189088 292396 189100
rect 291620 189060 292396 189088
rect 291620 189048 291626 189060
rect 292390 189048 292396 189060
rect 292448 189048 292454 189100
rect 293126 189048 293132 189100
rect 293184 189088 293190 189100
rect 293862 189088 293868 189100
rect 293184 189060 293868 189088
rect 293184 189048 293190 189060
rect 293862 189048 293868 189060
rect 293920 189048 293926 189100
rect 298094 189048 298100 189100
rect 298152 189088 298158 189100
rect 299382 189088 299388 189100
rect 298152 189060 299388 189088
rect 298152 189048 298158 189060
rect 299382 189048 299388 189060
rect 299440 189048 299446 189100
rect 301406 189048 301412 189100
rect 301464 189088 301470 189100
rect 302142 189088 302148 189100
rect 301464 189060 302148 189088
rect 301464 189048 301470 189060
rect 302142 189048 302148 189060
rect 302200 189048 302206 189100
rect 308030 189048 308036 189100
rect 308088 189088 308094 189100
rect 308950 189088 308956 189100
rect 308088 189060 308956 189088
rect 308088 189048 308094 189060
rect 308950 189048 308956 189060
rect 309008 189048 309014 189100
rect 324498 189048 324504 189100
rect 324556 189088 324562 189100
rect 327718 189088 327724 189100
rect 324556 189060 327724 189088
rect 324556 189048 324562 189060
rect 327718 189048 327724 189060
rect 327776 189048 327782 189100
rect 338482 189048 338488 189100
rect 338540 189088 338546 189100
rect 339310 189088 339316 189100
rect 338540 189060 339316 189088
rect 338540 189048 338546 189060
rect 339310 189048 339316 189060
rect 339368 189048 339374 189100
rect 342622 189048 342628 189100
rect 342680 189088 342686 189100
rect 344278 189088 344284 189100
rect 342680 189060 344284 189088
rect 342680 189048 342686 189060
rect 344278 189048 344284 189060
rect 344336 189048 344342 189100
rect 350902 189048 350908 189100
rect 350960 189088 350966 189100
rect 351730 189088 351736 189100
rect 350960 189060 351736 189088
rect 350960 189048 350966 189060
rect 351730 189048 351736 189060
rect 351788 189048 351794 189100
rect 357526 189048 357532 189100
rect 357584 189088 357590 189100
rect 358630 189088 358636 189100
rect 357584 189060 358636 189088
rect 357584 189048 357590 189060
rect 358630 189048 358636 189060
rect 358688 189048 358694 189100
rect 363230 189048 363236 189100
rect 363288 189088 363294 189100
rect 364242 189088 364248 189100
rect 363288 189060 364248 189088
rect 363288 189048 363294 189060
rect 364242 189048 364248 189060
rect 364300 189048 364306 189100
rect 381446 189048 381452 189100
rect 381504 189088 381510 189100
rect 382182 189088 382188 189100
rect 381504 189060 382188 189088
rect 381504 189048 381510 189060
rect 382182 189048 382188 189060
rect 382240 189048 382246 189100
rect 382274 189048 382280 189100
rect 382332 189088 382338 189100
rect 383470 189088 383476 189100
rect 382332 189060 383476 189088
rect 382332 189048 382338 189060
rect 383470 189048 383476 189060
rect 383528 189048 383534 189100
rect 385494 189048 385500 189100
rect 385552 189088 385558 189100
rect 386230 189088 386236 189100
rect 385552 189060 386236 189088
rect 385552 189048 385558 189060
rect 386230 189048 386236 189060
rect 386288 189048 386294 189100
rect 389634 189048 389640 189100
rect 389692 189088 389698 189100
rect 390462 189088 390468 189100
rect 389692 189060 390468 189088
rect 389692 189048 389698 189060
rect 390462 189048 390468 189060
rect 390520 189048 390526 189100
rect 392118 189048 392124 189100
rect 392176 189088 392182 189100
rect 393130 189088 393136 189100
rect 392176 189060 393136 189088
rect 392176 189048 392182 189060
rect 393130 189048 393136 189060
rect 393188 189048 393194 189100
rect 402054 189048 402060 189100
rect 402112 189088 402118 189100
rect 402882 189088 402888 189100
rect 402112 189060 402888 189088
rect 402112 189048 402118 189060
rect 402882 189048 402888 189060
rect 402940 189048 402946 189100
rect 404538 189048 404544 189100
rect 404596 189088 404602 189100
rect 405550 189088 405556 189100
rect 404596 189060 405556 189088
rect 404596 189048 404602 189060
rect 405550 189048 405556 189060
rect 405608 189048 405614 189100
rect 406102 189048 406108 189100
rect 406160 189088 406166 189100
rect 406930 189088 406936 189100
rect 406160 189060 406936 189088
rect 406160 189048 406166 189060
rect 406930 189048 406936 189060
rect 406988 189048 406994 189100
rect 414382 189048 414388 189100
rect 414440 189088 414446 189100
rect 416038 189088 416044 189100
rect 414440 189060 416044 189088
rect 414440 189048 414446 189060
rect 416038 189048 416044 189060
rect 416096 189048 416102 189100
rect 422662 189048 422668 189100
rect 422720 189088 422726 189100
rect 423582 189088 423588 189100
rect 422720 189060 423588 189088
rect 422720 189048 422726 189060
rect 423582 189048 423588 189060
rect 423640 189048 423646 189100
rect 425146 189048 425152 189100
rect 425204 189088 425210 189100
rect 426342 189088 426348 189100
rect 425204 189060 426348 189088
rect 425204 189048 425210 189060
rect 426342 189048 426348 189060
rect 426400 189048 426406 189100
rect 426802 189048 426808 189100
rect 426860 189088 426866 189100
rect 427630 189088 427636 189100
rect 426860 189060 427636 189088
rect 426860 189048 426866 189060
rect 427630 189048 427636 189060
rect 427688 189048 427694 189100
rect 429194 189048 429200 189100
rect 429252 189088 429258 189100
rect 430390 189088 430396 189100
rect 429252 189060 430396 189088
rect 429252 189048 429258 189060
rect 430390 189048 430396 189060
rect 430448 189048 430454 189100
rect 430850 189048 430856 189100
rect 430908 189088 430914 189100
rect 431770 189088 431776 189100
rect 430908 189060 431776 189088
rect 430908 189048 430914 189060
rect 431770 189048 431776 189060
rect 431828 189048 431834 189100
rect 436646 189048 436652 189100
rect 436704 189088 436710 189100
rect 437382 189088 437388 189100
rect 436704 189060 437388 189088
rect 436704 189048 436710 189060
rect 437382 189048 437388 189060
rect 437440 189048 437446 189100
rect 444926 189048 444932 189100
rect 444984 189088 444990 189100
rect 445662 189088 445668 189100
rect 444984 189060 445668 189088
rect 444984 189048 444990 189060
rect 445662 189048 445668 189060
rect 445720 189048 445726 189100
rect 235442 188300 235448 188352
rect 235500 188340 235506 188352
rect 271874 188340 271880 188352
rect 235500 188312 271880 188340
rect 235500 188300 235506 188312
rect 271874 188300 271880 188312
rect 271932 188300 271938 188352
rect 271966 188300 271972 188352
rect 272024 188340 272030 188352
rect 322934 188340 322940 188352
rect 272024 188312 322940 188340
rect 272024 188300 272030 188312
rect 322934 188300 322940 188312
rect 322992 188300 322998 188352
rect 386322 188300 386328 188352
rect 386380 188340 386386 188352
rect 489914 188340 489920 188352
rect 386380 188312 489920 188340
rect 386380 188300 386386 188312
rect 489914 188300 489920 188312
rect 489972 188300 489978 188352
rect 252738 186940 252744 186992
rect 252796 186980 252802 186992
rect 296714 186980 296720 186992
rect 252796 186952 296720 186980
rect 252796 186940 252802 186952
rect 296714 186940 296720 186952
rect 296772 186940 296778 186992
rect 388806 186940 388812 186992
rect 388864 186980 388870 186992
rect 494054 186980 494060 186992
rect 388864 186952 494060 186980
rect 388864 186940 388870 186952
rect 494054 186940 494060 186952
rect 494112 186940 494118 186992
rect 138014 185580 138020 185632
rect 138072 185620 138078 185632
rect 138566 185620 138572 185632
rect 138072 185592 138572 185620
rect 138072 185580 138078 185592
rect 138566 185580 138572 185592
rect 138624 185580 138630 185632
rect 139394 185580 139400 185632
rect 139452 185620 139458 185632
rect 140222 185620 140228 185632
rect 139452 185592 140228 185620
rect 139452 185580 139458 185592
rect 140222 185580 140228 185592
rect 140280 185580 140286 185632
rect 143534 185580 143540 185632
rect 143592 185620 143598 185632
rect 144454 185620 144460 185632
rect 143592 185592 144460 185620
rect 143592 185580 143598 185592
rect 144454 185580 144460 185592
rect 144512 185580 144518 185632
rect 146294 185580 146300 185632
rect 146352 185620 146358 185632
rect 146846 185620 146852 185632
rect 146352 185592 146852 185620
rect 146352 185580 146358 185592
rect 146846 185580 146852 185592
rect 146904 185580 146910 185632
rect 147674 185580 147680 185632
rect 147732 185620 147738 185632
rect 148502 185620 148508 185632
rect 147732 185592 148508 185620
rect 147732 185580 147738 185592
rect 148502 185580 148508 185592
rect 148560 185580 148566 185632
rect 393774 185580 393780 185632
rect 393832 185620 393838 185632
rect 500954 185620 500960 185632
rect 393832 185592 500960 185620
rect 393832 185580 393838 185592
rect 500954 185580 500960 185592
rect 501012 185580 501018 185632
rect 396258 184152 396264 184204
rect 396316 184192 396322 184204
rect 503714 184192 503720 184204
rect 396316 184164 503720 184192
rect 396316 184152 396322 184164
rect 503714 184152 503720 184164
rect 503772 184152 503778 184204
rect 398650 182792 398656 182844
rect 398708 182832 398714 182844
rect 507854 182832 507860 182844
rect 398708 182804 507860 182832
rect 398708 182792 398714 182804
rect 507854 182792 507860 182804
rect 507912 182792 507918 182844
rect 453666 182112 453672 182164
rect 453724 182152 453730 182164
rect 580166 182152 580172 182164
rect 453724 182124 580172 182152
rect 453724 182112 453730 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 133874 181432 133880 181484
rect 133932 181472 133938 181484
rect 134518 181472 134524 181484
rect 133932 181444 134524 181472
rect 133932 181432 133938 181444
rect 134518 181432 134524 181444
rect 134576 181432 134582 181484
rect 367370 181432 367376 181484
rect 367428 181472 367434 181484
rect 462314 181472 462320 181484
rect 367428 181444 462320 181472
rect 367428 181432 367434 181444
rect 462314 181432 462320 181444
rect 462372 181432 462378 181484
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 17218 180792 17224 180804
rect 3292 180764 17224 180792
rect 3292 180752 3298 180764
rect 17218 180752 17224 180764
rect 17276 180752 17282 180804
rect 401410 180072 401416 180124
rect 401468 180112 401474 180124
rect 511994 180112 512000 180124
rect 401468 180084 512000 180112
rect 401468 180072 401474 180084
rect 511994 180072 512000 180084
rect 512052 180072 512058 180124
rect 275830 178644 275836 178696
rect 275888 178684 275894 178696
rect 331214 178684 331220 178696
rect 275888 178656 331220 178684
rect 275888 178644 275894 178656
rect 331214 178644 331220 178656
rect 331272 178644 331278 178696
rect 406930 178644 406936 178696
rect 406988 178684 406994 178696
rect 518894 178684 518900 178696
rect 406988 178656 518900 178684
rect 406988 178644 406994 178656
rect 518894 178644 518900 178656
rect 518952 178644 518958 178696
rect 259270 177284 259276 177336
rect 259328 177324 259334 177336
rect 304994 177324 305000 177336
rect 259328 177296 305000 177324
rect 259328 177284 259334 177296
rect 304994 177284 305000 177296
rect 305052 177284 305058 177336
rect 314470 177284 314476 177336
rect 314528 177324 314534 177336
rect 385034 177324 385040 177336
rect 314528 177296 385040 177324
rect 314528 177284 314534 177296
rect 385034 177284 385040 177296
rect 385092 177284 385098 177336
rect 409690 177284 409696 177336
rect 409748 177324 409754 177336
rect 521654 177324 521660 177336
rect 409748 177296 521660 177324
rect 409748 177284 409754 177296
rect 521654 177284 521660 177296
rect 521712 177284 521718 177336
rect 411070 175924 411076 175976
rect 411128 175964 411134 175976
rect 525794 175964 525800 175976
rect 411128 175936 525800 175964
rect 411128 175924 411134 175936
rect 525794 175924 525800 175936
rect 525852 175924 525858 175976
rect 413830 174496 413836 174548
rect 413888 174536 413894 174548
rect 528554 174536 528560 174548
rect 413888 174508 528560 174536
rect 413888 174496 413894 174508
rect 528554 174496 528560 174508
rect 528612 174496 528618 174548
rect 135346 173884 135352 173936
rect 135404 173924 135410 173936
rect 135622 173924 135628 173936
rect 135404 173896 135628 173924
rect 135404 173884 135410 173896
rect 135622 173884 135628 173896
rect 135680 173884 135686 173936
rect 419350 173136 419356 173188
rect 419408 173176 419414 173188
rect 536834 173176 536840 173188
rect 419408 173148 536840 173176
rect 419408 173136 419414 173148
rect 536834 173136 536840 173148
rect 536892 173136 536898 173188
rect 422110 171776 422116 171828
rect 422168 171816 422174 171828
rect 539594 171816 539600 171828
rect 422168 171788 539600 171816
rect 422168 171776 422174 171788
rect 539594 171776 539600 171788
rect 539652 171776 539658 171828
rect 453574 171028 453580 171080
rect 453632 171068 453638 171080
rect 580166 171068 580172 171080
rect 453632 171040 580172 171068
rect 453632 171028 453638 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 423490 168988 423496 169040
rect 423548 169028 423554 169040
rect 543734 169028 543740 169040
rect 423548 169000 543740 169028
rect 423548 168988 423554 169000
rect 543734 168988 543740 169000
rect 543792 168988 543798 169040
rect 426250 167628 426256 167680
rect 426308 167668 426314 167680
rect 546494 167668 546500 167680
rect 426308 167640 546500 167668
rect 426308 167628 426314 167640
rect 546494 167628 546500 167640
rect 546552 167628 546558 167680
rect 431770 166268 431776 166320
rect 431828 166308 431834 166320
rect 554774 166308 554780 166320
rect 431828 166280 554780 166308
rect 431828 166268 431834 166280
rect 554774 166268 554780 166280
rect 554832 166268 554838 166320
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 126238 165560 126244 165572
rect 3568 165532 126244 165560
rect 3568 165520 3574 165532
rect 126238 165520 126244 165532
rect 126296 165520 126302 165572
rect 434530 164840 434536 164892
rect 434588 164880 434594 164892
rect 557534 164880 557540 164892
rect 434588 164852 557540 164880
rect 434588 164840 434594 164852
rect 557534 164840 557540 164852
rect 557592 164840 557598 164892
rect 135346 164160 135352 164212
rect 135404 164200 135410 164212
rect 135530 164200 135536 164212
rect 135404 164172 135536 164200
rect 135404 164160 135410 164172
rect 135530 164160 135536 164172
rect 135588 164160 135594 164212
rect 435910 163480 435916 163532
rect 435968 163520 435974 163532
rect 561674 163520 561680 163532
rect 435968 163492 561680 163520
rect 435968 163480 435974 163492
rect 561674 163480 561680 163492
rect 561732 163480 561738 163532
rect 438670 162120 438676 162172
rect 438728 162160 438734 162172
rect 564434 162160 564440 162172
rect 438728 162132 564440 162160
rect 438728 162120 438734 162132
rect 564434 162120 564440 162132
rect 564492 162120 564498 162172
rect 444190 160692 444196 160744
rect 444248 160732 444254 160744
rect 571334 160732 571340 160744
rect 444248 160704 571340 160732
rect 444248 160692 444254 160704
rect 571334 160692 571340 160704
rect 571392 160692 571398 160744
rect 364150 159332 364156 159384
rect 364208 159372 364214 159384
rect 458174 159372 458180 159384
rect 364208 159344 458180 159372
rect 364208 159332 364214 159344
rect 458174 159332 458180 159344
rect 458232 159332 458238 159384
rect 471238 158652 471244 158704
rect 471296 158692 471302 158704
rect 579798 158692 579804 158704
rect 471296 158664 579804 158692
rect 471296 158652 471302 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 366910 157972 366916 158024
rect 366968 158012 366974 158024
rect 460934 158012 460940 158024
rect 366968 157984 460940 158012
rect 366968 157972 366974 157984
rect 460934 157972 460940 157984
rect 460992 157972 460998 158024
rect 376570 156612 376576 156664
rect 376628 156652 376634 156664
rect 476114 156652 476120 156664
rect 376628 156624 476120 156652
rect 376628 156612 376634 156624
rect 476114 156612 476120 156624
rect 476172 156612 476178 156664
rect 383470 155184 383476 155236
rect 383528 155224 383534 155236
rect 484394 155224 484400 155236
rect 383528 155196 484400 155224
rect 383528 155184 383534 155196
rect 484394 155184 484400 155196
rect 484452 155184 484458 155236
rect 384942 153824 384948 153876
rect 385000 153864 385006 153876
rect 487154 153864 487160 153876
rect 385000 153836 487160 153864
rect 385000 153824 385006 153836
rect 487154 153824 487160 153836
rect 487212 153824 487218 153876
rect 393130 152464 393136 152516
rect 393188 152504 393194 152516
rect 498194 152504 498200 152516
rect 393188 152476 498200 152504
rect 393188 152464 393194 152476
rect 498194 152464 498200 152476
rect 498252 152464 498258 152516
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 129274 151756 129280 151768
rect 3200 151728 129280 151756
rect 3200 151716 3206 151728
rect 129274 151716 129280 151728
rect 129332 151716 129338 151768
rect 397362 151036 397368 151088
rect 397420 151076 397426 151088
rect 505094 151076 505100 151088
rect 397420 151048 505100 151076
rect 397420 151036 397426 151048
rect 505094 151036 505100 151048
rect 505152 151036 505158 151088
rect 405550 149676 405556 149728
rect 405608 149716 405614 149728
rect 516134 149716 516140 149728
rect 405608 149688 516140 149716
rect 405608 149676 405614 149688
rect 516134 149676 516140 149688
rect 516192 149676 516198 149728
rect 416038 148316 416044 148368
rect 416096 148356 416102 148368
rect 529934 148356 529940 148368
rect 416096 148328 529940 148356
rect 416096 148316 416102 148328
rect 529934 148316 529940 148328
rect 529992 148316 529998 148368
rect 417970 146888 417976 146940
rect 418028 146928 418034 146940
rect 534074 146928 534080 146940
rect 418028 146900 534080 146928
rect 418028 146888 418034 146900
rect 534074 146888 534080 146900
rect 534132 146888 534138 146940
rect 427630 145528 427636 145580
rect 427688 145568 427694 145580
rect 547874 145568 547880 145580
rect 427688 145540 547880 145568
rect 427688 145528 427694 145540
rect 547874 145528 547880 145540
rect 547932 145528 547938 145580
rect 430390 144168 430396 144220
rect 430448 144208 430454 144220
rect 552014 144208 552020 144220
rect 430448 144180 552020 144208
rect 430448 144168 430454 144180
rect 552014 144168 552020 144180
rect 552072 144168 552078 144220
rect 440050 142808 440056 142860
rect 440108 142848 440114 142860
rect 565814 142848 565820 142860
rect 440108 142820 565820 142848
rect 440108 142808 440114 142820
rect 565814 142808 565820 142820
rect 565872 142808 565878 142860
rect 442810 141380 442816 141432
rect 442868 141420 442874 141432
rect 569954 141420 569960 141432
rect 442868 141392 569960 141420
rect 442868 141380 442874 141392
rect 569954 141380 569960 141392
rect 570012 141380 570018 141432
rect 371050 140020 371056 140072
rect 371108 140060 371114 140072
rect 466454 140060 466460 140072
rect 371108 140032 466460 140060
rect 371108 140020 371114 140032
rect 466454 140020 466460 140032
rect 466512 140020 466518 140072
rect 375190 138660 375196 138712
rect 375248 138700 375254 138712
rect 473354 138700 473360 138712
rect 375248 138672 473360 138700
rect 375248 138660 375254 138672
rect 473354 138660 473360 138672
rect 473412 138660 473418 138712
rect 380710 137232 380716 137284
rect 380768 137272 380774 137284
rect 480254 137272 480260 137284
rect 380768 137244 480260 137272
rect 380768 137232 380774 137244
rect 480254 137232 480260 137244
rect 480312 137232 480318 137284
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 13078 136592 13084 136604
rect 3292 136564 13084 136592
rect 3292 136552 3298 136564
rect 13078 136552 13084 136564
rect 13136 136552 13142 136604
rect 390370 135872 390376 135924
rect 390428 135912 390434 135924
rect 495434 135912 495440 135924
rect 390428 135884 495440 135912
rect 390428 135872 390434 135884
rect 495434 135872 495440 135884
rect 495492 135872 495498 135924
rect 479518 135192 479524 135244
rect 479576 135232 479582 135244
rect 580166 135232 580172 135244
rect 479576 135204 580172 135232
rect 479576 135192 479582 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 313090 134512 313096 134564
rect 313148 134552 313154 134564
rect 383654 134552 383660 134564
rect 313148 134524 383660 134552
rect 313148 134512 313154 134524
rect 383654 134512 383660 134524
rect 383712 134512 383718 134564
rect 384298 134512 384304 134564
rect 384356 134552 384362 134564
rect 478874 134552 478880 134564
rect 384356 134524 478880 134552
rect 384356 134512 384362 134524
rect 478874 134512 478880 134524
rect 478932 134512 478938 134564
rect 402790 133152 402796 133204
rect 402848 133192 402854 133204
rect 513374 133192 513380 133204
rect 402848 133164 513380 133192
rect 402848 133152 402854 133164
rect 513374 133152 513380 133164
rect 513432 133152 513438 133204
rect 415302 131724 415308 131776
rect 415360 131764 415366 131776
rect 531314 131764 531320 131776
rect 415360 131736 531320 131764
rect 415360 131724 415366 131736
rect 531314 131724 531320 131736
rect 531372 131724 531378 131776
rect 433242 130364 433248 130416
rect 433300 130404 433306 130416
rect 556154 130404 556160 130416
rect 433300 130376 556160 130404
rect 433300 130364 433306 130376
rect 556154 130364 556160 130376
rect 556212 130364 556218 130416
rect 453482 124108 453488 124160
rect 453540 124148 453546 124160
rect 580166 124148 580172 124160
rect 453540 124120 580172 124148
rect 453540 124108 453546 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 14458 122788 14464 122800
rect 3476 122760 14464 122788
rect 3476 122748 3482 122760
rect 14458 122748 14464 122760
rect 14516 122748 14522 122800
rect 311710 117920 311716 117972
rect 311768 117960 311774 117972
rect 382274 117960 382280 117972
rect 311768 117932 382280 117960
rect 311768 117920 311774 117932
rect 382274 117920 382280 117932
rect 382332 117920 382338 117972
rect 307662 113772 307668 113824
rect 307720 113812 307726 113824
rect 373994 113812 374000 113824
rect 307720 113784 374000 113812
rect 307720 113772 307726 113784
rect 373994 113772 374000 113784
rect 374052 113772 374058 113824
rect 469858 111732 469864 111784
rect 469916 111772 469922 111784
rect 579798 111772 579804 111784
rect 469916 111744 579804 111772
rect 469916 111732 469922 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 372430 111052 372436 111104
rect 372488 111092 372494 111104
rect 469214 111092 469220 111104
rect 372488 111064 469220 111092
rect 372488 111052 372494 111064
rect 469214 111052 469220 111064
rect 469272 111052 469278 111104
rect 331030 109692 331036 109744
rect 331088 109732 331094 109744
rect 409874 109732 409880 109744
rect 331088 109704 409880 109732
rect 331088 109692 331094 109704
rect 409874 109692 409880 109704
rect 409932 109692 409938 109744
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 129182 108984 129188 108996
rect 3292 108956 129188 108984
rect 3292 108944 3298 108956
rect 129182 108944 129188 108956
rect 129240 108944 129246 108996
rect 321370 108264 321376 108316
rect 321428 108304 321434 108316
rect 394694 108304 394700 108316
rect 321428 108276 394700 108304
rect 321428 108264 321434 108276
rect 394694 108264 394700 108276
rect 394752 108264 394758 108316
rect 395982 108264 395988 108316
rect 396040 108304 396046 108316
rect 502334 108304 502340 108316
rect 396040 108276 502340 108304
rect 396040 108264 396046 108276
rect 502334 108264 502340 108276
rect 502392 108264 502398 108316
rect 354490 105544 354496 105596
rect 354548 105584 354554 105596
rect 442994 105584 443000 105596
rect 354548 105556 443000 105584
rect 354548 105544 354554 105556
rect 442994 105544 443000 105556
rect 443052 105544 443058 105596
rect 326890 104116 326896 104168
rect 326948 104156 326954 104168
rect 402974 104156 402980 104168
rect 326948 104128 402980 104156
rect 326948 104116 326954 104128
rect 402974 104116 402980 104128
rect 403032 104116 403038 104168
rect 351730 102756 351736 102808
rect 351788 102796 351794 102808
rect 438854 102796 438860 102808
rect 351788 102768 438860 102796
rect 351788 102756 351794 102768
rect 438854 102756 438860 102768
rect 438912 102756 438918 102808
rect 339310 101396 339316 101448
rect 339368 101436 339374 101448
rect 420914 101436 420920 101448
rect 339368 101408 420920 101436
rect 339368 101396 339374 101408
rect 420914 101396 420920 101408
rect 420972 101396 420978 101448
rect 346210 99968 346216 100020
rect 346268 100008 346274 100020
rect 431954 100008 431960 100020
rect 346268 99980 431960 100008
rect 346268 99968 346274 99980
rect 431954 99968 431960 99980
rect 432012 99968 432018 100020
rect 343542 98608 343548 98660
rect 343600 98648 343606 98660
rect 427814 98648 427820 98660
rect 343600 98620 427820 98648
rect 343600 98608 343606 98620
rect 427814 98608 427820 98620
rect 427872 98608 427878 98660
rect 342070 97248 342076 97300
rect 342128 97288 342134 97300
rect 425054 97288 425060 97300
rect 342128 97260 425060 97288
rect 342128 97248 342134 97260
rect 425054 97248 425060 97260
rect 425112 97248 425118 97300
rect 336642 95888 336648 95940
rect 336700 95928 336706 95940
rect 416774 95928 416780 95940
rect 336700 95900 416780 95928
rect 336700 95888 336706 95900
rect 416774 95888 416780 95900
rect 416832 95888 416838 95940
rect 333790 94460 333796 94512
rect 333848 94500 333854 94512
rect 414014 94500 414020 94512
rect 333848 94472 414020 94500
rect 333848 94460 333854 94472
rect 414014 94460 414020 94472
rect 414072 94460 414078 94512
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 19978 93820 19984 93832
rect 3476 93792 19984 93820
rect 3476 93780 3482 93792
rect 19978 93780 19984 93792
rect 20036 93780 20042 93832
rect 329650 93100 329656 93152
rect 329708 93140 329714 93152
rect 407114 93140 407120 93152
rect 329708 93112 407120 93140
rect 329708 93100 329714 93112
rect 407114 93100 407120 93112
rect 407172 93100 407178 93152
rect 324222 91740 324228 91792
rect 324280 91780 324286 91792
rect 400214 91780 400220 91792
rect 324280 91752 400220 91780
rect 324280 91740 324286 91752
rect 400214 91740 400220 91752
rect 400272 91740 400278 91792
rect 321462 90312 321468 90364
rect 321520 90352 321526 90364
rect 396074 90352 396080 90364
rect 321520 90324 396080 90352
rect 321520 90312 321526 90324
rect 396074 90312 396080 90324
rect 396132 90312 396138 90364
rect 318610 88952 318616 89004
rect 318668 88992 318674 89004
rect 391934 88992 391940 89004
rect 318668 88964 391940 88992
rect 318668 88952 318674 88964
rect 391934 88952 391940 88964
rect 391992 88952 391998 89004
rect 472618 88272 472624 88324
rect 472676 88312 472682 88324
rect 580166 88312 580172 88324
rect 472676 88284 580172 88312
rect 472676 88272 472682 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 375282 87592 375288 87644
rect 375340 87632 375346 87644
rect 471974 87632 471980 87644
rect 375340 87604 471980 87632
rect 375340 87592 375346 87604
rect 471974 87592 471980 87604
rect 472032 87592 472038 87644
rect 135349 86955 135407 86961
rect 135349 86921 135361 86955
rect 135395 86952 135407 86955
rect 135438 86952 135444 86964
rect 135395 86924 135444 86952
rect 135395 86921 135407 86924
rect 135349 86915 135407 86921
rect 135438 86912 135444 86924
rect 135496 86912 135502 86964
rect 317230 86232 317236 86284
rect 317288 86272 317294 86284
rect 389174 86272 389180 86284
rect 317288 86244 389180 86272
rect 317288 86232 317294 86244
rect 389174 86232 389180 86244
rect 389232 86232 389238 86284
rect 438762 86232 438768 86284
rect 438820 86272 438826 86284
rect 563054 86272 563060 86284
rect 438820 86244 563060 86272
rect 438820 86232 438826 86244
rect 563054 86232 563060 86244
rect 563112 86232 563118 86284
rect 304810 84804 304816 84856
rect 304868 84844 304874 84856
rect 371234 84844 371240 84856
rect 304868 84816 371240 84844
rect 304868 84804 304874 84816
rect 371234 84804 371240 84816
rect 371292 84804 371298 84856
rect 302142 83444 302148 83496
rect 302200 83484 302206 83496
rect 367094 83484 367100 83496
rect 302200 83456 367100 83484
rect 302200 83444 302206 83456
rect 367094 83444 367100 83456
rect 367152 83444 367158 83496
rect 430482 83444 430488 83496
rect 430540 83484 430546 83496
rect 553394 83484 553400 83496
rect 430540 83456 553400 83484
rect 430540 83444 430546 83456
rect 553394 83444 553400 83456
rect 553452 83444 553458 83496
rect 299290 82084 299296 82136
rect 299348 82124 299354 82136
rect 364334 82124 364340 82136
rect 299348 82096 364340 82124
rect 299348 82084 299354 82096
rect 364334 82084 364340 82096
rect 364392 82084 364398 82136
rect 398742 82084 398748 82136
rect 398800 82124 398806 82136
rect 506474 82124 506480 82136
rect 398800 82096 506480 82124
rect 398800 82084 398806 82096
rect 506474 82084 506480 82096
rect 506532 82084 506538 82136
rect 295242 80656 295248 80708
rect 295300 80696 295306 80708
rect 356054 80696 356060 80708
rect 295300 80668 356060 80696
rect 295300 80656 295306 80668
rect 356054 80656 356060 80668
rect 356112 80656 356118 80708
rect 365622 80656 365628 80708
rect 365680 80696 365686 80708
rect 459646 80696 459652 80708
rect 365680 80668 459652 80696
rect 365680 80656 365686 80668
rect 459646 80656 459652 80668
rect 459704 80656 459710 80708
rect 3510 79432 3516 79484
rect 3568 79472 3574 79484
rect 8938 79472 8944 79484
rect 3568 79444 8944 79472
rect 3568 79432 3574 79444
rect 8938 79432 8944 79444
rect 8996 79432 9002 79484
rect 292390 79296 292396 79348
rect 292448 79336 292454 79348
rect 353294 79336 353300 79348
rect 292448 79308 353300 79336
rect 292448 79296 292454 79308
rect 353294 79296 353300 79308
rect 353352 79296 353358 79348
rect 401502 79296 401508 79348
rect 401560 79336 401566 79348
rect 510614 79336 510620 79348
rect 401560 79308 510620 79336
rect 401560 79296 401566 79308
rect 510614 79296 510620 79308
rect 510672 79296 510678 79348
rect 289722 77936 289728 77988
rect 289780 77976 289786 77988
rect 349154 77976 349160 77988
rect 289780 77948 349160 77976
rect 289780 77936 289786 77948
rect 349154 77936 349160 77948
rect 349212 77936 349218 77988
rect 418062 77936 418068 77988
rect 418120 77976 418126 77988
rect 535454 77976 535460 77988
rect 418120 77948 535460 77976
rect 418120 77936 418126 77948
rect 535454 77936 535460 77948
rect 535512 77936 535518 77988
rect 135346 77296 135352 77308
rect 135307 77268 135352 77296
rect 135346 77256 135352 77268
rect 135404 77256 135410 77308
rect 453390 77188 453396 77240
rect 453448 77228 453454 77240
rect 580166 77228 580172 77240
rect 453448 77200 580172 77228
rect 453448 77188 453454 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 135346 77160 135352 77172
rect 135307 77132 135352 77160
rect 135346 77120 135352 77132
rect 135404 77120 135410 77172
rect 286870 76508 286876 76560
rect 286928 76548 286934 76560
rect 346394 76548 346400 76560
rect 286928 76520 346400 76548
rect 286928 76508 286934 76520
rect 346394 76508 346400 76520
rect 346452 76508 346458 76560
rect 349062 76508 349068 76560
rect 349120 76548 349126 76560
rect 434714 76548 434720 76560
rect 349120 76520 434720 76548
rect 349120 76508 349126 76520
rect 434714 76508 434720 76520
rect 434772 76508 434778 76560
rect 335170 75148 335176 75200
rect 335228 75188 335234 75200
rect 416866 75188 416872 75200
rect 335228 75160 416872 75188
rect 335228 75148 335234 75160
rect 416866 75148 416872 75160
rect 416924 75148 416930 75200
rect 423582 75148 423588 75200
rect 423640 75188 423646 75200
rect 542354 75188 542360 75200
rect 423640 75160 542360 75188
rect 423640 75148 423646 75160
rect 542354 75148 542360 75160
rect 542412 75148 542418 75200
rect 282730 73788 282736 73840
rect 282788 73828 282794 73840
rect 339494 73828 339500 73840
rect 282788 73800 339500 73828
rect 282788 73788 282794 73800
rect 339494 73788 339500 73800
rect 339552 73788 339558 73840
rect 355870 73788 355876 73840
rect 355928 73828 355934 73840
rect 444374 73828 444380 73840
rect 355928 73800 444380 73828
rect 355928 73788 355934 73800
rect 444374 73788 444380 73800
rect 444432 73788 444438 73840
rect 445662 73788 445668 73840
rect 445720 73828 445726 73840
rect 573358 73828 573364 73840
rect 445720 73800 573364 73828
rect 445720 73788 445726 73800
rect 573358 73788 573364 73800
rect 573416 73788 573422 73840
rect 333882 72428 333888 72480
rect 333940 72468 333946 72480
rect 412634 72468 412640 72480
rect 333940 72440 412640 72468
rect 333940 72428 333946 72440
rect 412634 72428 412640 72440
rect 412692 72428 412698 72480
rect 420822 72428 420828 72480
rect 420880 72468 420886 72480
rect 538214 72468 538220 72480
rect 420880 72440 538220 72468
rect 420880 72428 420886 72440
rect 538214 72428 538220 72440
rect 538272 72428 538278 72480
rect 279970 71000 279976 71052
rect 280028 71040 280034 71052
rect 335354 71040 335360 71052
rect 280028 71012 335360 71040
rect 280028 71000 280034 71012
rect 335354 71000 335360 71012
rect 335412 71000 335418 71052
rect 347590 71000 347596 71052
rect 347648 71040 347654 71052
rect 433334 71040 433340 71052
rect 347648 71012 433340 71040
rect 347648 71000 347654 71012
rect 433334 71000 433340 71012
rect 433392 71000 433398 71052
rect 436002 71000 436008 71052
rect 436060 71040 436066 71052
rect 560294 71040 560300 71052
rect 436060 71012 560300 71040
rect 436060 71000 436066 71012
rect 560294 71000 560300 71012
rect 560352 71000 560358 71052
rect 135349 70295 135407 70301
rect 135349 70261 135361 70295
rect 135395 70292 135407 70295
rect 135438 70292 135444 70304
rect 135395 70264 135444 70292
rect 135395 70261 135407 70264
rect 135349 70255 135407 70261
rect 135438 70252 135444 70264
rect 135496 70252 135502 70304
rect 331122 69640 331128 69692
rect 331180 69680 331186 69692
rect 408494 69680 408500 69692
rect 331180 69652 408500 69680
rect 331180 69640 331186 69652
rect 408494 69640 408500 69652
rect 408552 69640 408558 69692
rect 411162 69640 411168 69692
rect 411220 69680 411226 69692
rect 524414 69680 524420 69692
rect 411220 69652 524420 69680
rect 411220 69640 411226 69652
rect 524414 69640 524420 69652
rect 524472 69640 524478 69692
rect 271782 68280 271788 68332
rect 271840 68320 271846 68332
rect 324314 68320 324320 68332
rect 271840 68292 324320 68320
rect 271840 68280 271846 68292
rect 324314 68280 324320 68292
rect 324372 68280 324378 68332
rect 328362 68280 328368 68332
rect 328420 68320 328426 68332
rect 405734 68320 405740 68332
rect 328420 68292 405740 68320
rect 328420 68280 328426 68292
rect 405734 68280 405740 68292
rect 405792 68280 405798 68332
rect 408402 68280 408408 68332
rect 408460 68320 408466 68332
rect 520274 68320 520280 68332
rect 408460 68292 520280 68320
rect 408460 68280 408466 68292
rect 520274 68280 520280 68292
rect 520332 68280 520338 68332
rect 270310 66852 270316 66904
rect 270368 66892 270374 66904
rect 321554 66892 321560 66904
rect 270368 66864 321560 66892
rect 270368 66852 270374 66864
rect 321554 66852 321560 66864
rect 321612 66852 321618 66904
rect 325602 66852 325608 66904
rect 325660 66892 325666 66904
rect 401594 66892 401600 66904
rect 325660 66864 401600 66892
rect 325660 66852 325666 66864
rect 401594 66852 401600 66864
rect 401652 66852 401658 66904
rect 413922 66852 413928 66904
rect 413980 66892 413986 66904
rect 528646 66892 528652 66904
rect 413980 66864 528652 66892
rect 413980 66852 413986 66864
rect 528646 66852 528652 66864
rect 528704 66852 528710 66904
rect 267550 65492 267556 65544
rect 267608 65532 267614 65544
rect 317414 65532 317420 65544
rect 267608 65504 317420 65532
rect 267608 65492 267614 65504
rect 317414 65492 317420 65504
rect 317472 65492 317478 65544
rect 322750 65492 322756 65544
rect 322808 65532 322814 65544
rect 398834 65532 398840 65544
rect 322808 65504 398840 65532
rect 322808 65492 322814 65504
rect 398834 65492 398840 65504
rect 398892 65492 398898 65544
rect 405642 65492 405648 65544
rect 405700 65532 405706 65544
rect 517514 65532 517520 65544
rect 405700 65504 517520 65532
rect 405700 65492 405706 65504
rect 517514 65492 517520 65504
rect 517572 65492 517578 65544
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 129090 64852 129096 64864
rect 3384 64824 129096 64852
rect 3384 64812 3390 64824
rect 129090 64812 129096 64824
rect 129148 64812 129154 64864
rect 454678 64812 454684 64864
rect 454736 64852 454742 64864
rect 579798 64852 579804 64864
rect 454736 64824 579804 64852
rect 454736 64812 454742 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 262030 64132 262036 64184
rect 262088 64172 262094 64184
rect 310514 64172 310520 64184
rect 262088 64144 310520 64172
rect 262088 64132 262094 64144
rect 310514 64132 310520 64144
rect 310572 64132 310578 64184
rect 362770 64132 362776 64184
rect 362828 64172 362834 64184
rect 454034 64172 454040 64184
rect 362828 64144 454040 64172
rect 362828 64132 362834 64144
rect 454034 64132 454040 64144
rect 454092 64132 454098 64184
rect 259362 62772 259368 62824
rect 259420 62812 259426 62824
rect 306374 62812 306380 62824
rect 259420 62784 306380 62812
rect 259420 62772 259426 62784
rect 306374 62772 306380 62784
rect 306432 62772 306438 62824
rect 318702 62772 318708 62824
rect 318760 62812 318766 62824
rect 390554 62812 390560 62824
rect 318760 62784 390560 62812
rect 318760 62772 318766 62784
rect 390554 62772 390560 62784
rect 390612 62772 390618 62824
rect 393222 62772 393228 62824
rect 393280 62812 393286 62824
rect 499574 62812 499580 62824
rect 393280 62784 499580 62812
rect 393280 62772 393286 62784
rect 499574 62772 499580 62784
rect 499632 62772 499638 62824
rect 306282 61344 306288 61396
rect 306340 61384 306346 61396
rect 374086 61384 374092 61396
rect 306340 61356 374092 61384
rect 306340 61344 306346 61356
rect 374086 61344 374092 61356
rect 374144 61344 374150 61396
rect 389082 61344 389088 61396
rect 389140 61384 389146 61396
rect 492674 61384 492680 61396
rect 389140 61356 492680 61384
rect 389140 61344 389146 61356
rect 492674 61344 492680 61356
rect 492732 61344 492738 61396
rect 135438 60664 135444 60716
rect 135496 60704 135502 60716
rect 135622 60704 135628 60716
rect 135496 60676 135628 60704
rect 135496 60664 135502 60676
rect 135622 60664 135628 60676
rect 135680 60664 135686 60716
rect 257982 59984 257988 60036
rect 258040 60024 258046 60036
rect 303614 60024 303620 60036
rect 258040 59996 303620 60024
rect 258040 59984 258046 59996
rect 303614 59984 303620 59996
rect 303672 59984 303678 60036
rect 308950 59984 308956 60036
rect 309008 60024 309014 60036
rect 376754 60024 376760 60036
rect 309008 59996 376760 60024
rect 309008 59984 309014 59996
rect 376754 59984 376760 59996
rect 376812 59984 376818 60036
rect 386230 59984 386236 60036
rect 386288 60024 386294 60036
rect 488534 60024 488540 60036
rect 386288 59996 488540 60024
rect 386288 59984 386294 59996
rect 488534 59984 488540 59996
rect 488592 59984 488598 60036
rect 255130 58624 255136 58676
rect 255188 58664 255194 58676
rect 299474 58664 299480 58676
rect 255188 58636 299480 58664
rect 255188 58624 255194 58636
rect 299474 58624 299480 58636
rect 299532 58624 299538 58676
rect 303430 58624 303436 58676
rect 303488 58664 303494 58676
rect 369854 58664 369860 58676
rect 303488 58636 369860 58664
rect 303488 58624 303494 58636
rect 369854 58624 369860 58636
rect 369912 58624 369918 58676
rect 383562 58624 383568 58676
rect 383620 58664 383626 58676
rect 485866 58664 485872 58676
rect 383620 58636 485872 58664
rect 383620 58624 383626 58636
rect 485866 58624 485872 58636
rect 485924 58624 485930 58676
rect 135533 57919 135591 57925
rect 135533 57885 135545 57919
rect 135579 57916 135591 57919
rect 135622 57916 135628 57928
rect 135579 57888 135628 57916
rect 135579 57885 135591 57888
rect 135533 57879 135591 57885
rect 135622 57876 135628 57888
rect 135680 57876 135686 57928
rect 249610 57196 249616 57248
rect 249668 57236 249674 57248
rect 292574 57236 292580 57248
rect 249668 57208 292580 57236
rect 249668 57196 249674 57208
rect 292574 57196 292580 57208
rect 292632 57196 292638 57248
rect 300670 57196 300676 57248
rect 300728 57236 300734 57248
rect 365714 57236 365720 57248
rect 300728 57208 365720 57236
rect 300728 57196 300734 57208
rect 365714 57196 365720 57208
rect 365772 57196 365778 57248
rect 378042 57196 378048 57248
rect 378100 57236 378106 57248
rect 477586 57236 477592 57248
rect 378100 57208 477592 57236
rect 378100 57196 378106 57208
rect 477586 57196 477592 57208
rect 477644 57196 477650 57248
rect 299382 55904 299388 55956
rect 299440 55944 299446 55956
rect 362954 55944 362960 55956
rect 299440 55916 362960 55944
rect 299440 55904 299446 55916
rect 362954 55904 362960 55916
rect 363012 55904 363018 55956
rect 362862 55836 362868 55888
rect 362920 55876 362926 55888
rect 455414 55876 455420 55888
rect 362920 55848 455420 55876
rect 362920 55836 362926 55848
rect 455414 55836 455420 55848
rect 455472 55836 455478 55888
rect 246850 54476 246856 54528
rect 246908 54516 246914 54528
rect 288434 54516 288440 54528
rect 246908 54488 288440 54516
rect 246908 54476 246914 54488
rect 288434 54476 288440 54488
rect 288492 54476 288498 54528
rect 296530 54476 296536 54528
rect 296588 54516 296594 54528
rect 358814 54516 358820 54528
rect 296588 54488 358820 54516
rect 296588 54476 296594 54488
rect 358814 54476 358820 54488
rect 358872 54476 358878 54528
rect 360102 54476 360108 54528
rect 360160 54516 360166 54528
rect 451274 54516 451280 54528
rect 360160 54488 451280 54516
rect 360160 54476 360166 54488
rect 451274 54476 451280 54488
rect 451332 54476 451338 54528
rect 245470 53048 245476 53100
rect 245528 53088 245534 53100
rect 285674 53088 285680 53100
rect 245528 53060 285680 53088
rect 245528 53048 245534 53060
rect 285674 53048 285680 53060
rect 285732 53048 285738 53100
rect 293862 53048 293868 53100
rect 293920 53088 293926 53100
rect 356146 53088 356152 53100
rect 293920 53060 356152 53088
rect 293920 53048 293926 53060
rect 356146 53048 356152 53060
rect 356204 53048 356210 53100
rect 358630 53048 358636 53100
rect 358688 53088 358694 53100
rect 448514 53088 448520 53100
rect 358688 53060 448520 53088
rect 358688 53048 358694 53060
rect 448514 53048 448520 53060
rect 448572 53048 448578 53100
rect 242802 51688 242808 51740
rect 242860 51728 242866 51740
rect 281534 51728 281540 51740
rect 242860 51700 281540 51728
rect 242860 51688 242866 51700
rect 281534 51688 281540 51700
rect 281592 51688 281598 51740
rect 291010 51688 291016 51740
rect 291068 51728 291074 51740
rect 351914 51728 351920 51740
rect 291068 51700 351920 51728
rect 291068 51688 291074 51700
rect 351914 51688 351920 51700
rect 351972 51688 351978 51740
rect 353202 51688 353208 51740
rect 353260 51728 353266 51740
rect 441614 51728 441620 51740
rect 353260 51700 441620 51728
rect 353260 51688 353266 51700
rect 441614 51688 441620 51700
rect 441672 51688 441678 51740
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 15838 51048 15844 51060
rect 3476 51020 15844 51048
rect 3476 51008 3482 51020
rect 15838 51008 15844 51020
rect 15896 51008 15902 51060
rect 239950 50328 239956 50380
rect 240008 50368 240014 50380
rect 278774 50368 278780 50380
rect 240008 50340 278780 50368
rect 240008 50328 240014 50340
rect 278774 50328 278780 50340
rect 278832 50328 278838 50380
rect 288250 50328 288256 50380
rect 288308 50368 288314 50380
rect 347774 50368 347780 50380
rect 288308 50340 347780 50368
rect 288308 50328 288314 50340
rect 347774 50328 347780 50340
rect 347832 50328 347838 50380
rect 350350 50328 350356 50380
rect 350408 50368 350414 50380
rect 437474 50368 437480 50380
rect 350408 50340 437480 50368
rect 350408 50328 350414 50340
rect 437474 50328 437480 50340
rect 437532 50328 437538 50380
rect 442902 50328 442908 50380
rect 442960 50368 442966 50380
rect 571426 50368 571432 50380
rect 442960 50340 571432 50368
rect 442960 50328 442966 50340
rect 571426 50328 571432 50340
rect 571484 50328 571490 50380
rect 233050 48968 233056 49020
rect 233108 49008 233114 49020
rect 267734 49008 267740 49020
rect 233108 48980 267740 49008
rect 233108 48968 233114 48980
rect 267734 48968 267740 48980
rect 267792 48968 267798 49020
rect 284110 48968 284116 49020
rect 284168 49008 284174 49020
rect 340874 49008 340880 49020
rect 284168 48980 340880 49008
rect 284168 48968 284174 48980
rect 340874 48968 340880 48980
rect 340932 48968 340938 49020
rect 344278 48968 344284 49020
rect 344336 49008 344342 49020
rect 426434 49008 426440 49020
rect 344336 48980 426440 49008
rect 344336 48968 344342 48980
rect 426434 48968 426440 48980
rect 426492 48968 426498 49020
rect 427722 48968 427728 49020
rect 427780 49008 427786 49020
rect 549254 49008 549260 49020
rect 427780 48980 549260 49008
rect 427780 48968 427786 48980
rect 549254 48968 549260 48980
rect 549312 48968 549318 49020
rect 135530 48328 135536 48340
rect 135491 48300 135536 48328
rect 135530 48288 135536 48300
rect 135588 48288 135594 48340
rect 237190 47540 237196 47592
rect 237248 47580 237254 47592
rect 274634 47580 274640 47592
rect 237248 47552 274640 47580
rect 237248 47540 237254 47552
rect 274634 47540 274640 47552
rect 274692 47540 274698 47592
rect 281442 47540 281448 47592
rect 281500 47580 281506 47592
rect 338114 47580 338120 47592
rect 281500 47552 338120 47580
rect 281500 47540 281506 47552
rect 338114 47540 338120 47552
rect 338172 47540 338178 47592
rect 340782 47540 340788 47592
rect 340840 47580 340846 47592
rect 423674 47580 423680 47592
rect 340840 47552 423680 47580
rect 340840 47540 340846 47552
rect 423674 47540 423680 47552
rect 423732 47540 423738 47592
rect 447042 47540 447048 47592
rect 447100 47580 447106 47592
rect 574738 47580 574744 47592
rect 447100 47552 574744 47580
rect 447100 47540 447106 47552
rect 574738 47540 574744 47552
rect 574796 47540 574802 47592
rect 244090 46180 244096 46232
rect 244148 46220 244154 46232
rect 284294 46220 284300 46232
rect 244148 46192 284300 46220
rect 244148 46180 244154 46192
rect 284294 46180 284300 46192
rect 284352 46180 284358 46232
rect 286962 46180 286968 46232
rect 287020 46220 287026 46232
rect 345014 46220 345020 46232
rect 287020 46192 345020 46220
rect 287020 46180 287026 46192
rect 345014 46180 345020 46192
rect 345072 46180 345078 46232
rect 346302 46180 346308 46232
rect 346360 46220 346366 46232
rect 430574 46220 430580 46232
rect 346360 46192 430580 46220
rect 346360 46180 346366 46192
rect 430574 46180 430580 46192
rect 430632 46180 430638 46232
rect 440142 46180 440148 46232
rect 440200 46220 440206 46232
rect 567194 46220 567200 46232
rect 440200 46192 567200 46220
rect 440200 46180 440206 46192
rect 567194 46180 567200 46192
rect 567252 46180 567258 46232
rect 235810 44820 235816 44872
rect 235868 44860 235874 44872
rect 270494 44860 270500 44872
rect 235868 44832 270500 44860
rect 235868 44820 235874 44832
rect 270494 44820 270500 44832
rect 270552 44820 270558 44872
rect 278590 44820 278596 44872
rect 278648 44860 278654 44872
rect 333974 44860 333980 44872
rect 278648 44832 333980 44860
rect 278648 44820 278654 44832
rect 333974 44820 333980 44832
rect 334032 44820 334038 44872
rect 337930 44820 337936 44872
rect 337988 44860 337994 44872
rect 419534 44860 419540 44872
rect 337988 44832 419540 44860
rect 337988 44820 337994 44832
rect 419534 44820 419540 44832
rect 419592 44820 419598 44872
rect 426342 44820 426348 44872
rect 426400 44860 426406 44872
rect 546586 44860 546592 44872
rect 426400 44832 546592 44860
rect 426400 44820 426406 44832
rect 546586 44820 546592 44832
rect 546644 44820 546650 44872
rect 230382 43392 230388 43444
rect 230440 43432 230446 43444
rect 263594 43432 263600 43444
rect 230440 43404 263600 43432
rect 230440 43392 230446 43404
rect 263594 43392 263600 43404
rect 263652 43392 263658 43444
rect 274542 43392 274548 43444
rect 274600 43432 274606 43444
rect 327074 43432 327080 43444
rect 274600 43404 327080 43432
rect 274600 43392 274606 43404
rect 327074 43392 327080 43404
rect 327132 43392 327138 43444
rect 347682 43392 347688 43444
rect 347740 43432 347746 43444
rect 433426 43432 433432 43444
rect 347740 43404 433432 43432
rect 347740 43392 347746 43404
rect 433426 43392 433432 43404
rect 433484 43392 433490 43444
rect 434622 43392 434628 43444
rect 434680 43432 434686 43444
rect 558914 43432 558920 43444
rect 434680 43404 558920 43432
rect 434680 43392 434686 43404
rect 558914 43392 558920 43404
rect 558972 43392 558978 43444
rect 266170 42100 266176 42152
rect 266228 42140 266234 42152
rect 316034 42140 316040 42152
rect 266228 42112 316040 42140
rect 266228 42100 266234 42112
rect 316034 42100 316040 42112
rect 316092 42100 316098 42152
rect 227530 42032 227536 42084
rect 227588 42072 227594 42084
rect 260834 42072 260840 42084
rect 227588 42044 260840 42072
rect 227588 42032 227594 42044
rect 260834 42032 260840 42044
rect 260892 42032 260898 42084
rect 315942 42032 315948 42084
rect 316000 42072 316006 42084
rect 387794 42072 387800 42084
rect 316000 42044 387800 42072
rect 316000 42032 316006 42044
rect 387794 42032 387800 42044
rect 387852 42032 387858 42084
rect 424962 42032 424968 42084
rect 425020 42072 425026 42084
rect 545114 42072 545120 42084
rect 425020 42044 545120 42072
rect 425020 42032 425026 42044
rect 545114 42032 545120 42044
rect 545172 42032 545178 42084
rect 135438 41352 135444 41404
rect 135496 41392 135502 41404
rect 135622 41392 135628 41404
rect 135496 41364 135628 41392
rect 135496 41352 135502 41364
rect 135622 41352 135628 41364
rect 135680 41352 135686 41404
rect 478138 41352 478144 41404
rect 478196 41392 478202 41404
rect 580166 41392 580172 41404
rect 478196 41364 580172 41392
rect 478196 41352 478202 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 224770 40672 224776 40724
rect 224828 40712 224834 40724
rect 256694 40712 256700 40724
rect 224828 40684 256700 40712
rect 224828 40672 224834 40684
rect 256694 40672 256700 40684
rect 256752 40672 256758 40724
rect 263410 40672 263416 40724
rect 263468 40712 263474 40724
rect 313274 40712 313280 40724
rect 263468 40684 313280 40712
rect 263468 40672 263474 40684
rect 313274 40672 313280 40684
rect 313332 40672 313338 40724
rect 339402 40672 339408 40724
rect 339460 40712 339466 40724
rect 422294 40712 422300 40724
rect 339460 40684 422300 40712
rect 339460 40672 339466 40684
rect 422294 40672 422300 40684
rect 422352 40672 422358 40724
rect 296622 39380 296628 39432
rect 296680 39420 296686 39432
rect 360194 39420 360200 39432
rect 296680 39392 360200 39420
rect 296680 39380 296686 39392
rect 360194 39380 360200 39392
rect 360252 39380 360258 39432
rect 223482 39312 223488 39364
rect 223540 39352 223546 39364
rect 252554 39352 252560 39364
rect 223540 39324 252560 39352
rect 223540 39312 223546 39324
rect 252554 39312 252560 39324
rect 252612 39312 252618 39364
rect 262122 39312 262128 39364
rect 262180 39352 262186 39364
rect 309134 39352 309140 39364
rect 262180 39324 309140 39352
rect 262180 39312 262186 39324
rect 309134 39312 309140 39324
rect 309192 39312 309198 39364
rect 357342 39312 357348 39364
rect 357400 39352 357406 39364
rect 447134 39352 447140 39364
rect 357400 39324 447140 39352
rect 357400 39312 357406 39324
rect 447134 39312 447140 39324
rect 447192 39312 447198 39364
rect 449802 39312 449808 39364
rect 449860 39352 449866 39364
rect 574830 39352 574836 39364
rect 449860 39324 574836 39352
rect 449860 39312 449866 39324
rect 574830 39312 574836 39324
rect 574888 39312 574894 39364
rect 135533 38607 135591 38613
rect 135533 38573 135545 38607
rect 135579 38604 135591 38607
rect 135622 38604 135628 38616
rect 135579 38576 135628 38604
rect 135579 38573 135591 38576
rect 135533 38567 135591 38573
rect 135622 38564 135628 38576
rect 135680 38564 135686 38616
rect 220630 37884 220636 37936
rect 220688 37924 220694 37936
rect 249794 37924 249800 37936
rect 220688 37896 249800 37924
rect 220688 37884 220694 37896
rect 249794 37884 249800 37896
rect 249852 37884 249858 37936
rect 256602 37884 256608 37936
rect 256660 37924 256666 37936
rect 302234 37924 302240 37936
rect 256660 37896 302240 37924
rect 256660 37884 256666 37896
rect 302234 37884 302240 37896
rect 302292 37884 302298 37936
rect 335262 37884 335268 37936
rect 335320 37924 335326 37936
rect 415394 37924 415400 37936
rect 335320 37896 415400 37924
rect 335320 37884 335326 37896
rect 415394 37884 415400 37896
rect 415452 37884 415458 37936
rect 422202 37884 422208 37936
rect 422260 37924 422266 37936
rect 540974 37924 540980 37936
rect 422260 37896 540980 37924
rect 422260 37884 422266 37896
rect 540974 37884 540980 37896
rect 541032 37884 541038 37936
rect 250990 36592 250996 36644
rect 251048 36632 251054 36644
rect 295334 36632 295340 36644
rect 251048 36604 295340 36632
rect 251048 36592 251054 36604
rect 295334 36592 295340 36604
rect 295392 36592 295398 36644
rect 217962 36524 217968 36576
rect 218020 36564 218026 36576
rect 245654 36564 245660 36576
rect 218020 36536 245660 36564
rect 218020 36524 218026 36536
rect 245654 36524 245660 36536
rect 245712 36524 245718 36576
rect 284202 36524 284208 36576
rect 284260 36564 284266 36576
rect 342254 36564 342260 36576
rect 284260 36536 342260 36564
rect 284260 36524 284266 36536
rect 342254 36524 342260 36536
rect 342312 36524 342318 36576
rect 351822 36524 351828 36576
rect 351880 36564 351886 36576
rect 440234 36564 440240 36576
rect 351880 36536 440240 36564
rect 351880 36524 351886 36536
rect 440234 36524 440240 36536
rect 440292 36524 440298 36576
rect 444282 36524 444288 36576
rect 444340 36564 444346 36576
rect 572714 36564 572720 36576
rect 444340 36536 572720 36564
rect 444340 36524 444346 36536
rect 572714 36524 572720 36536
rect 572772 36524 572778 36576
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 11698 35884 11704 35896
rect 3476 35856 11704 35884
rect 3476 35844 3482 35856
rect 11698 35844 11704 35856
rect 11756 35844 11762 35896
rect 277302 35232 277308 35284
rect 277360 35272 277366 35284
rect 331306 35272 331312 35284
rect 277360 35244 331312 35272
rect 277360 35232 277366 35244
rect 331306 35232 331312 35244
rect 331364 35232 331370 35284
rect 215110 35164 215116 35216
rect 215168 35204 215174 35216
rect 242894 35204 242900 35216
rect 215168 35176 242900 35204
rect 215168 35164 215174 35176
rect 242894 35164 242900 35176
rect 242952 35164 242958 35216
rect 249702 35164 249708 35216
rect 249760 35204 249766 35216
rect 291194 35204 291200 35216
rect 249760 35176 291200 35204
rect 249760 35164 249766 35176
rect 291194 35164 291200 35176
rect 291252 35164 291258 35216
rect 327718 35164 327724 35216
rect 327776 35204 327782 35216
rect 400306 35204 400312 35216
rect 327776 35176 400312 35204
rect 327776 35164 327782 35176
rect 400306 35164 400312 35176
rect 400364 35164 400370 35216
rect 402882 35164 402888 35216
rect 402940 35204 402946 35216
rect 512086 35204 512092 35216
rect 402940 35176 512092 35204
rect 402940 35164 402946 35176
rect 512086 35164 512092 35176
rect 512144 35164 512150 35216
rect 241422 33736 241428 33788
rect 241480 33776 241486 33788
rect 280154 33776 280160 33788
rect 241480 33748 280160 33776
rect 241480 33736 241486 33748
rect 280154 33736 280160 33748
rect 280212 33736 280218 33788
rect 280798 33736 280804 33788
rect 280856 33776 280862 33788
rect 328454 33776 328460 33788
rect 280856 33748 328460 33776
rect 280856 33736 280862 33748
rect 328454 33736 328460 33748
rect 328512 33736 328518 33788
rect 329742 33736 329748 33788
rect 329800 33776 329806 33788
rect 408586 33776 408592 33788
rect 329800 33748 408592 33776
rect 329800 33736 329806 33748
rect 408586 33736 408592 33748
rect 408644 33736 408650 33788
rect 409782 33736 409788 33788
rect 409840 33776 409846 33788
rect 523034 33776 523040 33788
rect 409840 33748 523040 33776
rect 409840 33736 409846 33748
rect 523034 33736 523040 33748
rect 523092 33736 523098 33788
rect 240042 32444 240048 32496
rect 240100 32484 240106 32496
rect 277394 32484 277400 32496
rect 240100 32456 277400 32484
rect 240100 32444 240106 32456
rect 277394 32444 277400 32456
rect 277452 32444 277458 32496
rect 264882 32376 264888 32428
rect 264940 32416 264946 32428
rect 313366 32416 313372 32428
rect 264940 32388 313372 32416
rect 264940 32376 264946 32388
rect 313366 32376 313372 32388
rect 313424 32376 313430 32428
rect 314562 32376 314568 32428
rect 314620 32416 314626 32428
rect 386414 32416 386420 32428
rect 314620 32388 386420 32416
rect 314620 32376 314626 32388
rect 386414 32376 386420 32388
rect 386472 32376 386478 32428
rect 387702 32376 387708 32428
rect 387760 32416 387766 32428
rect 491294 32416 491300 32428
rect 387760 32388 491300 32416
rect 387760 32376 387766 32388
rect 491294 32376 491300 32388
rect 491352 32376 491358 32428
rect 237282 31084 237288 31136
rect 237340 31124 237346 31136
rect 273254 31124 273260 31136
rect 237340 31096 273260 31124
rect 237340 31084 237346 31096
rect 273254 31084 273260 31096
rect 273312 31084 273318 31136
rect 269022 31016 269028 31068
rect 269080 31056 269086 31068
rect 320174 31056 320180 31068
rect 269080 31028 320180 31056
rect 269080 31016 269086 31028
rect 320174 31016 320180 31028
rect 320232 31016 320238 31068
rect 326982 31016 326988 31068
rect 327040 31056 327046 31068
rect 404354 31056 404360 31068
rect 327040 31028 404360 31056
rect 327040 31016 327046 31028
rect 404354 31016 404360 31028
rect 404412 31016 404418 31068
rect 407022 31016 407028 31068
rect 407080 31056 407086 31068
rect 520366 31056 520372 31068
rect 407080 31028 520372 31056
rect 407080 31016 407086 31028
rect 520366 31016 520372 31028
rect 520424 31016 520430 31068
rect 453298 30268 453304 30320
rect 453356 30308 453362 30320
rect 580166 30308 580172 30320
rect 453356 30280 580172 30308
rect 453356 30268 453362 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 227622 29656 227628 29708
rect 227680 29696 227686 29708
rect 259454 29696 259460 29708
rect 227680 29668 259460 29696
rect 227680 29656 227686 29668
rect 259454 29656 259460 29668
rect 259512 29656 259518 29708
rect 252462 29588 252468 29640
rect 252520 29628 252526 29640
rect 296806 29628 296812 29640
rect 252520 29600 296812 29628
rect 252520 29588 252526 29600
rect 296806 29588 296812 29600
rect 296864 29588 296870 29640
rect 304902 29588 304908 29640
rect 304960 29628 304966 29640
rect 372614 29628 372620 29640
rect 304960 29600 372620 29628
rect 304960 29588 304966 29600
rect 372614 29588 372620 29600
rect 372672 29588 372678 29640
rect 135530 29016 135536 29028
rect 135491 28988 135536 29016
rect 135530 28976 135536 28988
rect 135588 28976 135594 29028
rect 224862 28228 224868 28280
rect 224920 28268 224926 28280
rect 255314 28268 255320 28280
rect 224920 28240 255320 28268
rect 224920 28228 224926 28240
rect 255314 28228 255320 28240
rect 255372 28228 255378 28280
rect 257338 28228 257344 28280
rect 257396 28268 257402 28280
rect 298094 28268 298100 28280
rect 257396 28240 298100 28268
rect 257396 28228 257402 28240
rect 298094 28228 298100 28240
rect 298152 28228 298158 28280
rect 303522 28228 303528 28280
rect 303580 28268 303586 28280
rect 368474 28268 368480 28280
rect 303580 28240 368480 28268
rect 303580 28228 303586 28240
rect 368474 28228 368480 28240
rect 368532 28228 368538 28280
rect 369762 28228 369768 28280
rect 369820 28268 369826 28280
rect 465074 28268 465080 28280
rect 369820 28240 465080 28268
rect 369820 28228 369826 28240
rect 465074 28228 465080 28240
rect 465132 28228 465138 28280
rect 216490 26868 216496 26920
rect 216548 26908 216554 26920
rect 244274 26908 244280 26920
rect 216548 26880 244280 26908
rect 216548 26868 216554 26880
rect 244274 26868 244280 26880
rect 244332 26868 244338 26920
rect 246942 26868 246948 26920
rect 247000 26908 247006 26920
rect 287054 26908 287060 26920
rect 247000 26880 287060 26908
rect 247000 26868 247006 26880
rect 287054 26868 287060 26880
rect 287112 26868 287118 26920
rect 298002 26868 298008 26920
rect 298060 26908 298066 26920
rect 361574 26908 361580 26920
rect 298060 26880 361580 26908
rect 298060 26868 298066 26880
rect 361574 26868 361580 26880
rect 361632 26868 361638 26920
rect 372522 26868 372528 26920
rect 372580 26908 372586 26920
rect 467926 26908 467932 26920
rect 372580 26880 467932 26908
rect 372580 26868 372586 26880
rect 467926 26868 467932 26880
rect 467984 26868 467990 26920
rect 212350 25576 212356 25628
rect 212408 25616 212414 25628
rect 237374 25616 237380 25628
rect 212408 25588 237380 25616
rect 212408 25576 212414 25588
rect 237374 25576 237380 25588
rect 237432 25576 237438 25628
rect 234522 25508 234528 25560
rect 234580 25548 234586 25560
rect 270586 25548 270592 25560
rect 234580 25520 270592 25548
rect 234580 25508 234586 25520
rect 270586 25508 270592 25520
rect 270644 25508 270650 25560
rect 292482 25508 292488 25560
rect 292540 25548 292546 25560
rect 354674 25548 354680 25560
rect 292540 25520 354680 25548
rect 292540 25508 292546 25520
rect 354674 25508 354680 25520
rect 354732 25508 354738 25560
rect 441522 25508 441528 25560
rect 441580 25548 441586 25560
rect 568574 25548 568580 25560
rect 441580 25520 568580 25548
rect 441580 25508 441586 25520
rect 568574 25508 568580 25520
rect 568632 25508 568638 25560
rect 206830 24080 206836 24132
rect 206888 24120 206894 24132
rect 230474 24120 230480 24132
rect 206888 24092 230480 24120
rect 206888 24080 206894 24092
rect 230474 24080 230480 24092
rect 230532 24080 230538 24132
rect 231670 24080 231676 24132
rect 231728 24120 231734 24132
rect 266354 24120 266360 24132
rect 231728 24092 266360 24120
rect 231728 24080 231734 24092
rect 266354 24080 266360 24092
rect 266412 24080 266418 24132
rect 282822 24080 282828 24132
rect 282880 24120 282886 24132
rect 339586 24120 339592 24132
rect 282880 24092 339592 24120
rect 282880 24080 282886 24092
rect 339586 24080 339592 24092
rect 339644 24080 339650 24132
rect 342162 24080 342168 24132
rect 342220 24120 342226 24132
rect 425146 24120 425152 24132
rect 342220 24092 425152 24120
rect 342220 24080 342226 24092
rect 425146 24080 425152 24092
rect 425204 24080 425210 24132
rect 431862 24080 431868 24132
rect 431920 24120 431926 24132
rect 554866 24120 554872 24132
rect 431920 24092 554872 24120
rect 431920 24080 431926 24092
rect 554866 24080 554872 24092
rect 554924 24080 554930 24132
rect 204070 22720 204076 22772
rect 204128 22760 204134 22772
rect 227806 22760 227812 22772
rect 204128 22732 227812 22760
rect 204128 22720 204134 22732
rect 227806 22720 227812 22732
rect 227864 22720 227870 22772
rect 228910 22720 228916 22772
rect 228968 22760 228974 22772
rect 262214 22760 262220 22772
rect 228968 22732 262220 22760
rect 228968 22720 228974 22732
rect 262214 22720 262220 22732
rect 262272 22720 262278 22772
rect 280062 22720 280068 22772
rect 280120 22760 280126 22772
rect 336734 22760 336740 22772
rect 280120 22732 336740 22760
rect 280120 22720 280126 22732
rect 336734 22720 336740 22732
rect 336792 22720 336798 22772
rect 338022 22720 338028 22772
rect 338080 22760 338086 22772
rect 418154 22760 418160 22772
rect 338080 22732 418160 22760
rect 338080 22720 338086 22732
rect 418154 22720 418160 22732
rect 418212 22720 418218 22772
rect 419442 22720 419448 22772
rect 419500 22760 419506 22772
rect 536926 22760 536932 22772
rect 419500 22732 536932 22760
rect 419500 22720 419506 22732
rect 536926 22720 536932 22732
rect 536984 22720 536990 22772
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 128998 22080 129004 22092
rect 3200 22052 129004 22080
rect 3200 22040 3206 22052
rect 128998 22040 129004 22052
rect 129056 22040 129062 22092
rect 135438 22040 135444 22092
rect 135496 22080 135502 22092
rect 135622 22080 135628 22092
rect 135496 22052 135628 22080
rect 135496 22040 135502 22052
rect 135622 22040 135628 22052
rect 135680 22040 135686 22092
rect 202690 21428 202696 21480
rect 202748 21468 202754 21480
rect 223574 21468 223580 21480
rect 202748 21440 223580 21468
rect 202748 21428 202754 21440
rect 223574 21428 223580 21440
rect 223632 21428 223638 21480
rect 278682 21428 278688 21480
rect 278740 21468 278746 21480
rect 332594 21468 332600 21480
rect 278740 21440 332600 21468
rect 278740 21428 278746 21440
rect 332594 21428 332600 21440
rect 332652 21428 332658 21480
rect 222838 21360 222844 21412
rect 222896 21400 222902 21412
rect 252646 21400 252652 21412
rect 222896 21372 252652 21400
rect 222896 21360 222902 21372
rect 252646 21360 252652 21372
rect 252704 21360 252710 21412
rect 332502 21360 332508 21412
rect 332560 21400 332566 21412
rect 411254 21400 411260 21412
rect 332560 21372 411260 21400
rect 332560 21360 332566 21372
rect 411254 21360 411260 21372
rect 411312 21360 411318 21412
rect 412542 21360 412548 21412
rect 412600 21400 412606 21412
rect 527174 21400 527180 21412
rect 412600 21372 527180 21400
rect 412600 21360 412606 21372
rect 527174 21360 527180 21372
rect 527232 21360 527238 21412
rect 200758 20000 200764 20052
rect 200816 20040 200822 20052
rect 219434 20040 219440 20052
rect 200816 20012 219440 20040
rect 200816 20000 200822 20012
rect 219434 20000 219440 20012
rect 219492 20000 219498 20052
rect 219250 19932 219256 19984
rect 219308 19972 219314 19984
rect 248414 19972 248420 19984
rect 219308 19944 248420 19972
rect 219308 19932 219314 19944
rect 248414 19932 248420 19944
rect 248472 19932 248478 19984
rect 266262 19932 266268 19984
rect 266320 19972 266326 19984
rect 314654 19972 314660 19984
rect 266320 19944 314660 19972
rect 266320 19932 266326 19944
rect 314654 19932 314660 19944
rect 314712 19932 314718 19984
rect 317322 19932 317328 19984
rect 317380 19972 317386 19984
rect 390646 19972 390652 19984
rect 317380 19944 390652 19972
rect 317380 19932 317386 19944
rect 390646 19932 390652 19944
rect 390704 19932 390710 19984
rect 429102 19932 429108 19984
rect 429160 19972 429166 19984
rect 550634 19972 550640 19984
rect 429160 19944 550640 19972
rect 429160 19932 429166 19944
rect 550634 19932 550640 19944
rect 550692 19932 550698 19984
rect 135622 19292 135628 19304
rect 135583 19264 135628 19292
rect 135622 19252 135628 19264
rect 135680 19252 135686 19304
rect 301498 19252 301504 19304
rect 301556 19292 301562 19304
rect 305086 19292 305092 19304
rect 301556 19264 305092 19292
rect 301556 19252 301562 19264
rect 305086 19252 305092 19264
rect 305144 19252 305150 19304
rect 197262 18640 197268 18692
rect 197320 18680 197326 18692
rect 216674 18680 216680 18692
rect 197320 18652 216680 18680
rect 197320 18640 197326 18652
rect 216674 18640 216680 18652
rect 216732 18640 216738 18692
rect 215202 18572 215208 18624
rect 215260 18612 215266 18624
rect 241514 18612 241520 18624
rect 215260 18584 241520 18612
rect 215260 18572 215266 18584
rect 241514 18572 241520 18584
rect 241572 18572 241578 18624
rect 251082 18572 251088 18624
rect 251140 18612 251146 18624
rect 293954 18612 293960 18624
rect 251140 18584 293960 18612
rect 251140 18572 251146 18584
rect 293954 18572 293960 18584
rect 294012 18572 294018 18624
rect 310422 18572 310428 18624
rect 310480 18612 310486 18624
rect 379514 18612 379520 18624
rect 310480 18584 379520 18612
rect 310480 18572 310486 18584
rect 379514 18572 379520 18584
rect 379572 18572 379578 18624
rect 400122 18572 400128 18624
rect 400180 18612 400186 18624
rect 509234 18612 509240 18624
rect 400180 18584 509240 18612
rect 400180 18572 400186 18584
rect 509234 18572 509240 18584
rect 509292 18572 509298 18624
rect 483658 17892 483664 17944
rect 483716 17932 483722 17944
rect 579798 17932 579804 17944
rect 483716 17904 579804 17932
rect 483716 17892 483722 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 194410 17280 194416 17332
rect 194468 17320 194474 17332
rect 212534 17320 212540 17332
rect 194468 17292 212540 17320
rect 194468 17280 194474 17292
rect 212534 17280 212540 17292
rect 212592 17280 212598 17332
rect 209682 17212 209688 17264
rect 209740 17252 209746 17264
rect 234614 17252 234620 17264
rect 209740 17224 234620 17252
rect 209740 17212 209746 17224
rect 234614 17212 234620 17224
rect 234672 17212 234678 17264
rect 244182 17212 244188 17264
rect 244240 17252 244246 17264
rect 282914 17252 282920 17264
rect 244240 17224 282920 17252
rect 244240 17212 244246 17224
rect 282914 17212 282920 17224
rect 282972 17212 282978 17264
rect 285582 17212 285588 17264
rect 285640 17252 285646 17264
rect 343634 17252 343640 17264
rect 285640 17224 343640 17252
rect 285640 17212 285646 17224
rect 343634 17212 343640 17224
rect 343692 17212 343698 17264
rect 344922 17212 344928 17264
rect 344980 17252 344986 17264
rect 429194 17252 429200 17264
rect 344980 17224 429200 17252
rect 344980 17212 344986 17224
rect 429194 17212 429200 17224
rect 429252 17212 429258 17264
rect 255222 15920 255228 15972
rect 255280 15960 255286 15972
rect 300854 15960 300860 15972
rect 255280 15932 300860 15960
rect 255280 15920 255286 15932
rect 300854 15920 300860 15932
rect 300912 15920 300918 15972
rect 191650 15852 191656 15904
rect 191708 15892 191714 15904
rect 209866 15892 209872 15904
rect 191708 15864 209872 15892
rect 191708 15852 191714 15864
rect 209866 15852 209872 15864
rect 209924 15852 209930 15904
rect 220722 15852 220728 15904
rect 220780 15892 220786 15904
rect 251174 15892 251180 15904
rect 220780 15864 251180 15892
rect 220780 15852 220786 15864
rect 251174 15852 251180 15864
rect 251232 15852 251238 15904
rect 300762 15852 300768 15904
rect 300820 15892 300826 15904
rect 365806 15892 365812 15904
rect 300820 15864 365812 15892
rect 300820 15852 300826 15864
rect 365806 15852 365812 15864
rect 365864 15852 365870 15904
rect 390462 15852 390468 15904
rect 390520 15892 390526 15904
rect 494146 15892 494152 15904
rect 390520 15864 494152 15892
rect 390520 15852 390526 15864
rect 494146 15852 494152 15864
rect 494204 15852 494210 15904
rect 190270 14424 190276 14476
rect 190328 14464 190334 14476
rect 205634 14464 205640 14476
rect 190328 14436 205640 14464
rect 190328 14424 190334 14436
rect 205634 14424 205640 14436
rect 205692 14424 205698 14476
rect 216582 14424 216588 14476
rect 216640 14464 216646 14476
rect 244366 14464 244372 14476
rect 216640 14436 244372 14464
rect 216640 14424 216646 14436
rect 244366 14424 244372 14436
rect 244424 14424 244430 14476
rect 245562 14424 245568 14476
rect 245620 14464 245626 14476
rect 287146 14464 287152 14476
rect 245620 14436 287152 14464
rect 245620 14424 245626 14436
rect 287146 14424 287152 14436
rect 287204 14424 287210 14476
rect 288342 14424 288348 14476
rect 288400 14464 288406 14476
rect 347866 14464 347872 14476
rect 288400 14436 347872 14464
rect 288400 14424 288406 14436
rect 347866 14424 347872 14436
rect 347924 14424 347930 14476
rect 350442 14424 350448 14476
rect 350500 14464 350506 14476
rect 436094 14464 436100 14476
rect 350500 14436 436100 14464
rect 350500 14424 350506 14436
rect 436094 14424 436100 14436
rect 436152 14424 436158 14476
rect 437382 14424 437388 14476
rect 437440 14464 437446 14476
rect 563146 14464 563152 14476
rect 437440 14436 563152 14464
rect 437440 14424 437446 14436
rect 563146 14424 563152 14436
rect 563204 14424 563210 14476
rect 208210 13132 208216 13184
rect 208268 13172 208274 13184
rect 233234 13172 233240 13184
rect 208268 13144 233240 13172
rect 208268 13132 208274 13144
rect 233234 13132 233240 13144
rect 233292 13132 233298 13184
rect 187510 13064 187516 13116
rect 187568 13104 187574 13116
rect 201494 13104 201500 13116
rect 187568 13076 201500 13104
rect 187568 13064 187574 13076
rect 201494 13064 201500 13076
rect 201552 13064 201558 13116
rect 233142 13064 233148 13116
rect 233200 13104 233206 13116
rect 269114 13104 269120 13116
rect 233200 13076 269120 13104
rect 233200 13064 233206 13076
rect 269114 13064 269120 13076
rect 269172 13064 269178 13116
rect 270402 13064 270408 13116
rect 270460 13104 270466 13116
rect 321646 13104 321652 13116
rect 270460 13076 321652 13104
rect 270460 13064 270466 13076
rect 321646 13064 321652 13076
rect 321704 13064 321710 13116
rect 322842 13064 322848 13116
rect 322900 13104 322906 13116
rect 397454 13104 397460 13116
rect 322900 13076 397460 13104
rect 322900 13064 322906 13076
rect 397454 13064 397460 13076
rect 397512 13064 397518 13116
rect 416682 13064 416688 13116
rect 416740 13104 416746 13116
rect 532694 13104 532700 13116
rect 416740 13076 532700 13104
rect 416740 13064 416746 13076
rect 532694 13064 532700 13076
rect 532752 13064 532758 13116
rect 135622 12288 135628 12300
rect 135583 12260 135628 12288
rect 135622 12248 135628 12260
rect 135680 12248 135686 12300
rect 184842 11704 184848 11756
rect 184900 11744 184906 11756
rect 198734 11744 198740 11756
rect 184900 11716 198740 11744
rect 184900 11704 184906 11716
rect 198734 11704 198740 11716
rect 198792 11704 198798 11756
rect 204162 11704 204168 11756
rect 204220 11744 204226 11756
rect 226334 11744 226340 11756
rect 204220 11716 226340 11744
rect 204220 11704 204226 11716
rect 226334 11704 226340 11716
rect 226392 11704 226398 11756
rect 229002 11704 229008 11756
rect 229060 11744 229066 11756
rect 262306 11744 262312 11756
rect 229060 11716 262312 11744
rect 229060 11704 229066 11716
rect 262306 11704 262312 11716
rect 262364 11704 262370 11756
rect 263502 11704 263508 11756
rect 263560 11744 263566 11756
rect 311894 11744 311900 11756
rect 263560 11716 311900 11744
rect 263560 11704 263566 11716
rect 311894 11704 311900 11716
rect 311952 11704 311958 11756
rect 313182 11704 313188 11756
rect 313240 11744 313246 11756
rect 382366 11744 382372 11756
rect 313240 11716 382372 11744
rect 313240 11704 313246 11716
rect 382366 11704 382372 11716
rect 382424 11704 382430 11756
rect 404262 11704 404268 11756
rect 404320 11744 404326 11756
rect 514754 11744 514760 11756
rect 404320 11716 514760 11744
rect 404320 11704 404326 11716
rect 514754 11704 514760 11716
rect 514812 11704 514818 11756
rect 188982 10276 188988 10328
rect 189040 10316 189046 10328
rect 204254 10316 204260 10328
rect 189040 10288 204260 10316
rect 189040 10276 189046 10288
rect 204254 10276 204260 10288
rect 204312 10276 204318 10328
rect 206922 10276 206928 10328
rect 206980 10316 206986 10328
rect 229094 10316 229100 10328
rect 206980 10288 229100 10316
rect 206980 10276 206986 10288
rect 229094 10276 229100 10288
rect 229152 10276 229158 10328
rect 231762 10276 231768 10328
rect 231820 10316 231826 10328
rect 264974 10316 264980 10328
rect 231820 10288 264980 10316
rect 231820 10276 231826 10288
rect 264974 10276 264980 10288
rect 265032 10276 265038 10328
rect 267642 10276 267648 10328
rect 267700 10316 267706 10328
rect 318794 10316 318800 10328
rect 267700 10288 318800 10316
rect 267700 10276 267706 10288
rect 318794 10276 318800 10288
rect 318852 10276 318858 10328
rect 320082 10276 320088 10328
rect 320140 10316 320146 10328
rect 393314 10316 393320 10328
rect 320140 10288 393320 10316
rect 320140 10276 320146 10288
rect 393314 10276 393320 10288
rect 393372 10276 393378 10328
rect 394602 10276 394608 10328
rect 394660 10316 394666 10328
rect 502426 10316 502432 10328
rect 394660 10288 502432 10316
rect 394660 10276 394666 10288
rect 502426 10276 502432 10288
rect 502484 10276 502490 10328
rect 186130 8984 186136 9036
rect 186188 9024 186194 9036
rect 201586 9024 201592 9036
rect 186188 8996 201592 9024
rect 186188 8984 186194 8996
rect 201586 8984 201592 8996
rect 201644 8984 201650 9036
rect 201402 8916 201408 8968
rect 201460 8956 201466 8968
rect 222930 8956 222936 8968
rect 201460 8928 222936 8956
rect 201460 8916 201466 8928
rect 222930 8916 222936 8928
rect 222988 8916 222994 8968
rect 226242 8916 226248 8968
rect 226300 8956 226306 8968
rect 258626 8956 258632 8968
rect 226300 8928 258632 8956
rect 226300 8916 226306 8928
rect 258626 8916 258632 8928
rect 258684 8916 258690 8968
rect 260742 8916 260748 8968
rect 260800 8956 260806 8968
rect 308582 8956 308588 8968
rect 260800 8928 308588 8956
rect 260800 8916 260806 8928
rect 308582 8916 308588 8928
rect 308640 8916 308646 8968
rect 309778 8916 309784 8968
rect 309836 8956 309842 8968
rect 376386 8956 376392 8968
rect 309836 8928 376392 8956
rect 309836 8916 309842 8928
rect 376386 8916 376392 8928
rect 376444 8916 376450 8968
rect 381538 8916 381544 8968
rect 381596 8956 381602 8968
rect 451366 8956 451372 8968
rect 381596 8928 451372 8956
rect 381596 8916 381602 8928
rect 451366 8916 451372 8928
rect 451424 8916 451430 8968
rect 456058 8916 456064 8968
rect 456116 8956 456122 8968
rect 579798 8956 579804 8968
rect 456116 8928 579804 8956
rect 456116 8916 456122 8928
rect 579798 8916 579804 8928
rect 579856 8916 579862 8968
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 10318 8276 10324 8288
rect 3476 8248 10324 8276
rect 3476 8236 3482 8248
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 183370 7556 183376 7608
rect 183428 7596 183434 7608
rect 197998 7596 198004 7608
rect 183428 7568 198004 7596
rect 183428 7556 183434 7568
rect 197998 7556 198004 7568
rect 198056 7556 198062 7608
rect 198550 7556 198556 7608
rect 198608 7596 198614 7608
rect 198608 7568 209820 7596
rect 198608 7556 198614 7568
rect 209792 7528 209820 7568
rect 219342 7556 219348 7608
rect 219400 7596 219406 7608
rect 247954 7596 247960 7608
rect 219400 7568 247960 7596
rect 219400 7556 219406 7568
rect 247954 7556 247960 7568
rect 248012 7556 248018 7608
rect 248322 7556 248328 7608
rect 248380 7596 248386 7608
rect 290734 7596 290740 7608
rect 248380 7568 290740 7596
rect 248380 7556 248386 7568
rect 290734 7556 290740 7568
rect 290792 7556 290798 7608
rect 291102 7556 291108 7608
rect 291160 7596 291166 7608
rect 351362 7596 351368 7608
rect 291160 7568 351368 7596
rect 291160 7556 291166 7568
rect 351362 7556 351368 7568
rect 351420 7556 351426 7608
rect 354582 7556 354588 7608
rect 354640 7596 354646 7608
rect 444190 7596 444196 7608
rect 354640 7568 444196 7596
rect 354640 7556 354646 7568
rect 444190 7556 444196 7568
rect 444248 7556 444254 7608
rect 451918 7556 451924 7608
rect 451976 7596 451982 7608
rect 576210 7596 576216 7608
rect 451976 7568 576216 7596
rect 451976 7556 451982 7568
rect 576210 7556 576216 7568
rect 576268 7556 576274 7608
rect 209792 7500 219480 7528
rect 219342 7352 219348 7404
rect 219400 7392 219406 7404
rect 219452 7392 219480 7500
rect 219400 7364 219480 7392
rect 219400 7352 219406 7364
rect 273162 6196 273168 6248
rect 273220 6236 273226 6248
rect 326430 6236 326436 6248
rect 273220 6208 326436 6236
rect 273220 6196 273226 6208
rect 326430 6196 326436 6208
rect 326488 6196 326494 6248
rect 179230 6128 179236 6180
rect 179288 6168 179294 6180
rect 190822 6168 190828 6180
rect 179288 6140 190828 6168
rect 179288 6128 179294 6140
rect 190822 6128 190828 6140
rect 190880 6128 190886 6180
rect 191742 6128 191748 6180
rect 191800 6168 191806 6180
rect 208670 6168 208676 6180
rect 191800 6140 208676 6168
rect 191800 6128 191806 6140
rect 208670 6128 208676 6140
rect 208728 6128 208734 6180
rect 210970 6128 210976 6180
rect 211028 6168 211034 6180
rect 237190 6168 237196 6180
rect 211028 6140 237196 6168
rect 211028 6128 211034 6140
rect 237190 6128 237196 6140
rect 237248 6128 237254 6180
rect 238662 6128 238668 6180
rect 238720 6168 238726 6180
rect 276474 6168 276480 6180
rect 238720 6140 276480 6168
rect 238720 6128 238726 6140
rect 276474 6128 276480 6140
rect 276532 6128 276538 6180
rect 311802 6128 311808 6180
rect 311860 6168 311866 6180
rect 381170 6168 381176 6180
rect 311860 6140 381176 6168
rect 311860 6128 311866 6140
rect 381170 6128 381176 6140
rect 381228 6128 381234 6180
rect 391842 6128 391848 6180
rect 391900 6168 391906 6180
rect 497734 6168 497740 6180
rect 391900 6140 497740 6168
rect 391900 6128 391906 6140
rect 497734 6128 497740 6140
rect 497792 6128 497798 6180
rect 275922 4836 275928 4888
rect 275980 4876 275986 4888
rect 330018 4876 330024 4888
rect 275980 4848 330024 4876
rect 275980 4836 275986 4848
rect 330018 4836 330024 4848
rect 330076 4836 330082 4888
rect 352558 4836 352564 4888
rect 352616 4876 352622 4888
rect 358538 4876 358544 4888
rect 352616 4848 358544 4876
rect 352616 4836 352622 4848
rect 358538 4836 358544 4848
rect 358596 4836 358602 4888
rect 173710 4768 173716 4820
rect 173768 4808 173774 4820
rect 183738 4808 183744 4820
rect 173768 4780 183744 4808
rect 173768 4768 173774 4780
rect 183738 4768 183744 4780
rect 183796 4768 183802 4820
rect 194502 4768 194508 4820
rect 194560 4808 194566 4820
rect 212258 4808 212264 4820
rect 194560 4780 212264 4808
rect 194560 4768 194566 4780
rect 212258 4768 212264 4780
rect 212316 4768 212322 4820
rect 221458 4768 221464 4820
rect 221516 4808 221522 4820
rect 240778 4808 240784 4820
rect 221516 4780 240784 4808
rect 221516 4768 221522 4780
rect 240778 4768 240784 4780
rect 240836 4768 240842 4820
rect 242158 4768 242164 4820
rect 242216 4808 242222 4820
rect 255038 4808 255044 4820
rect 242216 4780 255044 4808
rect 242216 4768 242222 4780
rect 255038 4768 255044 4780
rect 255096 4768 255102 4820
rect 255958 4768 255964 4820
rect 256016 4808 256022 4820
rect 280062 4808 280068 4820
rect 256016 4780 280068 4808
rect 256016 4768 256022 4780
rect 280062 4768 280068 4780
rect 280120 4768 280126 4820
rect 309042 4768 309048 4820
rect 309100 4808 309106 4820
rect 378778 4808 378784 4820
rect 309100 4780 378784 4808
rect 309100 4768 309106 4780
rect 378778 4768 378784 4780
rect 378836 4768 378842 4820
rect 382182 4768 382188 4820
rect 382240 4808 382246 4820
rect 483474 4808 483480 4820
rect 382240 4780 483480 4808
rect 382240 4768 382246 4780
rect 483474 4768 483480 4780
rect 483532 4768 483538 4820
rect 184198 4156 184204 4208
rect 184256 4196 184262 4208
rect 187234 4196 187240 4208
rect 184256 4168 187240 4196
rect 184256 4156 184262 4168
rect 187234 4156 187240 4168
rect 187292 4156 187298 4208
rect 192478 4156 192484 4208
rect 192536 4196 192542 4208
rect 194410 4196 194416 4208
rect 192536 4168 194416 4196
rect 192536 4156 192542 4168
rect 194410 4156 194416 4168
rect 194468 4156 194474 4208
rect 213178 4156 213184 4208
rect 213236 4196 213242 4208
rect 215846 4196 215852 4208
rect 213236 4168 215852 4196
rect 213236 4156 213242 4168
rect 215846 4156 215852 4168
rect 215904 4156 215910 4208
rect 408494 4156 408500 4208
rect 408552 4196 408558 4208
rect 409690 4196 409696 4208
rect 408552 4168 409696 4196
rect 408552 4156 408558 4168
rect 409690 4156 409696 4168
rect 409748 4156 409754 4208
rect 425146 4156 425152 4208
rect 425204 4196 425210 4208
rect 426342 4196 426348 4208
rect 425204 4168 426348 4196
rect 425204 4156 425210 4168
rect 426342 4156 426348 4168
rect 426400 4156 426406 4208
rect 451274 4156 451280 4208
rect 451332 4196 451338 4208
rect 452470 4196 452476 4208
rect 451332 4168 452476 4196
rect 451332 4156 451338 4168
rect 452470 4156 452476 4168
rect 452528 4156 452534 4208
rect 127802 4088 127808 4140
rect 127860 4128 127866 4140
rect 133874 4128 133880 4140
rect 127860 4100 133880 4128
rect 127860 4088 127866 4100
rect 133874 4088 133880 4100
rect 133932 4088 133938 4140
rect 142062 4088 142068 4140
rect 142120 4128 142126 4140
rect 143534 4128 143540 4140
rect 142120 4100 143540 4128
rect 142120 4088 142126 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
rect 160002 4088 160008 4140
rect 160060 4128 160066 4140
rect 163498 4128 163504 4140
rect 160060 4100 163504 4128
rect 160060 4088 160066 4100
rect 163498 4088 163504 4100
rect 163556 4088 163562 4140
rect 166902 4088 166908 4140
rect 166960 4128 166966 4140
rect 172974 4128 172980 4140
rect 166960 4100 172980 4128
rect 166960 4088 166966 4100
rect 172974 4088 172980 4100
rect 173032 4088 173038 4140
rect 212537 4131 212595 4137
rect 212537 4097 212549 4131
rect 212583 4128 212595 4131
rect 217321 4131 217379 4137
rect 217321 4128 217333 4131
rect 212583 4100 217333 4128
rect 212583 4097 212595 4100
rect 212537 4091 212595 4097
rect 217321 4097 217333 4100
rect 217367 4097 217379 4131
rect 217321 4091 217379 4097
rect 361482 4088 361488 4140
rect 361540 4128 361546 4140
rect 453666 4128 453672 4140
rect 361540 4100 453672 4128
rect 361540 4088 361546 4100
rect 453666 4088 453672 4100
rect 453724 4088 453730 4140
rect 574738 4088 574744 4140
rect 574796 4128 574802 4140
rect 577406 4128 577412 4140
rect 574796 4100 577412 4128
rect 574796 4088 574802 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 130194 4020 130200 4072
rect 130252 4060 130258 4072
rect 135622 4060 135628 4072
rect 130252 4032 135628 4060
rect 130252 4020 130258 4032
rect 135622 4020 135628 4032
rect 135680 4020 135686 4072
rect 139670 4020 139676 4072
rect 139728 4060 139734 4072
rect 142430 4060 142436 4072
rect 139728 4032 142436 4060
rect 139728 4020 139734 4032
rect 142430 4020 142436 4032
rect 142488 4020 142494 4072
rect 159910 4020 159916 4072
rect 159968 4060 159974 4072
rect 162302 4060 162308 4072
rect 159968 4032 162308 4060
rect 159968 4020 159974 4032
rect 162302 4020 162308 4032
rect 162360 4020 162366 4072
rect 176562 4020 176568 4072
rect 176620 4060 176626 4072
rect 186038 4060 186044 4072
rect 176620 4032 186044 4060
rect 176620 4020 176626 4032
rect 186038 4020 186044 4032
rect 186096 4020 186102 4072
rect 367002 4020 367008 4072
rect 367060 4060 367066 4072
rect 460842 4060 460848 4072
rect 367060 4032 460848 4060
rect 367060 4020 367066 4032
rect 460842 4020 460848 4032
rect 460900 4020 460906 4072
rect 128998 3952 129004 4004
rect 129056 3992 129062 4004
rect 135254 3992 135260 4004
rect 129056 3964 135260 3992
rect 129056 3952 129062 3964
rect 135254 3952 135260 3964
rect 135312 3952 135318 4004
rect 140866 3952 140872 4004
rect 140924 3992 140930 4004
rect 143626 3992 143632 4004
rect 140924 3964 143632 3992
rect 140924 3952 140930 3964
rect 143626 3952 143632 3964
rect 143684 3952 143690 4004
rect 175182 3952 175188 4004
rect 175240 3992 175246 4004
rect 184842 3992 184848 4004
rect 175240 3964 184848 3992
rect 175240 3952 175246 3964
rect 184842 3952 184848 3964
rect 184900 3952 184906 4004
rect 205542 3952 205548 4004
rect 205600 3992 205606 4004
rect 212537 3995 212595 4001
rect 212537 3992 212549 3995
rect 205600 3964 212549 3992
rect 205600 3952 205606 3964
rect 212537 3961 212549 3964
rect 212583 3961 212595 3995
rect 212537 3955 212595 3961
rect 364242 3952 364248 4004
rect 364300 3992 364306 4004
rect 457254 3992 457260 4004
rect 364300 3964 457260 3992
rect 364300 3952 364306 3964
rect 457254 3952 457260 3964
rect 457312 3952 457318 4004
rect 138474 3884 138480 3936
rect 138532 3924 138538 3936
rect 142154 3924 142160 3936
rect 138532 3896 142160 3924
rect 138532 3884 138538 3896
rect 142154 3884 142160 3896
rect 142212 3884 142218 3936
rect 169570 3884 169576 3936
rect 169628 3924 169634 3936
rect 176562 3924 176568 3936
rect 169628 3896 176568 3924
rect 169628 3884 169634 3896
rect 176562 3884 176568 3896
rect 176620 3884 176626 3936
rect 177850 3884 177856 3936
rect 177908 3924 177914 3936
rect 188430 3924 188436 3936
rect 177908 3896 188436 3924
rect 177908 3884 177914 3896
rect 188430 3884 188436 3896
rect 188488 3884 188494 3936
rect 195882 3884 195888 3936
rect 195940 3924 195946 3936
rect 214650 3924 214656 3936
rect 195940 3896 214656 3924
rect 195940 3884 195946 3896
rect 214650 3884 214656 3896
rect 214708 3884 214714 3936
rect 368382 3884 368388 3936
rect 368440 3924 368446 3936
rect 464430 3924 464436 3936
rect 368440 3896 464436 3924
rect 368440 3884 368446 3896
rect 464430 3884 464436 3896
rect 464488 3884 464494 3936
rect 168190 3816 168196 3868
rect 168248 3856 168254 3868
rect 174170 3856 174176 3868
rect 168248 3828 174176 3856
rect 168248 3816 168254 3828
rect 174170 3816 174176 3828
rect 174228 3816 174234 3868
rect 182082 3816 182088 3868
rect 182140 3856 182146 3868
rect 195606 3856 195612 3868
rect 182140 3828 195612 3856
rect 182140 3816 182146 3828
rect 195606 3816 195612 3828
rect 195664 3816 195670 3868
rect 198642 3816 198648 3868
rect 198700 3856 198706 3868
rect 218146 3856 218152 3868
rect 198700 3828 218152 3856
rect 198700 3816 198706 3828
rect 218146 3816 218152 3828
rect 218204 3816 218210 3868
rect 371142 3816 371148 3868
rect 371200 3856 371206 3868
rect 467834 3856 467840 3868
rect 371200 3828 467840 3856
rect 371200 3816 371206 3828
rect 467834 3816 467840 3828
rect 467892 3816 467898 3868
rect 169662 3748 169668 3800
rect 169720 3788 169726 3800
rect 177758 3788 177764 3800
rect 169720 3760 177764 3788
rect 169720 3748 169726 3760
rect 177758 3748 177764 3760
rect 177816 3748 177822 3800
rect 183462 3748 183468 3800
rect 183520 3788 183526 3800
rect 196802 3788 196808 3800
rect 183520 3760 196808 3788
rect 183520 3748 183526 3760
rect 196802 3748 196808 3760
rect 196860 3748 196866 3800
rect 200022 3748 200028 3800
rect 200080 3788 200086 3800
rect 213089 3791 213147 3797
rect 213089 3788 213101 3791
rect 200080 3760 213101 3788
rect 200080 3748 200086 3760
rect 213089 3757 213101 3760
rect 213135 3757 213147 3791
rect 213089 3751 213147 3757
rect 373902 3748 373908 3800
rect 373960 3788 373966 3800
rect 471514 3788 471520 3800
rect 373960 3760 471520 3788
rect 373960 3748 373966 3760
rect 471514 3748 471520 3760
rect 471572 3748 471578 3800
rect 126606 3680 126612 3732
rect 126664 3720 126670 3732
rect 133966 3720 133972 3732
rect 126664 3692 133972 3720
rect 126664 3680 126670 3692
rect 133966 3680 133972 3692
rect 134024 3680 134030 3732
rect 180702 3680 180708 3732
rect 180760 3720 180766 3732
rect 193214 3720 193220 3732
rect 180760 3692 193220 3720
rect 180760 3680 180766 3692
rect 193214 3680 193220 3692
rect 193272 3680 193278 3732
rect 202782 3680 202788 3732
rect 202840 3720 202846 3732
rect 202840 3692 204024 3720
rect 202840 3680 202846 3692
rect 172422 3612 172428 3664
rect 172480 3652 172486 3664
rect 181346 3652 181352 3664
rect 172480 3624 181352 3652
rect 172480 3612 172486 3624
rect 181346 3612 181352 3624
rect 181404 3612 181410 3664
rect 186222 3612 186228 3664
rect 186280 3652 186286 3664
rect 200390 3652 200396 3664
rect 186280 3624 200396 3652
rect 186280 3612 186286 3624
rect 200390 3612 200396 3624
rect 200448 3612 200454 3664
rect 203886 3652 203892 3664
rect 201420 3624 203892 3652
rect 146846 3544 146852 3596
rect 146904 3584 146910 3596
rect 147766 3584 147772 3596
rect 146904 3556 147772 3584
rect 146904 3544 146910 3556
rect 147766 3544 147772 3556
rect 147824 3544 147830 3596
rect 161382 3544 161388 3596
rect 161440 3584 161446 3596
rect 164694 3584 164700 3596
rect 161440 3556 164700 3584
rect 161440 3544 161446 3556
rect 164694 3544 164700 3556
rect 164752 3544 164758 3596
rect 173802 3544 173808 3596
rect 173860 3584 173866 3596
rect 182542 3584 182548 3596
rect 173860 3556 182548 3584
rect 173860 3544 173866 3556
rect 182542 3544 182548 3556
rect 182600 3544 182606 3596
rect 187602 3544 187608 3596
rect 187660 3584 187666 3596
rect 201420 3584 201448 3624
rect 203886 3612 203892 3624
rect 203944 3612 203950 3664
rect 203996 3652 204024 3692
rect 208302 3680 208308 3732
rect 208360 3720 208366 3732
rect 217321 3723 217379 3729
rect 208360 3692 214604 3720
rect 208360 3680 208366 3692
rect 214469 3655 214527 3661
rect 214469 3652 214481 3655
rect 203996 3624 214481 3652
rect 214469 3621 214481 3624
rect 214515 3621 214527 3655
rect 214469 3615 214527 3621
rect 187660 3556 201448 3584
rect 187660 3544 187666 3556
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 214576 3584 214604 3692
rect 217321 3689 217333 3723
rect 217367 3720 217379 3723
rect 228910 3720 228916 3732
rect 217367 3692 228916 3720
rect 217367 3689 217379 3692
rect 217321 3683 217379 3689
rect 228910 3680 228916 3692
rect 228968 3680 228974 3732
rect 376662 3680 376668 3732
rect 376720 3720 376726 3732
rect 475102 3720 475108 3732
rect 376720 3692 475108 3720
rect 376720 3680 376726 3692
rect 475102 3680 475108 3692
rect 475160 3680 475166 3732
rect 214653 3655 214711 3661
rect 214653 3621 214665 3655
rect 214699 3652 214711 3655
rect 225322 3652 225328 3664
rect 214699 3624 225328 3652
rect 214699 3621 214711 3624
rect 214653 3615 214711 3621
rect 225322 3612 225328 3624
rect 225380 3612 225386 3664
rect 379422 3612 379428 3664
rect 379480 3652 379486 3664
rect 478690 3652 478696 3664
rect 379480 3624 478696 3652
rect 379480 3612 379486 3624
rect 478690 3612 478696 3624
rect 478748 3612 478754 3664
rect 574830 3612 574836 3664
rect 574888 3652 574894 3664
rect 580994 3652 581000 3664
rect 574888 3624 581000 3652
rect 574888 3612 574894 3624
rect 580994 3612 581000 3624
rect 581052 3612 581058 3664
rect 232498 3584 232504 3596
rect 214576 3556 232504 3584
rect 232498 3544 232504 3556
rect 232556 3544 232562 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 263410 3584 263416 3596
rect 262272 3556 263416 3584
rect 262272 3544 262278 3556
rect 263410 3544 263416 3556
rect 263468 3544 263474 3596
rect 270494 3544 270500 3596
rect 270552 3584 270558 3596
rect 271690 3584 271696 3596
rect 270552 3556 271696 3584
rect 270552 3544 270558 3556
rect 271690 3544 271696 3556
rect 271748 3544 271754 3596
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 365714 3544 365720 3596
rect 365772 3584 365778 3596
rect 366910 3584 366916 3596
rect 365772 3556 366916 3584
rect 365772 3544 365778 3556
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 373994 3544 374000 3596
rect 374052 3584 374058 3596
rect 375190 3584 375196 3596
rect 374052 3556 375196 3584
rect 374052 3544 374058 3556
rect 375190 3544 375196 3556
rect 375248 3544 375254 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 482278 3584 482284 3596
rect 380860 3556 482284 3584
rect 380860 3544 380866 3556
rect 482278 3544 482284 3556
rect 482336 3544 482342 3596
rect 485774 3544 485780 3596
rect 485832 3584 485838 3596
rect 486970 3584 486976 3596
rect 485832 3556 486976 3584
rect 485832 3544 485838 3556
rect 486970 3544 486976 3556
rect 487028 3544 487034 3596
rect 494146 3544 494152 3596
rect 494204 3584 494210 3596
rect 495342 3584 495348 3596
rect 494204 3556 495348 3584
rect 494204 3544 494210 3556
rect 495342 3544 495348 3556
rect 495400 3544 495406 3596
rect 520274 3544 520280 3596
rect 520332 3584 520338 3596
rect 521470 3584 521476 3596
rect 520332 3556 521476 3584
rect 520332 3544 520338 3556
rect 521470 3544 521476 3556
rect 521528 3544 521534 3596
rect 528554 3544 528560 3596
rect 528612 3584 528618 3596
rect 529842 3584 529848 3596
rect 528612 3556 529848 3584
rect 528612 3544 528618 3556
rect 529842 3544 529848 3556
rect 529900 3544 529906 3596
rect 536926 3544 536932 3596
rect 536984 3584 536990 3596
rect 538122 3584 538128 3596
rect 536984 3556 538128 3584
rect 536984 3544 536990 3556
rect 538122 3544 538128 3556
rect 538180 3544 538186 3596
rect 546494 3544 546500 3596
rect 546552 3584 546558 3596
rect 547690 3584 547696 3596
rect 546552 3556 547696 3584
rect 546552 3544 546558 3556
rect 547690 3544 547696 3556
rect 547748 3544 547754 3596
rect 573358 3544 573364 3596
rect 573416 3584 573422 3596
rect 575014 3584 575020 3596
rect 573416 3556 575020 3584
rect 573416 3544 573422 3556
rect 575014 3544 575020 3556
rect 575072 3544 575078 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 131114 3516 131120 3528
rect 624 3488 131120 3516
rect 624 3476 630 3488
rect 131114 3476 131120 3488
rect 131172 3476 131178 3528
rect 137278 3476 137284 3528
rect 137336 3516 137342 3528
rect 140774 3516 140780 3528
rect 137336 3488 140780 3516
rect 137336 3476 137342 3488
rect 140774 3476 140780 3488
rect 140832 3476 140838 3528
rect 145650 3476 145656 3528
rect 145708 3516 145714 3528
rect 146294 3516 146300 3528
rect 145708 3488 146300 3516
rect 145708 3476 145714 3488
rect 146294 3476 146300 3488
rect 146352 3476 146358 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151538 3516 151544 3528
rect 150676 3488 151544 3516
rect 150676 3476 150682 3488
rect 151538 3476 151544 3488
rect 151596 3476 151602 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 152734 3516 152740 3528
rect 151872 3488 152740 3516
rect 151872 3476 151878 3488
rect 152734 3476 152740 3488
rect 152792 3476 152798 3528
rect 153102 3476 153108 3528
rect 153160 3516 153166 3528
rect 153930 3516 153936 3528
rect 153160 3488 153936 3516
rect 153160 3476 153166 3488
rect 153930 3476 153936 3488
rect 153988 3476 153994 3528
rect 155770 3476 155776 3528
rect 155828 3516 155834 3528
rect 156322 3516 156328 3528
rect 155828 3488 156328 3516
rect 155828 3476 155834 3488
rect 156322 3476 156328 3488
rect 156380 3476 156386 3528
rect 157242 3476 157248 3528
rect 157300 3516 157306 3528
rect 158714 3516 158720 3528
rect 157300 3488 158720 3516
rect 157300 3476 157306 3488
rect 158714 3476 158720 3488
rect 158772 3476 158778 3528
rect 165522 3476 165528 3528
rect 165580 3516 165586 3528
rect 170582 3516 170588 3528
rect 165580 3488 170588 3516
rect 165580 3476 165586 3488
rect 170582 3476 170588 3488
rect 170640 3476 170646 3528
rect 171042 3476 171048 3528
rect 171100 3516 171106 3528
rect 178954 3516 178960 3528
rect 171100 3488 178960 3516
rect 171100 3476 171106 3488
rect 178954 3476 178960 3488
rect 179012 3476 179018 3528
rect 179322 3476 179328 3528
rect 179380 3516 179386 3528
rect 192018 3516 192024 3528
rect 179380 3488 192024 3516
rect 179380 3476 179386 3488
rect 192018 3476 192024 3488
rect 192076 3476 192082 3528
rect 193122 3476 193128 3528
rect 193180 3516 193186 3528
rect 211062 3516 211068 3528
rect 193180 3488 211068 3516
rect 193180 3476 193186 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 235994 3516 236000 3528
rect 211172 3488 236000 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 132494 3448 132500 3460
rect 1728 3420 132500 3448
rect 1728 3408 1734 3420
rect 132494 3408 132500 3420
rect 132552 3408 132558 3460
rect 134886 3408 134892 3460
rect 134944 3448 134950 3460
rect 139486 3448 139492 3460
rect 134944 3420 139492 3448
rect 134944 3408 134950 3420
rect 139486 3408 139492 3420
rect 139544 3408 139550 3460
rect 144454 3408 144460 3460
rect 144512 3448 144518 3460
rect 146386 3448 146392 3460
rect 144512 3420 146392 3448
rect 144512 3408 144518 3420
rect 146386 3408 146392 3420
rect 146444 3408 146450 3460
rect 154482 3408 154488 3460
rect 154540 3448 154546 3460
rect 155126 3448 155132 3460
rect 154540 3420 155132 3448
rect 154540 3408 154546 3420
rect 155126 3408 155132 3420
rect 155184 3408 155190 3460
rect 158622 3408 158628 3460
rect 158680 3448 158686 3460
rect 161106 3448 161112 3460
rect 158680 3420 161112 3448
rect 158680 3408 158686 3420
rect 161106 3408 161112 3420
rect 161164 3408 161170 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 165890 3448 165896 3460
rect 161348 3420 165896 3448
rect 161348 3408 161354 3420
rect 165890 3408 165896 3420
rect 165948 3408 165954 3460
rect 168282 3408 168288 3460
rect 168340 3448 168346 3460
rect 175366 3448 175372 3460
rect 168340 3420 175372 3448
rect 168340 3408 168346 3420
rect 175366 3408 175372 3420
rect 175424 3408 175430 3460
rect 177942 3408 177948 3460
rect 178000 3448 178006 3460
rect 189626 3448 189632 3460
rect 178000 3420 189632 3448
rect 178000 3408 178006 3420
rect 189626 3408 189632 3420
rect 189684 3408 189690 3460
rect 190362 3408 190368 3460
rect 190420 3448 190426 3460
rect 207474 3448 207480 3460
rect 190420 3420 207480 3448
rect 190420 3408 190426 3420
rect 207474 3408 207480 3420
rect 207532 3408 207538 3460
rect 210970 3408 210976 3460
rect 211028 3448 211034 3460
rect 211172 3448 211200 3488
rect 235994 3476 236000 3488
rect 236052 3476 236058 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 252554 3476 252560 3528
rect 252612 3516 252618 3528
rect 253842 3516 253848 3528
rect 252612 3488 253848 3516
rect 252612 3476 252618 3488
rect 253842 3476 253848 3488
rect 253900 3476 253906 3528
rect 287054 3476 287060 3528
rect 287112 3516 287118 3528
rect 288342 3516 288348 3528
rect 287112 3488 288348 3516
rect 287112 3476 287118 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 296714 3476 296720 3528
rect 296772 3516 296778 3528
rect 297910 3516 297916 3528
rect 296772 3488 297916 3516
rect 296772 3476 296778 3488
rect 297910 3476 297916 3488
rect 297968 3476 297974 3528
rect 304994 3476 305000 3528
rect 305052 3516 305058 3528
rect 306190 3516 306196 3528
rect 305052 3488 306196 3516
rect 305052 3476 305058 3488
rect 306190 3476 306196 3488
rect 306248 3476 306254 3528
rect 313366 3476 313372 3528
rect 313424 3516 313430 3528
rect 314562 3516 314568 3528
rect 313424 3488 314568 3516
rect 313424 3476 313430 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 347774 3476 347780 3528
rect 347832 3516 347838 3528
rect 349062 3516 349068 3528
rect 347832 3488 349068 3516
rect 347832 3476 347838 3488
rect 349062 3476 349068 3488
rect 349120 3476 349126 3528
rect 356054 3476 356060 3528
rect 356112 3516 356118 3528
rect 357342 3516 357348 3528
rect 356112 3488 357348 3516
rect 356112 3476 356118 3488
rect 357342 3476 357348 3488
rect 357400 3476 357406 3528
rect 358722 3476 358728 3528
rect 358780 3516 358786 3528
rect 450170 3516 450176 3528
rect 358780 3488 450176 3516
rect 358780 3476 358786 3488
rect 450170 3476 450176 3488
rect 450228 3476 450234 3528
rect 451182 3476 451188 3528
rect 451240 3516 451246 3528
rect 582190 3516 582196 3528
rect 451240 3488 582196 3516
rect 451240 3476 451246 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 211028 3420 211200 3448
rect 211028 3408 211034 3420
rect 212442 3408 212448 3460
rect 212500 3448 212506 3460
rect 239582 3448 239588 3460
rect 212500 3420 239588 3448
rect 212500 3408 212506 3420
rect 239582 3408 239588 3420
rect 239640 3408 239646 3460
rect 355962 3408 355968 3460
rect 356020 3448 356026 3460
rect 446582 3448 446588 3460
rect 356020 3420 446588 3448
rect 356020 3408 356026 3420
rect 446582 3408 446588 3420
rect 446640 3408 446646 3460
rect 448422 3408 448428 3460
rect 448480 3448 448486 3460
rect 578602 3448 578608 3460
rect 448480 3420 578608 3448
rect 448480 3408 448486 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 164050 3340 164056 3392
rect 164108 3380 164114 3392
rect 169386 3380 169392 3392
rect 164108 3352 169392 3380
rect 164108 3340 164114 3352
rect 169386 3340 169392 3352
rect 169444 3340 169450 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 416774 3340 416780 3392
rect 416832 3380 416838 3392
rect 417970 3380 417976 3392
rect 416832 3352 417976 3380
rect 416832 3340 416838 3352
rect 417970 3340 417976 3352
rect 418028 3340 418034 3392
rect 433334 3340 433340 3392
rect 433392 3380 433398 3392
rect 434622 3380 434628 3392
rect 433392 3352 434628 3380
rect 433392 3340 433398 3352
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 133782 3272 133788 3324
rect 133840 3312 133846 3324
rect 138014 3312 138020 3324
rect 133840 3284 138020 3312
rect 133840 3272 133846 3284
rect 138014 3272 138020 3284
rect 138072 3272 138078 3324
rect 155862 3272 155868 3324
rect 155920 3312 155926 3324
rect 157518 3312 157524 3324
rect 155920 3284 157524 3312
rect 155920 3272 155926 3284
rect 157518 3272 157524 3284
rect 157576 3272 157582 3324
rect 162762 3272 162768 3324
rect 162820 3312 162826 3324
rect 167086 3312 167092 3324
rect 162820 3284 167092 3312
rect 162820 3272 162826 3284
rect 167086 3272 167092 3284
rect 167144 3272 167150 3324
rect 172330 3272 172336 3324
rect 172388 3312 172394 3324
rect 180150 3312 180156 3324
rect 172388 3284 180156 3312
rect 172388 3272 172394 3284
rect 180150 3272 180156 3284
rect 180208 3272 180214 3324
rect 136082 3204 136088 3256
rect 136140 3244 136146 3256
rect 139394 3244 139400 3256
rect 136140 3216 139400 3244
rect 136140 3204 136146 3216
rect 139394 3204 139400 3216
rect 139452 3204 139458 3256
rect 164142 3204 164148 3256
rect 164200 3244 164206 3256
rect 168190 3244 168196 3256
rect 164200 3216 168196 3244
rect 164200 3204 164206 3216
rect 168190 3204 168196 3216
rect 168248 3204 168254 3256
rect 132586 3136 132592 3188
rect 132644 3176 132650 3188
rect 138106 3176 138112 3188
rect 132644 3148 138112 3176
rect 132644 3136 132650 3148
rect 138106 3136 138112 3148
rect 138164 3136 138170 3188
rect 131390 3068 131396 3120
rect 131448 3108 131454 3120
rect 136634 3108 136640 3120
rect 131448 3080 136640 3108
rect 131448 3068 131454 3080
rect 136634 3068 136640 3080
rect 136692 3068 136698 3120
rect 213089 3111 213147 3117
rect 213089 3077 213101 3111
rect 213135 3108 213147 3111
rect 221734 3108 221740 3120
rect 213135 3080 221740 3108
rect 213135 3077 213147 3080
rect 213089 3071 213147 3077
rect 221734 3068 221740 3080
rect 221792 3068 221798 3120
rect 157150 3000 157156 3052
rect 157208 3040 157214 3052
rect 159910 3040 159916 3052
rect 157208 3012 159916 3040
rect 157208 3000 157214 3012
rect 159910 3000 159916 3012
rect 159968 3000 159974 3052
rect 143258 2864 143264 2916
rect 143316 2904 143322 2916
rect 144914 2904 144920 2916
rect 143316 2876 144920 2904
rect 143316 2864 143322 2876
rect 144914 2864 144920 2876
rect 144972 2864 144978 2916
rect 165430 2864 165436 2916
rect 165488 2904 165494 2916
rect 171778 2904 171784 2916
rect 165488 2876 171784 2904
rect 165488 2864 165494 2876
rect 171778 2864 171784 2876
rect 171836 2864 171842 2916
rect 502334 2728 502340 2780
rect 502392 2768 502398 2780
rect 503622 2768 503628 2780
rect 502392 2740 503628 2768
rect 502392 2728 502398 2740
rect 503622 2728 503628 2740
rect 503680 2728 503686 2780
rect 563054 2728 563060 2780
rect 563112 2768 563118 2780
rect 564342 2768 564348 2780
rect 563112 2740 564348 2768
rect 563112 2728 563118 2740
rect 564342 2728 564348 2740
rect 564400 2728 564406 2780
rect 571334 2728 571340 2780
rect 571392 2768 571398 2780
rect 572622 2768 572628 2780
rect 571392 2740 572628 2768
rect 571392 2728 571398 2740
rect 572622 2728 572628 2740
rect 572680 2728 572686 2780
rect 364334 552 364340 604
rect 364392 592 364398 604
rect 364518 592 364524 604
rect 364392 564 364524 592
rect 364392 552 364398 564
rect 364518 552 364524 564
rect 364576 552 364582 604
rect 367094 552 367100 604
rect 367152 592 367158 604
rect 368014 592 368020 604
rect 367152 564 368020 592
rect 367152 552 367158 564
rect 368014 552 368020 564
rect 368072 552 368078 604
rect 368474 552 368480 604
rect 368532 592 368538 604
rect 369210 592 369216 604
rect 368532 564 369216 592
rect 368532 552 368538 564
rect 369210 552 369216 564
rect 369268 552 369274 604
rect 369854 552 369860 604
rect 369912 592 369918 604
rect 370406 592 370412 604
rect 369912 564 370412 592
rect 369912 552 369918 564
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 372614 552 372620 604
rect 372672 592 372678 604
rect 372798 592 372804 604
rect 372672 564 372804 592
rect 372672 552 372678 564
rect 372798 552 372804 564
rect 372856 552 372862 604
<< via1 >>
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 413008 698232 413060 698284
rect 413744 698232 413796 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 331220 697552 331272 697604
rect 332508 697552 332560 697604
rect 472624 696940 472676 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 694084 72752 694136
rect 412824 694084 412876 694136
rect 413008 694084 413060 694136
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 347780 692792 347832 692844
rect 348884 692792 348936 692844
rect 364340 692792 364392 692844
rect 365076 692792 365128 692844
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 412824 692724 412876 692776
rect 542544 692724 542596 692776
rect 542728 692724 542780 692776
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 494244 685856 494296 685908
rect 494888 685856 494940 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 429200 684428 429252 684480
rect 429844 684428 429896 684480
rect 558920 684428 558972 684480
rect 559656 684428 559708 684480
rect 412640 683247 412692 683256
rect 412640 683213 412649 683247
rect 412649 683213 412683 683247
rect 412683 683213 412692 683247
rect 412640 683204 412692 683213
rect 412640 683068 412692 683120
rect 429200 683068 429252 683120
rect 542360 683068 542412 683120
rect 558920 683068 558972 683120
rect 3516 681708 3568 681760
rect 8944 681708 8996 681760
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 347780 673480 347832 673532
rect 347964 673480 348016 673532
rect 364340 673480 364392 673532
rect 364524 673480 364576 673532
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 490564 673480 490616 673532
rect 580172 673480 580224 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 3424 667904 3476 667956
rect 17224 667904 17276 667956
rect 219072 666544 219124 666596
rect 413100 666544 413152 666596
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 73068 656820 73120 656872
rect 219348 656820 219400 656872
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 284024 654100 284076 654152
rect 284208 654100 284260 654152
rect 347780 654100 347832 654152
rect 347964 654100 348016 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 14464 652740 14516 652792
rect 471244 650020 471296 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 412824 647232 412876 647284
rect 412916 647232 412968 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 72976 640364 73028 640416
rect 219256 640364 219308 640416
rect 412824 640364 412876 640416
rect 412916 640364 412968 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 72792 640228 72844 640280
rect 219072 640228 219124 640280
rect 72792 637508 72844 637560
rect 72884 637508 72936 637560
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 137744 634788 137796 634840
rect 137928 634788 137980 634840
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 284024 634788 284076 634840
rect 284208 634788 284260 634840
rect 347780 634788 347832 634840
rect 347964 634788 348016 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 412732 630640 412784 630692
rect 412916 630640 412968 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 479524 626560 479576 626612
rect 580172 626560 580224 626612
rect 73068 626535 73120 626544
rect 73068 626501 73077 626535
rect 73077 626501 73111 626535
rect 73111 626501 73120 626535
rect 73068 626492 73120 626501
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 3424 623772 3476 623824
rect 10324 623772 10376 623824
rect 73068 616879 73120 616888
rect 73068 616845 73077 616879
rect 73077 616845 73111 616879
rect 73111 616845 73120 616879
rect 73068 616836 73120 616845
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 137744 615476 137796 615528
rect 137928 615476 137980 615528
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 284024 615476 284076 615528
rect 284208 615476 284260 615528
rect 347780 615476 347832 615528
rect 347964 615476 348016 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 477500 615476 477552 615528
rect 477684 615476 477736 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 73068 611396 73120 611448
rect 219348 611396 219400 611448
rect 412732 611328 412784 611380
rect 412916 611328 412968 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 72884 611260 72936 611312
rect 3424 609968 3476 610020
rect 19984 609968 20036 610020
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 412824 608583 412876 608592
rect 412824 608549 412833 608583
rect 412833 608549 412867 608583
rect 412867 608549 412876 608583
rect 412824 608540 412876 608549
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 542544 608583 542596 608592
rect 542544 608549 542553 608583
rect 542553 608549 542587 608583
rect 542587 608549 542596 608583
rect 542544 608540 542596 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 467104 603100 467156 603152
rect 580172 603100 580224 603152
rect 413008 601672 413060 601724
rect 429568 601672 429620 601724
rect 542728 601672 542780 601724
rect 559288 601672 559340 601724
rect 72976 601536 73028 601588
rect 73160 601536 73212 601588
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 72976 598884 73028 598936
rect 219256 598884 219308 598936
rect 413008 598927 413060 598936
rect 413008 598893 413017 598927
rect 413017 598893 413051 598927
rect 413051 598893 413060 598927
rect 413008 598884 413060 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 542728 598927 542780 598936
rect 542728 598893 542737 598927
rect 542737 598893 542771 598927
rect 542771 598893 542780 598927
rect 542728 598884 542780 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 137744 596164 137796 596216
rect 137928 596164 137980 596216
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 284024 596164 284076 596216
rect 284208 596164 284260 596216
rect 347780 596164 347832 596216
rect 347964 596164 348016 596216
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 477500 596164 477552 596216
rect 477684 596164 477736 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 13084 594804 13136 594856
rect 476764 592016 476816 592068
rect 579896 592016 579948 592068
rect 72884 589339 72936 589348
rect 72884 589305 72893 589339
rect 72893 589305 72927 589339
rect 72927 589305 72936 589339
rect 72884 589296 72936 589305
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 413100 589296 413152 589348
rect 429660 589296 429712 589348
rect 542820 589296 542872 589348
rect 559380 589296 559432 589348
rect 8024 589271 8076 589280
rect 8024 589237 8033 589271
rect 8033 589237 8067 589271
rect 8067 589237 8076 589271
rect 8024 589228 8076 589237
rect 137744 589271 137796 589280
rect 137744 589237 137753 589271
rect 137753 589237 137787 589271
rect 137787 589237 137796 589271
rect 137744 589228 137796 589237
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 284024 589271 284076 589280
rect 284024 589237 284033 589271
rect 284033 589237 284067 589271
rect 284067 589237 284076 589271
rect 284024 589228 284076 589237
rect 347872 589228 347924 589280
rect 364432 589228 364484 589280
rect 477592 589228 477644 589280
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 72700 582360 72752 582412
rect 72884 582360 72936 582412
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 413100 582428 413152 582480
rect 429660 582428 429712 582480
rect 542820 582428 542872 582480
rect 559380 582428 559432 582480
rect 413008 582292 413060 582344
rect 429568 582292 429620 582344
rect 542728 582292 542780 582344
rect 559288 582292 559340 582344
rect 8024 579751 8076 579760
rect 8024 579717 8033 579751
rect 8033 579717 8067 579751
rect 8067 579717 8076 579751
rect 8024 579708 8076 579717
rect 137744 579751 137796 579760
rect 137744 579717 137753 579751
rect 137753 579717 137787 579751
rect 137787 579717 137796 579751
rect 137744 579708 137796 579717
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 284024 579751 284076 579760
rect 284024 579717 284033 579751
rect 284033 579717 284067 579751
rect 284067 579717 284076 579751
rect 284024 579708 284076 579717
rect 347780 579683 347832 579692
rect 347780 579649 347789 579683
rect 347789 579649 347823 579683
rect 347823 579649 347832 579683
rect 364340 579683 364392 579692
rect 347780 579640 347832 579649
rect 364340 579649 364349 579683
rect 364349 579649 364383 579683
rect 364383 579649 364392 579683
rect 364340 579640 364392 579649
rect 477500 579683 477552 579692
rect 477500 579649 477509 579683
rect 477509 579649 477543 579683
rect 477543 579649 477552 579683
rect 477500 579640 477552 579649
rect 489184 579640 489236 579692
rect 580172 579640 580224 579692
rect 7932 579572 7984 579624
rect 8116 579572 8168 579624
rect 72700 579572 72752 579624
rect 137652 579572 137704 579624
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 283932 579572 283984 579624
rect 284116 579572 284168 579624
rect 72608 569959 72660 569968
rect 72608 569925 72617 569959
rect 72617 569925 72651 569959
rect 72651 569925 72660 569959
rect 72608 569916 72660 569925
rect 137560 569959 137612 569968
rect 137560 569925 137569 569959
rect 137569 569925 137603 569959
rect 137603 569925 137612 569959
rect 137560 569916 137612 569925
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 347872 569891 347924 569900
rect 347872 569857 347881 569891
rect 347881 569857 347915 569891
rect 347915 569857 347924 569891
rect 347872 569848 347924 569857
rect 364432 569891 364484 569900
rect 364432 569857 364441 569891
rect 364441 569857 364475 569891
rect 364475 569857 364484 569891
rect 364432 569848 364484 569857
rect 477592 569891 477644 569900
rect 477592 569857 477601 569891
rect 477601 569857 477635 569891
rect 477635 569857 477644 569891
rect 477592 569848 477644 569857
rect 494152 569891 494204 569900
rect 494152 569857 494161 569891
rect 494161 569857 494195 569891
rect 494195 569857 494204 569891
rect 494152 569848 494204 569857
rect 13084 567808 13136 567860
rect 129004 567808 129056 567860
rect 4068 567264 4120 567316
rect 11704 567264 11756 567316
rect 412732 563116 412784 563168
rect 429292 563116 429344 563168
rect 542452 563116 542504 563168
rect 559012 563116 559064 563168
rect 72608 563048 72660 563100
rect 137560 563048 137612 563100
rect 218888 563048 218940 563100
rect 348056 563048 348108 563100
rect 364616 563048 364668 563100
rect 7932 562912 7984 562964
rect 8116 562912 8168 562964
rect 72700 562912 72752 562964
rect 137652 562912 137704 562964
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 477776 563048 477828 563100
rect 494336 563048 494388 563100
rect 412732 562980 412784 563032
rect 429292 562980 429344 563032
rect 542452 562980 542504 563032
rect 559012 562980 559064 563032
rect 218980 562912 219032 562964
rect 283932 562912 283984 562964
rect 284116 562912 284168 562964
rect 72700 560235 72752 560244
rect 72700 560201 72709 560235
rect 72709 560201 72743 560235
rect 72743 560201 72752 560235
rect 72700 560192 72752 560201
rect 137652 560235 137704 560244
rect 137652 560201 137661 560235
rect 137661 560201 137695 560235
rect 137695 560201 137704 560235
rect 137652 560192 137704 560201
rect 218980 560235 219032 560244
rect 218980 560201 218989 560235
rect 218989 560201 219023 560235
rect 219023 560201 219032 560235
rect 218980 560192 219032 560201
rect 412732 560235 412784 560244
rect 412732 560201 412741 560235
rect 412741 560201 412775 560235
rect 412775 560201 412784 560235
rect 412732 560192 412784 560201
rect 429292 560235 429344 560244
rect 429292 560201 429301 560235
rect 429301 560201 429335 560235
rect 429335 560201 429344 560235
rect 429292 560192 429344 560201
rect 542452 560235 542504 560244
rect 542452 560201 542461 560235
rect 542461 560201 542495 560235
rect 542495 560201 542504 560235
rect 542452 560192 542504 560201
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 483664 556180 483716 556232
rect 580172 556180 580224 556232
rect 72884 550604 72936 550656
rect 137836 550604 137888 550656
rect 219164 550604 219216 550656
rect 347872 550604 347924 550656
rect 348148 550604 348200 550656
rect 364432 550604 364484 550656
rect 364708 550604 364760 550656
rect 412916 550604 412968 550656
rect 429476 550604 429528 550656
rect 477592 550604 477644 550656
rect 477868 550604 477920 550656
rect 494152 550604 494204 550656
rect 494428 550604 494480 550656
rect 542636 550604 542688 550656
rect 559196 550604 559248 550656
rect 8024 550579 8076 550588
rect 8024 550545 8033 550579
rect 8033 550545 8067 550579
rect 8067 550545 8076 550579
rect 8024 550536 8076 550545
rect 154304 550579 154356 550588
rect 154304 550545 154313 550579
rect 154313 550545 154347 550579
rect 154347 550545 154356 550579
rect 154304 550536 154356 550545
rect 284024 550579 284076 550588
rect 284024 550545 284033 550579
rect 284033 550545 284067 550579
rect 284067 550545 284076 550579
rect 284024 550536 284076 550545
rect 475384 545096 475436 545148
rect 579896 545096 579948 545148
rect 8208 543736 8260 543788
rect 154488 543736 154540 543788
rect 284208 543736 284260 543788
rect 348148 543804 348200 543856
rect 364708 543804 364760 543856
rect 477868 543804 477920 543856
rect 494428 543804 494480 543856
rect 348056 543668 348108 543720
rect 364616 543668 364668 543720
rect 477776 543668 477828 543720
rect 494336 543668 494388 543720
rect 72700 543600 72752 543652
rect 72884 543600 72936 543652
rect 137652 543600 137704 543652
rect 137836 543600 137888 543652
rect 218980 543600 219032 543652
rect 219164 543600 219216 543652
rect 412732 543600 412784 543652
rect 412916 543600 412968 543652
rect 429292 543600 429344 543652
rect 429476 543600 429528 543652
rect 542452 543600 542504 543652
rect 542636 543600 542688 543652
rect 559012 543600 559064 543652
rect 559196 543600 559248 543652
rect 3700 538228 3752 538280
rect 15844 538228 15896 538280
rect 72700 534012 72752 534064
rect 72884 534012 72936 534064
rect 137652 534012 137704 534064
rect 137836 534012 137888 534064
rect 218980 534012 219032 534064
rect 219164 534012 219216 534064
rect 485044 532720 485096 532772
rect 580172 532720 580224 532772
rect 7932 531292 7984 531344
rect 8024 531292 8076 531344
rect 154212 531292 154264 531344
rect 154304 531292 154356 531344
rect 347872 531292 347924 531344
rect 348148 531292 348200 531344
rect 364432 531292 364484 531344
rect 364708 531292 364760 531344
rect 477592 531292 477644 531344
rect 477868 531292 477920 531344
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 72792 524467 72844 524476
rect 72792 524433 72801 524467
rect 72801 524433 72835 524467
rect 72835 524433 72844 524467
rect 72792 524424 72844 524433
rect 137744 524467 137796 524476
rect 137744 524433 137753 524467
rect 137753 524433 137787 524467
rect 137787 524433 137796 524467
rect 137744 524424 137796 524433
rect 154304 524424 154356 524476
rect 219072 524467 219124 524476
rect 219072 524433 219081 524467
rect 219081 524433 219115 524467
rect 219115 524433 219124 524467
rect 219072 524424 219124 524433
rect 8116 524288 8168 524340
rect 8300 524288 8352 524340
rect 154396 524288 154448 524340
rect 284116 524288 284168 524340
rect 284300 524288 284352 524340
rect 72792 521679 72844 521688
rect 72792 521645 72801 521679
rect 72801 521645 72835 521679
rect 72835 521645 72844 521679
rect 72792 521636 72844 521645
rect 137744 521679 137796 521688
rect 137744 521645 137753 521679
rect 137753 521645 137787 521679
rect 137787 521645 137796 521679
rect 137744 521636 137796 521645
rect 219072 521679 219124 521688
rect 219072 521645 219081 521679
rect 219081 521645 219115 521679
rect 219115 521645 219124 521679
rect 219072 521636 219124 521645
rect 347964 521636 348016 521688
rect 348148 521636 348200 521688
rect 364524 521636 364576 521688
rect 364708 521636 364760 521688
rect 477684 521636 477736 521688
rect 477868 521636 477920 521688
rect 494244 521636 494296 521688
rect 494428 521636 494480 521688
rect 284116 516060 284168 516112
rect 291108 516060 291160 516112
rect 106188 515720 106240 515772
rect 196808 515720 196860 515772
rect 385500 515720 385552 515772
rect 462320 515720 462372 515772
rect 89628 515652 89680 515704
rect 185032 515652 185084 515704
rect 397276 515652 397328 515704
rect 477684 515652 477736 515704
rect 72792 515584 72844 515636
rect 173256 515584 173308 515636
rect 202788 515584 202840 515636
rect 244004 515584 244056 515636
rect 409052 515584 409104 515636
rect 494244 515584 494296 515636
rect 41328 515516 41380 515568
rect 161480 515516 161532 515568
rect 171048 515516 171100 515568
rect 232228 515516 232280 515568
rect 350080 515516 350132 515568
rect 397460 515516 397512 515568
rect 420828 515516 420880 515568
rect 527180 515516 527232 515568
rect 24768 515448 24820 515500
rect 149704 515448 149756 515500
rect 154396 515448 154448 515500
rect 220452 515448 220504 515500
rect 235908 515448 235960 515500
rect 267556 515448 267608 515500
rect 326528 515448 326580 515500
rect 347964 515448 348016 515500
rect 361856 515448 361908 515500
rect 412916 515448 412968 515500
rect 432604 515448 432656 515500
rect 542636 515448 542688 515500
rect 8116 515380 8168 515432
rect 137928 515380 137980 515432
rect 138020 515380 138072 515432
rect 208584 515380 208636 515432
rect 219072 515380 219124 515432
rect 255780 515380 255832 515432
rect 267648 515380 267700 515432
rect 279332 515380 279384 515432
rect 314752 515380 314804 515432
rect 331220 515380 331272 515432
rect 338304 515380 338356 515432
rect 364524 515380 364576 515432
rect 373632 515380 373684 515432
rect 429476 515380 429528 515432
rect 444380 515380 444432 515432
rect 559196 515380 559248 515432
rect 300768 514836 300820 514888
rect 302976 514836 303028 514888
rect 2872 509260 2924 509312
rect 13084 509260 13136 509312
rect 462964 509260 463016 509312
rect 580172 509260 580224 509312
rect 8944 509192 8996 509244
rect 128360 509192 128412 509244
rect 453212 509192 453264 509244
rect 472624 509192 472676 509244
rect 17224 502256 17276 502308
rect 128360 502256 128412 502308
rect 453396 502256 453448 502308
rect 580264 502256 580316 502308
rect 460204 498176 460256 498228
rect 580172 498176 580224 498228
rect 453948 495388 454000 495440
rect 490564 495388 490616 495440
rect 14464 493960 14516 494012
rect 128360 493960 128412 494012
rect 453764 488452 453816 488504
rect 471244 488452 471296 488504
rect 456064 485800 456116 485852
rect 580172 485800 580224 485852
rect 10324 485732 10376 485784
rect 128360 485732 128412 485784
rect 453764 481584 453816 481636
rect 580356 481584 580408 481636
rect 3332 480224 3384 480276
rect 8944 480224 8996 480276
rect 19984 478796 20036 478848
rect 128360 478796 128412 478848
rect 453948 473288 454000 473340
rect 479524 473288 479576 473340
rect 452752 466352 452804 466404
rect 467104 466352 467156 466404
rect 11704 463632 11756 463684
rect 128360 463632 128412 463684
rect 454684 462340 454736 462392
rect 580172 462340 580224 462392
rect 453396 459484 453448 459536
rect 476764 459484 476816 459536
rect 3424 455336 3476 455388
rect 128360 455336 128412 455388
rect 453948 452548 454000 452600
rect 489184 452548 489236 452600
rect 3148 451256 3200 451308
rect 58624 451256 58676 451308
rect 15844 448468 15896 448520
rect 128360 448468 128412 448520
rect 453672 445680 453724 445732
rect 483664 445680 483716 445732
rect 13084 440172 13136 440224
rect 128360 440172 128412 440224
rect 453304 438880 453356 438932
rect 579896 438880 579948 438932
rect 453764 438812 453816 438864
rect 475384 438812 475436 438864
rect 3516 433236 3568 433288
rect 128360 433236 128412 433288
rect 453948 430516 454000 430568
rect 485044 430516 485096 430568
rect 8944 425008 8996 425060
rect 128360 425008 128412 425060
rect 453948 423580 454000 423632
rect 462964 423580 463016 423632
rect 58624 418072 58676 418124
rect 128360 418072 128412 418124
rect 453948 416372 454000 416424
rect 460204 416372 460256 416424
rect 543004 414672 543056 414724
rect 580172 414672 580224 414724
rect 3424 409776 3476 409828
rect 128360 409776 128412 409828
rect 453396 409368 453448 409420
rect 456064 409368 456116 409420
rect 3516 402908 3568 402960
rect 128360 402908 128412 402960
rect 452844 402500 452896 402552
rect 454684 402500 454736 402552
rect 453764 395972 453816 396024
rect 580264 395972 580316 396024
rect 3424 394612 3476 394664
rect 128360 394612 128412 394664
rect 454684 391960 454736 392012
rect 580172 391960 580224 392012
rect 3240 380808 3292 380860
rect 129004 380808 129056 380860
rect 453948 380808 454000 380860
rect 543004 380808 543056 380860
rect 453396 373940 453448 373992
rect 580356 373940 580408 373992
rect 3148 367004 3200 367056
rect 129004 367004 129056 367056
rect 452660 367004 452712 367056
rect 454684 367004 454736 367056
rect 453948 360136 454000 360188
rect 580264 360136 580316 360188
rect 453764 353200 453816 353252
rect 580264 353200 580316 353252
rect 8944 347760 8996 347812
rect 128360 347760 128412 347812
rect 453948 345652 454000 345704
rect 580172 345652 580224 345704
rect 3424 338036 3476 338088
rect 129280 338036 129332 338088
rect 13084 332596 13136 332648
rect 128360 332596 128412 332648
rect 11704 324300 11756 324352
rect 128360 324300 128412 324352
rect 3240 324232 3292 324284
rect 129004 324232 129056 324284
rect 453488 322872 453540 322924
rect 580172 322872 580224 322924
rect 453396 311788 453448 311840
rect 580172 311788 580224 311840
rect 15844 309136 15896 309188
rect 128360 309136 128412 309188
rect 3332 309068 3384 309120
rect 129188 309068 129240 309120
rect 452936 302336 452988 302388
rect 454684 302336 454736 302388
rect 10324 302200 10376 302252
rect 128360 302200 128412 302252
rect 453304 299412 453356 299464
rect 579804 299412 579856 299464
rect 3516 294856 3568 294908
rect 8944 294856 8996 294908
rect 17224 287036 17276 287088
rect 128360 287036 128412 287088
rect 453028 280168 453080 280220
rect 456064 280168 456116 280220
rect 3424 280100 3476 280152
rect 129096 280100 129148 280152
rect 126244 278740 126296 278792
rect 129096 278740 129148 278792
rect 453580 275952 453632 276004
rect 580172 275952 580224 276004
rect 3148 266296 3200 266348
rect 13084 266296 13136 266348
rect 453488 264868 453540 264920
rect 580172 264868 580224 264920
rect 13084 263576 13136 263628
rect 128360 263576 128412 263628
rect 453948 259428 454000 259480
rect 471244 259428 471296 259480
rect 14464 256708 14516 256760
rect 128360 256708 128412 256760
rect 3424 252492 3476 252544
rect 11704 252492 11756 252544
rect 454684 252492 454736 252544
rect 579804 252492 579856 252544
rect 452844 250452 452896 250504
rect 479524 250452 479576 250504
rect 19984 241476 20036 241528
rect 128360 241476 128412 241528
rect 453948 237396 454000 237448
rect 469864 237396 469916 237448
rect 3424 237328 3476 237380
rect 129004 237328 129056 237380
rect 8944 233248 8996 233300
rect 128360 233248 128412 233300
rect 453120 230460 453172 230512
rect 472624 230460 472676 230512
rect 453396 229032 453448 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 15844 223524 15896 223576
rect 15844 218016 15896 218068
rect 128360 218016 128412 218068
rect 453304 217948 453356 218000
rect 580172 217948 580224 218000
rect 452936 216792 452988 216844
rect 454684 216792 454736 216844
rect 11704 211148 11756 211200
rect 128360 211148 128412 211200
rect 453948 209788 454000 209840
rect 478144 209788 478196 209840
rect 3424 208292 3476 208344
rect 10324 208292 10376 208344
rect 456064 205572 456116 205624
rect 579804 205572 579856 205624
rect 10324 194556 10376 194608
rect 128636 194556 128688 194608
rect 453948 194556 454000 194608
rect 483664 194556 483716 194608
rect 3148 194488 3200 194540
rect 129372 194488 129424 194540
rect 295616 190340 295668 190392
rect 296536 190340 296588 190392
rect 303896 190340 303948 190392
rect 304816 190340 304868 190392
rect 439136 190340 439188 190392
rect 440056 190340 440108 190392
rect 168656 190272 168708 190324
rect 169576 190272 169628 190324
rect 320364 190272 320416 190324
rect 321376 190272 321428 190324
rect 328644 190272 328696 190324
rect 329656 190272 329708 190324
rect 219808 190204 219860 190256
rect 220636 190204 220688 190256
rect 332784 190204 332836 190256
rect 333888 190204 333940 190256
rect 355048 190204 355100 190256
rect 355876 190204 355928 190256
rect 443276 190204 443328 190256
rect 444196 190204 444248 190256
rect 201592 190136 201644 190188
rect 202696 190136 202748 190188
rect 281632 190136 281684 190188
rect 282736 190136 282788 190188
rect 408592 190136 408644 190188
rect 409696 190136 409748 190188
rect 416872 190136 416924 190188
rect 417976 190136 418028 190188
rect 154672 190068 154724 190120
rect 155776 190068 155828 190120
rect 244556 190068 244608 190120
rect 245476 190068 245528 190120
rect 253572 190068 253624 190120
rect 257344 190068 257396 190120
rect 316224 190068 316276 190120
rect 317236 190068 317288 190120
rect 353392 190068 353444 190120
rect 354496 190068 354548 190120
rect 379796 190068 379848 190120
rect 380716 190068 380768 190120
rect 441620 190068 441672 190120
rect 442816 190068 442868 190120
rect 361580 190000 361632 190052
rect 362776 190000 362828 190052
rect 369860 190000 369912 190052
rect 371056 190000 371108 190052
rect 433340 190000 433392 190052
rect 434536 190000 434588 190052
rect 237932 189932 237984 189984
rect 238668 189932 238720 189984
rect 269212 189932 269264 189984
rect 270316 189932 270368 189984
rect 270868 189932 270920 189984
rect 271972 189932 272024 189984
rect 340972 189932 341024 189984
rect 342076 189932 342128 189984
rect 373172 189932 373224 189984
rect 373908 189932 373960 189984
rect 421012 189932 421064 189984
rect 422116 189932 422168 189984
rect 158720 189796 158772 189848
rect 159916 189796 159968 189848
rect 176108 189796 176160 189848
rect 184204 189796 184256 189848
rect 240416 189796 240468 189848
rect 255964 189796 256016 189848
rect 257712 189796 257764 189848
rect 301504 189796 301556 189848
rect 448244 189796 448296 189848
rect 456064 189796 456116 189848
rect 180984 189728 181036 189780
rect 192484 189728 192536 189780
rect 195888 189728 195940 189780
rect 213184 189728 213236 189780
rect 223120 189728 223172 189780
rect 242164 189728 242216 189780
rect 274180 189728 274232 189780
rect 280804 189728 280856 189780
rect 294788 189728 294840 189780
rect 352564 189728 352616 189780
rect 359188 189728 359240 189780
rect 381544 189728 381596 189780
rect 383844 189728 383896 189780
rect 485780 189728 485832 189780
rect 229652 189660 229704 189712
rect 230388 189660 230440 189712
rect 309692 189660 309744 189712
rect 310428 189660 310480 189712
rect 334440 189660 334492 189712
rect 335268 189660 335320 189712
rect 364892 189660 364944 189712
rect 365628 189660 365680 189712
rect 428372 189660 428424 189712
rect 429108 189660 429160 189712
rect 234620 189524 234672 189576
rect 235816 189524 235868 189576
rect 397920 189524 397972 189576
rect 398748 189524 398800 189576
rect 449900 189524 449952 189576
rect 451188 189524 451240 189576
rect 222292 189456 222344 189508
rect 223488 189456 223540 189508
rect 250260 189456 250312 189508
rect 251088 189456 251140 189508
rect 285772 189456 285824 189508
rect 286968 189456 287020 189508
rect 322020 189456 322072 189508
rect 322848 189456 322900 189508
rect 330300 189456 330352 189508
rect 331128 189456 331180 189508
rect 387984 189456 388036 189508
rect 389088 189456 389140 189508
rect 175280 189388 175332 189440
rect 176568 189388 176620 189440
rect 182640 189388 182692 189440
rect 183468 189388 183520 189440
rect 203248 189388 203300 189440
rect 204168 189388 204220 189440
rect 275008 189388 275060 189440
rect 275928 189388 275980 189440
rect 293960 189388 294012 189440
rect 295248 189388 295300 189440
rect 317880 189388 317932 189440
rect 318708 189388 318760 189440
rect 346768 189388 346820 189440
rect 347688 189388 347740 189440
rect 410248 189388 410300 189440
rect 411168 189388 411220 189440
rect 447416 189388 447468 189440
rect 448428 189388 448480 189440
rect 156236 189320 156288 189372
rect 157248 189320 157300 189372
rect 164516 189320 164568 189372
rect 165528 189320 165580 189372
rect 172796 189320 172848 189372
rect 173808 189320 173860 189372
rect 197544 189320 197596 189372
rect 198648 189320 198700 189372
rect 214012 189320 214064 189372
rect 215208 189320 215260 189372
rect 236276 189320 236328 189372
rect 237288 189320 237340 189372
rect 261024 189320 261076 189372
rect 262128 189320 262180 189372
rect 277492 189320 277544 189372
rect 278688 189320 278740 189372
rect 299756 189320 299808 189372
rect 300768 189320 300820 189372
rect 349252 189320 349304 189372
rect 350448 189320 350500 189372
rect 371516 189320 371568 189372
rect 372528 189320 372580 189372
rect 412732 189320 412784 189372
rect 413928 189320 413980 189372
rect 434996 189320 435048 189372
rect 436008 189320 436060 189372
rect 185124 189252 185176 189304
rect 186228 189252 186280 189304
rect 193404 189252 193456 189304
rect 194508 189252 194560 189304
rect 205732 189252 205784 189304
rect 206928 189252 206980 189304
rect 209872 189252 209924 189304
rect 211068 189252 211120 189304
rect 223856 189252 223908 189304
rect 224868 189252 224920 189304
rect 230480 189252 230532 189304
rect 231768 189252 231820 189304
rect 238760 189252 238812 189304
rect 240048 189252 240100 189304
rect 248604 189252 248656 189304
rect 249708 189252 249760 189304
rect 265164 189252 265216 189304
rect 266268 189252 266320 189304
rect 302240 189252 302292 189304
rect 303528 189252 303580 189304
rect 306380 189252 306432 189304
rect 307668 189252 307720 189304
rect 310520 189252 310572 189304
rect 311808 189252 311860 189304
rect 312176 189252 312228 189304
rect 313188 189252 313240 189304
rect 336924 189252 336976 189304
rect 338028 189252 338080 189304
rect 345112 189252 345164 189304
rect 346308 189252 346360 189304
rect 365720 189252 365772 189304
rect 367008 189252 367060 189304
rect 374000 189252 374052 189304
rect 375288 189252 375340 189304
rect 375656 189252 375708 189304
rect 376668 189252 376720 189304
rect 378140 189252 378192 189304
rect 379428 189252 379480 189304
rect 400404 189252 400456 189304
rect 401508 189252 401560 189304
rect 437480 189252 437532 189304
rect 438768 189252 438820 189304
rect 160376 189116 160428 189168
rect 161388 189116 161440 189168
rect 213552 189116 213604 189168
rect 221280 189116 221332 189168
rect 283288 189116 283340 189168
rect 284116 189116 284168 189168
rect 307208 189116 307260 189168
rect 309784 189116 309836 189168
rect 378968 189116 379020 189168
rect 384304 189116 384356 189168
rect 418528 189116 418580 189168
rect 419356 189116 419408 189168
rect 445760 189116 445812 189168
rect 451924 189116 451976 189168
rect 157892 189048 157944 189100
rect 158628 189048 158680 189100
rect 162860 189048 162912 189100
rect 164148 189048 164200 189100
rect 166172 189048 166224 189100
rect 166908 189048 166960 189100
rect 167000 189048 167052 189100
rect 168196 189048 168248 189100
rect 171140 189048 171192 189100
rect 172336 189048 172388 189100
rect 174452 189048 174504 189100
rect 175188 189048 175240 189100
rect 176936 189048 176988 189100
rect 177856 189048 177908 189100
rect 178500 189048 178552 189100
rect 179236 189048 179288 189100
rect 186780 189048 186832 189100
rect 187516 189048 187568 189100
rect 189264 189048 189316 189100
rect 190276 189048 190328 189100
rect 190920 189048 190972 189100
rect 191748 189048 191800 189100
rect 195060 189048 195112 189100
rect 195888 189048 195940 189100
rect 199200 189048 199252 189100
rect 200764 189048 200816 189100
rect 207388 189048 207440 189100
rect 208308 189048 208360 189100
rect 211528 189048 211580 189100
rect 212356 189048 212408 189100
rect 215668 189048 215720 189100
rect 216588 189048 216640 189100
rect 218152 189048 218204 189100
rect 219348 189048 219400 189100
rect 221464 189048 221516 189100
rect 222844 189048 222896 189100
rect 226340 189048 226392 189100
rect 227628 189048 227680 189100
rect 227996 189048 228048 189100
rect 229008 189048 229060 189100
rect 232136 189048 232188 189100
rect 233056 189048 233108 189100
rect 242900 189048 242952 189100
rect 244188 189048 244240 189100
rect 246120 189048 246172 189100
rect 246948 189048 247000 189100
rect 256884 189048 256936 189100
rect 257988 189048 258040 189100
rect 258540 189048 258592 189100
rect 259276 189048 259328 189100
rect 262680 189048 262732 189100
rect 263508 189048 263560 189100
rect 266820 189048 266872 189100
rect 267556 189048 267608 189100
rect 273352 189048 273404 189100
rect 274548 189048 274600 189100
rect 279148 189048 279200 189100
rect 279976 189048 280028 189100
rect 287428 189048 287480 189100
rect 288348 189048 288400 189100
rect 289912 189048 289964 189100
rect 291108 189048 291160 189100
rect 291568 189048 291620 189100
rect 292396 189048 292448 189100
rect 293132 189048 293184 189100
rect 293868 189048 293920 189100
rect 298100 189048 298152 189100
rect 299388 189048 299440 189100
rect 301412 189048 301464 189100
rect 302148 189048 302200 189100
rect 308036 189048 308088 189100
rect 308956 189048 309008 189100
rect 324504 189048 324556 189100
rect 327724 189048 327776 189100
rect 338488 189048 338540 189100
rect 339316 189048 339368 189100
rect 342628 189048 342680 189100
rect 344284 189048 344336 189100
rect 350908 189048 350960 189100
rect 351736 189048 351788 189100
rect 357532 189048 357584 189100
rect 358636 189048 358688 189100
rect 363236 189048 363288 189100
rect 364248 189048 364300 189100
rect 381452 189048 381504 189100
rect 382188 189048 382240 189100
rect 382280 189048 382332 189100
rect 383476 189048 383528 189100
rect 385500 189048 385552 189100
rect 386236 189048 386288 189100
rect 389640 189048 389692 189100
rect 390468 189048 390520 189100
rect 392124 189048 392176 189100
rect 393136 189048 393188 189100
rect 402060 189048 402112 189100
rect 402888 189048 402940 189100
rect 404544 189048 404596 189100
rect 405556 189048 405608 189100
rect 406108 189048 406160 189100
rect 406936 189048 406988 189100
rect 414388 189048 414440 189100
rect 416044 189048 416096 189100
rect 422668 189048 422720 189100
rect 423588 189048 423640 189100
rect 425152 189048 425204 189100
rect 426348 189048 426400 189100
rect 426808 189048 426860 189100
rect 427636 189048 427688 189100
rect 429200 189048 429252 189100
rect 430396 189048 430448 189100
rect 430856 189048 430908 189100
rect 431776 189048 431828 189100
rect 436652 189048 436704 189100
rect 437388 189048 437440 189100
rect 444932 189048 444984 189100
rect 445668 189048 445720 189100
rect 235448 188300 235500 188352
rect 271880 188300 271932 188352
rect 271972 188300 272024 188352
rect 322940 188300 322992 188352
rect 386328 188300 386380 188352
rect 489920 188300 489972 188352
rect 252744 186940 252796 186992
rect 296720 186940 296772 186992
rect 388812 186940 388864 186992
rect 494060 186940 494112 186992
rect 138020 185580 138072 185632
rect 138572 185580 138624 185632
rect 139400 185580 139452 185632
rect 140228 185580 140280 185632
rect 143540 185580 143592 185632
rect 144460 185580 144512 185632
rect 146300 185580 146352 185632
rect 146852 185580 146904 185632
rect 147680 185580 147732 185632
rect 148508 185580 148560 185632
rect 393780 185580 393832 185632
rect 500960 185580 501012 185632
rect 396264 184152 396316 184204
rect 503720 184152 503772 184204
rect 398656 182792 398708 182844
rect 507860 182792 507912 182844
rect 453672 182112 453724 182164
rect 580172 182112 580224 182164
rect 133880 181432 133932 181484
rect 134524 181432 134576 181484
rect 367376 181432 367428 181484
rect 462320 181432 462372 181484
rect 3240 180752 3292 180804
rect 17224 180752 17276 180804
rect 401416 180072 401468 180124
rect 512000 180072 512052 180124
rect 275836 178644 275888 178696
rect 331220 178644 331272 178696
rect 406936 178644 406988 178696
rect 518900 178644 518952 178696
rect 259276 177284 259328 177336
rect 305000 177284 305052 177336
rect 314476 177284 314528 177336
rect 385040 177284 385092 177336
rect 409696 177284 409748 177336
rect 521660 177284 521712 177336
rect 411076 175924 411128 175976
rect 525800 175924 525852 175976
rect 413836 174496 413888 174548
rect 528560 174496 528612 174548
rect 135352 173884 135404 173936
rect 135628 173884 135680 173936
rect 419356 173136 419408 173188
rect 536840 173136 536892 173188
rect 422116 171776 422168 171828
rect 539600 171776 539652 171828
rect 453580 171028 453632 171080
rect 580172 171028 580224 171080
rect 423496 168988 423548 169040
rect 543740 168988 543792 169040
rect 426256 167628 426308 167680
rect 546500 167628 546552 167680
rect 431776 166268 431828 166320
rect 554780 166268 554832 166320
rect 3516 165520 3568 165572
rect 126244 165520 126296 165572
rect 434536 164840 434588 164892
rect 557540 164840 557592 164892
rect 135352 164160 135404 164212
rect 135536 164160 135588 164212
rect 435916 163480 435968 163532
rect 561680 163480 561732 163532
rect 438676 162120 438728 162172
rect 564440 162120 564492 162172
rect 444196 160692 444248 160744
rect 571340 160692 571392 160744
rect 364156 159332 364208 159384
rect 458180 159332 458232 159384
rect 471244 158652 471296 158704
rect 579804 158652 579856 158704
rect 366916 157972 366968 158024
rect 460940 157972 460992 158024
rect 376576 156612 376628 156664
rect 476120 156612 476172 156664
rect 383476 155184 383528 155236
rect 484400 155184 484452 155236
rect 384948 153824 385000 153876
rect 487160 153824 487212 153876
rect 393136 152464 393188 152516
rect 498200 152464 498252 152516
rect 3148 151716 3200 151768
rect 129280 151716 129332 151768
rect 397368 151036 397420 151088
rect 505100 151036 505152 151088
rect 405556 149676 405608 149728
rect 516140 149676 516192 149728
rect 416044 148316 416096 148368
rect 529940 148316 529992 148368
rect 417976 146888 418028 146940
rect 534080 146888 534132 146940
rect 427636 145528 427688 145580
rect 547880 145528 547932 145580
rect 430396 144168 430448 144220
rect 552020 144168 552072 144220
rect 440056 142808 440108 142860
rect 565820 142808 565872 142860
rect 442816 141380 442868 141432
rect 569960 141380 570012 141432
rect 371056 140020 371108 140072
rect 466460 140020 466512 140072
rect 375196 138660 375248 138712
rect 473360 138660 473412 138712
rect 380716 137232 380768 137284
rect 480260 137232 480312 137284
rect 3240 136552 3292 136604
rect 13084 136552 13136 136604
rect 390376 135872 390428 135924
rect 495440 135872 495492 135924
rect 479524 135192 479576 135244
rect 580172 135192 580224 135244
rect 313096 134512 313148 134564
rect 383660 134512 383712 134564
rect 384304 134512 384356 134564
rect 478880 134512 478932 134564
rect 402796 133152 402848 133204
rect 513380 133152 513432 133204
rect 415308 131724 415360 131776
rect 531320 131724 531372 131776
rect 433248 130364 433300 130416
rect 556160 130364 556212 130416
rect 453488 124108 453540 124160
rect 580172 124108 580224 124160
rect 3424 122748 3476 122800
rect 14464 122748 14516 122800
rect 311716 117920 311768 117972
rect 382280 117920 382332 117972
rect 307668 113772 307720 113824
rect 374000 113772 374052 113824
rect 469864 111732 469916 111784
rect 579804 111732 579856 111784
rect 372436 111052 372488 111104
rect 469220 111052 469272 111104
rect 331036 109692 331088 109744
rect 409880 109692 409932 109744
rect 3240 108944 3292 108996
rect 129188 108944 129240 108996
rect 321376 108264 321428 108316
rect 394700 108264 394752 108316
rect 395988 108264 396040 108316
rect 502340 108264 502392 108316
rect 354496 105544 354548 105596
rect 443000 105544 443052 105596
rect 326896 104116 326948 104168
rect 402980 104116 403032 104168
rect 351736 102756 351788 102808
rect 438860 102756 438912 102808
rect 339316 101396 339368 101448
rect 420920 101396 420972 101448
rect 346216 99968 346268 100020
rect 431960 99968 432012 100020
rect 343548 98608 343600 98660
rect 427820 98608 427872 98660
rect 342076 97248 342128 97300
rect 425060 97248 425112 97300
rect 336648 95888 336700 95940
rect 416780 95888 416832 95940
rect 333796 94460 333848 94512
rect 414020 94460 414072 94512
rect 3424 93780 3476 93832
rect 19984 93780 20036 93832
rect 329656 93100 329708 93152
rect 407120 93100 407172 93152
rect 324228 91740 324280 91792
rect 400220 91740 400272 91792
rect 321468 90312 321520 90364
rect 396080 90312 396132 90364
rect 318616 88952 318668 89004
rect 391940 88952 391992 89004
rect 472624 88272 472676 88324
rect 580172 88272 580224 88324
rect 375288 87592 375340 87644
rect 471980 87592 472032 87644
rect 135444 86912 135496 86964
rect 317236 86232 317288 86284
rect 389180 86232 389232 86284
rect 438768 86232 438820 86284
rect 563060 86232 563112 86284
rect 304816 84804 304868 84856
rect 371240 84804 371292 84856
rect 302148 83444 302200 83496
rect 367100 83444 367152 83496
rect 430488 83444 430540 83496
rect 553400 83444 553452 83496
rect 299296 82084 299348 82136
rect 364340 82084 364392 82136
rect 398748 82084 398800 82136
rect 506480 82084 506532 82136
rect 295248 80656 295300 80708
rect 356060 80656 356112 80708
rect 365628 80656 365680 80708
rect 459652 80656 459704 80708
rect 3516 79432 3568 79484
rect 8944 79432 8996 79484
rect 292396 79296 292448 79348
rect 353300 79296 353352 79348
rect 401508 79296 401560 79348
rect 510620 79296 510672 79348
rect 289728 77936 289780 77988
rect 349160 77936 349212 77988
rect 418068 77936 418120 77988
rect 535460 77936 535512 77988
rect 135352 77299 135404 77308
rect 135352 77265 135361 77299
rect 135361 77265 135395 77299
rect 135395 77265 135404 77299
rect 135352 77256 135404 77265
rect 453396 77188 453448 77240
rect 580172 77188 580224 77240
rect 135352 77163 135404 77172
rect 135352 77129 135361 77163
rect 135361 77129 135395 77163
rect 135395 77129 135404 77163
rect 135352 77120 135404 77129
rect 286876 76508 286928 76560
rect 346400 76508 346452 76560
rect 349068 76508 349120 76560
rect 434720 76508 434772 76560
rect 335176 75148 335228 75200
rect 416872 75148 416924 75200
rect 423588 75148 423640 75200
rect 542360 75148 542412 75200
rect 282736 73788 282788 73840
rect 339500 73788 339552 73840
rect 355876 73788 355928 73840
rect 444380 73788 444432 73840
rect 445668 73788 445720 73840
rect 573364 73788 573416 73840
rect 333888 72428 333940 72480
rect 412640 72428 412692 72480
rect 420828 72428 420880 72480
rect 538220 72428 538272 72480
rect 279976 71000 280028 71052
rect 335360 71000 335412 71052
rect 347596 71000 347648 71052
rect 433340 71000 433392 71052
rect 436008 71000 436060 71052
rect 560300 71000 560352 71052
rect 135444 70252 135496 70304
rect 331128 69640 331180 69692
rect 408500 69640 408552 69692
rect 411168 69640 411220 69692
rect 524420 69640 524472 69692
rect 271788 68280 271840 68332
rect 324320 68280 324372 68332
rect 328368 68280 328420 68332
rect 405740 68280 405792 68332
rect 408408 68280 408460 68332
rect 520280 68280 520332 68332
rect 270316 66852 270368 66904
rect 321560 66852 321612 66904
rect 325608 66852 325660 66904
rect 401600 66852 401652 66904
rect 413928 66852 413980 66904
rect 528652 66852 528704 66904
rect 267556 65492 267608 65544
rect 317420 65492 317472 65544
rect 322756 65492 322808 65544
rect 398840 65492 398892 65544
rect 405648 65492 405700 65544
rect 517520 65492 517572 65544
rect 3332 64812 3384 64864
rect 129096 64812 129148 64864
rect 454684 64812 454736 64864
rect 579804 64812 579856 64864
rect 262036 64132 262088 64184
rect 310520 64132 310572 64184
rect 362776 64132 362828 64184
rect 454040 64132 454092 64184
rect 259368 62772 259420 62824
rect 306380 62772 306432 62824
rect 318708 62772 318760 62824
rect 390560 62772 390612 62824
rect 393228 62772 393280 62824
rect 499580 62772 499632 62824
rect 306288 61344 306340 61396
rect 374092 61344 374144 61396
rect 389088 61344 389140 61396
rect 492680 61344 492732 61396
rect 135444 60664 135496 60716
rect 135628 60664 135680 60716
rect 257988 59984 258040 60036
rect 303620 59984 303672 60036
rect 308956 59984 309008 60036
rect 376760 59984 376812 60036
rect 386236 59984 386288 60036
rect 488540 59984 488592 60036
rect 255136 58624 255188 58676
rect 299480 58624 299532 58676
rect 303436 58624 303488 58676
rect 369860 58624 369912 58676
rect 383568 58624 383620 58676
rect 485872 58624 485924 58676
rect 135628 57876 135680 57928
rect 249616 57196 249668 57248
rect 292580 57196 292632 57248
rect 300676 57196 300728 57248
rect 365720 57196 365772 57248
rect 378048 57196 378100 57248
rect 477592 57196 477644 57248
rect 299388 55904 299440 55956
rect 362960 55904 363012 55956
rect 362868 55836 362920 55888
rect 455420 55836 455472 55888
rect 246856 54476 246908 54528
rect 288440 54476 288492 54528
rect 296536 54476 296588 54528
rect 358820 54476 358872 54528
rect 360108 54476 360160 54528
rect 451280 54476 451332 54528
rect 245476 53048 245528 53100
rect 285680 53048 285732 53100
rect 293868 53048 293920 53100
rect 356152 53048 356204 53100
rect 358636 53048 358688 53100
rect 448520 53048 448572 53100
rect 242808 51688 242860 51740
rect 281540 51688 281592 51740
rect 291016 51688 291068 51740
rect 351920 51688 351972 51740
rect 353208 51688 353260 51740
rect 441620 51688 441672 51740
rect 3424 51008 3476 51060
rect 15844 51008 15896 51060
rect 239956 50328 240008 50380
rect 278780 50328 278832 50380
rect 288256 50328 288308 50380
rect 347780 50328 347832 50380
rect 350356 50328 350408 50380
rect 437480 50328 437532 50380
rect 442908 50328 442960 50380
rect 571432 50328 571484 50380
rect 233056 48968 233108 49020
rect 267740 48968 267792 49020
rect 284116 48968 284168 49020
rect 340880 48968 340932 49020
rect 344284 48968 344336 49020
rect 426440 48968 426492 49020
rect 427728 48968 427780 49020
rect 549260 48968 549312 49020
rect 135536 48331 135588 48340
rect 135536 48297 135545 48331
rect 135545 48297 135579 48331
rect 135579 48297 135588 48331
rect 135536 48288 135588 48297
rect 237196 47540 237248 47592
rect 274640 47540 274692 47592
rect 281448 47540 281500 47592
rect 338120 47540 338172 47592
rect 340788 47540 340840 47592
rect 423680 47540 423732 47592
rect 447048 47540 447100 47592
rect 574744 47540 574796 47592
rect 244096 46180 244148 46232
rect 284300 46180 284352 46232
rect 286968 46180 287020 46232
rect 345020 46180 345072 46232
rect 346308 46180 346360 46232
rect 430580 46180 430632 46232
rect 440148 46180 440200 46232
rect 567200 46180 567252 46232
rect 235816 44820 235868 44872
rect 270500 44820 270552 44872
rect 278596 44820 278648 44872
rect 333980 44820 334032 44872
rect 337936 44820 337988 44872
rect 419540 44820 419592 44872
rect 426348 44820 426400 44872
rect 546592 44820 546644 44872
rect 230388 43392 230440 43444
rect 263600 43392 263652 43444
rect 274548 43392 274600 43444
rect 327080 43392 327132 43444
rect 347688 43392 347740 43444
rect 433432 43392 433484 43444
rect 434628 43392 434680 43444
rect 558920 43392 558972 43444
rect 266176 42100 266228 42152
rect 316040 42100 316092 42152
rect 227536 42032 227588 42084
rect 260840 42032 260892 42084
rect 315948 42032 316000 42084
rect 387800 42032 387852 42084
rect 424968 42032 425020 42084
rect 545120 42032 545172 42084
rect 135444 41352 135496 41404
rect 135628 41352 135680 41404
rect 478144 41352 478196 41404
rect 580172 41352 580224 41404
rect 224776 40672 224828 40724
rect 256700 40672 256752 40724
rect 263416 40672 263468 40724
rect 313280 40672 313332 40724
rect 339408 40672 339460 40724
rect 422300 40672 422352 40724
rect 296628 39380 296680 39432
rect 360200 39380 360252 39432
rect 223488 39312 223540 39364
rect 252560 39312 252612 39364
rect 262128 39312 262180 39364
rect 309140 39312 309192 39364
rect 357348 39312 357400 39364
rect 447140 39312 447192 39364
rect 449808 39312 449860 39364
rect 574836 39312 574888 39364
rect 135628 38564 135680 38616
rect 220636 37884 220688 37936
rect 249800 37884 249852 37936
rect 256608 37884 256660 37936
rect 302240 37884 302292 37936
rect 335268 37884 335320 37936
rect 415400 37884 415452 37936
rect 422208 37884 422260 37936
rect 540980 37884 541032 37936
rect 250996 36592 251048 36644
rect 295340 36592 295392 36644
rect 217968 36524 218020 36576
rect 245660 36524 245712 36576
rect 284208 36524 284260 36576
rect 342260 36524 342312 36576
rect 351828 36524 351880 36576
rect 440240 36524 440292 36576
rect 444288 36524 444340 36576
rect 572720 36524 572772 36576
rect 3424 35844 3476 35896
rect 11704 35844 11756 35896
rect 277308 35232 277360 35284
rect 331312 35232 331364 35284
rect 215116 35164 215168 35216
rect 242900 35164 242952 35216
rect 249708 35164 249760 35216
rect 291200 35164 291252 35216
rect 327724 35164 327776 35216
rect 400312 35164 400364 35216
rect 402888 35164 402940 35216
rect 512092 35164 512144 35216
rect 241428 33736 241480 33788
rect 280160 33736 280212 33788
rect 280804 33736 280856 33788
rect 328460 33736 328512 33788
rect 329748 33736 329800 33788
rect 408592 33736 408644 33788
rect 409788 33736 409840 33788
rect 523040 33736 523092 33788
rect 240048 32444 240100 32496
rect 277400 32444 277452 32496
rect 264888 32376 264940 32428
rect 313372 32376 313424 32428
rect 314568 32376 314620 32428
rect 386420 32376 386472 32428
rect 387708 32376 387760 32428
rect 491300 32376 491352 32428
rect 237288 31084 237340 31136
rect 273260 31084 273312 31136
rect 269028 31016 269080 31068
rect 320180 31016 320232 31068
rect 326988 31016 327040 31068
rect 404360 31016 404412 31068
rect 407028 31016 407080 31068
rect 520372 31016 520424 31068
rect 453304 30268 453356 30320
rect 580172 30268 580224 30320
rect 227628 29656 227680 29708
rect 259460 29656 259512 29708
rect 252468 29588 252520 29640
rect 296812 29588 296864 29640
rect 304908 29588 304960 29640
rect 372620 29588 372672 29640
rect 135536 29019 135588 29028
rect 135536 28985 135545 29019
rect 135545 28985 135579 29019
rect 135579 28985 135588 29019
rect 135536 28976 135588 28985
rect 224868 28228 224920 28280
rect 255320 28228 255372 28280
rect 257344 28228 257396 28280
rect 298100 28228 298152 28280
rect 303528 28228 303580 28280
rect 368480 28228 368532 28280
rect 369768 28228 369820 28280
rect 465080 28228 465132 28280
rect 216496 26868 216548 26920
rect 244280 26868 244332 26920
rect 246948 26868 247000 26920
rect 287060 26868 287112 26920
rect 298008 26868 298060 26920
rect 361580 26868 361632 26920
rect 372528 26868 372580 26920
rect 467932 26868 467984 26920
rect 212356 25576 212408 25628
rect 237380 25576 237432 25628
rect 234528 25508 234580 25560
rect 270592 25508 270644 25560
rect 292488 25508 292540 25560
rect 354680 25508 354732 25560
rect 441528 25508 441580 25560
rect 568580 25508 568632 25560
rect 206836 24080 206888 24132
rect 230480 24080 230532 24132
rect 231676 24080 231728 24132
rect 266360 24080 266412 24132
rect 282828 24080 282880 24132
rect 339592 24080 339644 24132
rect 342168 24080 342220 24132
rect 425152 24080 425204 24132
rect 431868 24080 431920 24132
rect 554872 24080 554924 24132
rect 204076 22720 204128 22772
rect 227812 22720 227864 22772
rect 228916 22720 228968 22772
rect 262220 22720 262272 22772
rect 280068 22720 280120 22772
rect 336740 22720 336792 22772
rect 338028 22720 338080 22772
rect 418160 22720 418212 22772
rect 419448 22720 419500 22772
rect 536932 22720 536984 22772
rect 3148 22040 3200 22092
rect 129004 22040 129056 22092
rect 135444 22040 135496 22092
rect 135628 22040 135680 22092
rect 202696 21428 202748 21480
rect 223580 21428 223632 21480
rect 278688 21428 278740 21480
rect 332600 21428 332652 21480
rect 222844 21360 222896 21412
rect 252652 21360 252704 21412
rect 332508 21360 332560 21412
rect 411260 21360 411312 21412
rect 412548 21360 412600 21412
rect 527180 21360 527232 21412
rect 200764 20000 200816 20052
rect 219440 20000 219492 20052
rect 219256 19932 219308 19984
rect 248420 19932 248472 19984
rect 266268 19932 266320 19984
rect 314660 19932 314712 19984
rect 317328 19932 317380 19984
rect 390652 19932 390704 19984
rect 429108 19932 429160 19984
rect 550640 19932 550692 19984
rect 135628 19295 135680 19304
rect 135628 19261 135637 19295
rect 135637 19261 135671 19295
rect 135671 19261 135680 19295
rect 135628 19252 135680 19261
rect 301504 19252 301556 19304
rect 305092 19252 305144 19304
rect 197268 18640 197320 18692
rect 216680 18640 216732 18692
rect 215208 18572 215260 18624
rect 241520 18572 241572 18624
rect 251088 18572 251140 18624
rect 293960 18572 294012 18624
rect 310428 18572 310480 18624
rect 379520 18572 379572 18624
rect 400128 18572 400180 18624
rect 509240 18572 509292 18624
rect 483664 17892 483716 17944
rect 579804 17892 579856 17944
rect 194416 17280 194468 17332
rect 212540 17280 212592 17332
rect 209688 17212 209740 17264
rect 234620 17212 234672 17264
rect 244188 17212 244240 17264
rect 282920 17212 282972 17264
rect 285588 17212 285640 17264
rect 343640 17212 343692 17264
rect 344928 17212 344980 17264
rect 429200 17212 429252 17264
rect 255228 15920 255280 15972
rect 300860 15920 300912 15972
rect 191656 15852 191708 15904
rect 209872 15852 209924 15904
rect 220728 15852 220780 15904
rect 251180 15852 251232 15904
rect 300768 15852 300820 15904
rect 365812 15852 365864 15904
rect 390468 15852 390520 15904
rect 494152 15852 494204 15904
rect 190276 14424 190328 14476
rect 205640 14424 205692 14476
rect 216588 14424 216640 14476
rect 244372 14424 244424 14476
rect 245568 14424 245620 14476
rect 287152 14424 287204 14476
rect 288348 14424 288400 14476
rect 347872 14424 347924 14476
rect 350448 14424 350500 14476
rect 436100 14424 436152 14476
rect 437388 14424 437440 14476
rect 563152 14424 563204 14476
rect 208216 13132 208268 13184
rect 233240 13132 233292 13184
rect 187516 13064 187568 13116
rect 201500 13064 201552 13116
rect 233148 13064 233200 13116
rect 269120 13064 269172 13116
rect 270408 13064 270460 13116
rect 321652 13064 321704 13116
rect 322848 13064 322900 13116
rect 397460 13064 397512 13116
rect 416688 13064 416740 13116
rect 532700 13064 532752 13116
rect 135628 12291 135680 12300
rect 135628 12257 135637 12291
rect 135637 12257 135671 12291
rect 135671 12257 135680 12291
rect 135628 12248 135680 12257
rect 184848 11704 184900 11756
rect 198740 11704 198792 11756
rect 204168 11704 204220 11756
rect 226340 11704 226392 11756
rect 229008 11704 229060 11756
rect 262312 11704 262364 11756
rect 263508 11704 263560 11756
rect 311900 11704 311952 11756
rect 313188 11704 313240 11756
rect 382372 11704 382424 11756
rect 404268 11704 404320 11756
rect 514760 11704 514812 11756
rect 188988 10276 189040 10328
rect 204260 10276 204312 10328
rect 206928 10276 206980 10328
rect 229100 10276 229152 10328
rect 231768 10276 231820 10328
rect 264980 10276 265032 10328
rect 267648 10276 267700 10328
rect 318800 10276 318852 10328
rect 320088 10276 320140 10328
rect 393320 10276 393372 10328
rect 394608 10276 394660 10328
rect 502432 10276 502484 10328
rect 186136 8984 186188 9036
rect 201592 8984 201644 9036
rect 201408 8916 201460 8968
rect 222936 8916 222988 8968
rect 226248 8916 226300 8968
rect 258632 8916 258684 8968
rect 260748 8916 260800 8968
rect 308588 8916 308640 8968
rect 309784 8916 309836 8968
rect 376392 8916 376444 8968
rect 381544 8916 381596 8968
rect 451372 8916 451424 8968
rect 456064 8916 456116 8968
rect 579804 8916 579856 8968
rect 3424 8236 3476 8288
rect 10324 8236 10376 8288
rect 183376 7556 183428 7608
rect 198004 7556 198056 7608
rect 198556 7556 198608 7608
rect 219348 7556 219400 7608
rect 247960 7556 248012 7608
rect 248328 7556 248380 7608
rect 290740 7556 290792 7608
rect 291108 7556 291160 7608
rect 351368 7556 351420 7608
rect 354588 7556 354640 7608
rect 444196 7556 444248 7608
rect 451924 7556 451976 7608
rect 576216 7556 576268 7608
rect 219348 7352 219400 7404
rect 273168 6196 273220 6248
rect 326436 6196 326488 6248
rect 179236 6128 179288 6180
rect 190828 6128 190880 6180
rect 191748 6128 191800 6180
rect 208676 6128 208728 6180
rect 210976 6128 211028 6180
rect 237196 6128 237248 6180
rect 238668 6128 238720 6180
rect 276480 6128 276532 6180
rect 311808 6128 311860 6180
rect 381176 6128 381228 6180
rect 391848 6128 391900 6180
rect 497740 6128 497792 6180
rect 275928 4836 275980 4888
rect 330024 4836 330076 4888
rect 352564 4836 352616 4888
rect 358544 4836 358596 4888
rect 173716 4768 173768 4820
rect 183744 4768 183796 4820
rect 194508 4768 194560 4820
rect 212264 4768 212316 4820
rect 221464 4768 221516 4820
rect 240784 4768 240836 4820
rect 242164 4768 242216 4820
rect 255044 4768 255096 4820
rect 255964 4768 256016 4820
rect 280068 4768 280120 4820
rect 309048 4768 309100 4820
rect 378784 4768 378836 4820
rect 382188 4768 382240 4820
rect 483480 4768 483532 4820
rect 184204 4156 184256 4208
rect 187240 4156 187292 4208
rect 192484 4156 192536 4208
rect 194416 4156 194468 4208
rect 213184 4156 213236 4208
rect 215852 4156 215904 4208
rect 408500 4156 408552 4208
rect 409696 4156 409748 4208
rect 425152 4156 425204 4208
rect 426348 4156 426400 4208
rect 451280 4156 451332 4208
rect 452476 4156 452528 4208
rect 127808 4088 127860 4140
rect 133880 4088 133932 4140
rect 142068 4088 142120 4140
rect 143540 4088 143592 4140
rect 160008 4088 160060 4140
rect 163504 4088 163556 4140
rect 166908 4088 166960 4140
rect 172980 4088 173032 4140
rect 361488 4088 361540 4140
rect 453672 4088 453724 4140
rect 574744 4088 574796 4140
rect 577412 4088 577464 4140
rect 130200 4020 130252 4072
rect 135628 4020 135680 4072
rect 139676 4020 139728 4072
rect 142436 4020 142488 4072
rect 159916 4020 159968 4072
rect 162308 4020 162360 4072
rect 176568 4020 176620 4072
rect 186044 4020 186096 4072
rect 367008 4020 367060 4072
rect 460848 4020 460900 4072
rect 129004 3952 129056 4004
rect 135260 3952 135312 4004
rect 140872 3952 140924 4004
rect 143632 3952 143684 4004
rect 175188 3952 175240 4004
rect 184848 3952 184900 4004
rect 205548 3952 205600 4004
rect 364248 3952 364300 4004
rect 457260 3952 457312 4004
rect 138480 3884 138532 3936
rect 142160 3884 142212 3936
rect 169576 3884 169628 3936
rect 176568 3884 176620 3936
rect 177856 3884 177908 3936
rect 188436 3884 188488 3936
rect 195888 3884 195940 3936
rect 214656 3884 214708 3936
rect 368388 3884 368440 3936
rect 464436 3884 464488 3936
rect 168196 3816 168248 3868
rect 174176 3816 174228 3868
rect 182088 3816 182140 3868
rect 195612 3816 195664 3868
rect 198648 3816 198700 3868
rect 218152 3816 218204 3868
rect 371148 3816 371200 3868
rect 467840 3816 467892 3868
rect 169668 3748 169720 3800
rect 177764 3748 177816 3800
rect 183468 3748 183520 3800
rect 196808 3748 196860 3800
rect 200028 3748 200080 3800
rect 373908 3748 373960 3800
rect 471520 3748 471572 3800
rect 126612 3680 126664 3732
rect 133972 3680 134024 3732
rect 180708 3680 180760 3732
rect 193220 3680 193272 3732
rect 202788 3680 202840 3732
rect 172428 3612 172480 3664
rect 181352 3612 181404 3664
rect 186228 3612 186280 3664
rect 200396 3612 200448 3664
rect 146852 3544 146904 3596
rect 147772 3544 147824 3596
rect 161388 3544 161440 3596
rect 164700 3544 164752 3596
rect 173808 3544 173860 3596
rect 182548 3544 182600 3596
rect 187608 3544 187660 3596
rect 203892 3612 203944 3664
rect 208308 3680 208360 3732
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 228916 3680 228968 3732
rect 376668 3680 376720 3732
rect 475108 3680 475160 3732
rect 225328 3612 225380 3664
rect 379428 3612 379480 3664
rect 478696 3612 478748 3664
rect 574836 3612 574888 3664
rect 581000 3612 581052 3664
rect 232504 3544 232556 3596
rect 262220 3544 262272 3596
rect 263416 3544 263468 3596
rect 270500 3544 270552 3596
rect 271696 3544 271748 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 365720 3544 365772 3596
rect 366916 3544 366968 3596
rect 374000 3544 374052 3596
rect 375196 3544 375248 3596
rect 380808 3544 380860 3596
rect 482284 3544 482336 3596
rect 485780 3544 485832 3596
rect 486976 3544 487028 3596
rect 494152 3544 494204 3596
rect 495348 3544 495400 3596
rect 520280 3544 520332 3596
rect 521476 3544 521528 3596
rect 528560 3544 528612 3596
rect 529848 3544 529900 3596
rect 536932 3544 536984 3596
rect 538128 3544 538180 3596
rect 546500 3544 546552 3596
rect 547696 3544 547748 3596
rect 573364 3544 573416 3596
rect 575020 3544 575072 3596
rect 572 3476 624 3528
rect 131120 3476 131172 3528
rect 137284 3476 137336 3528
rect 140780 3476 140832 3528
rect 145656 3476 145708 3528
rect 146300 3476 146352 3528
rect 150624 3476 150676 3528
rect 151544 3476 151596 3528
rect 151820 3476 151872 3528
rect 152740 3476 152792 3528
rect 153108 3476 153160 3528
rect 153936 3476 153988 3528
rect 155776 3476 155828 3528
rect 156328 3476 156380 3528
rect 157248 3476 157300 3528
rect 158720 3476 158772 3528
rect 165528 3476 165580 3528
rect 170588 3476 170640 3528
rect 171048 3476 171100 3528
rect 178960 3476 179012 3528
rect 179328 3476 179380 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 211068 3476 211120 3528
rect 1676 3408 1728 3460
rect 132500 3408 132552 3460
rect 134892 3408 134944 3460
rect 139492 3408 139544 3460
rect 144460 3408 144512 3460
rect 146392 3408 146444 3460
rect 154488 3408 154540 3460
rect 155132 3408 155184 3460
rect 158628 3408 158680 3460
rect 161112 3408 161164 3460
rect 161296 3408 161348 3460
rect 165896 3408 165948 3460
rect 168288 3408 168340 3460
rect 175372 3408 175424 3460
rect 177948 3408 178000 3460
rect 189632 3408 189684 3460
rect 190368 3408 190420 3460
rect 207480 3408 207532 3460
rect 210976 3408 211028 3460
rect 236000 3476 236052 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 252560 3476 252612 3528
rect 253848 3476 253900 3528
rect 287060 3476 287112 3528
rect 288348 3476 288400 3528
rect 296720 3476 296772 3528
rect 297916 3476 297968 3528
rect 305000 3476 305052 3528
rect 306196 3476 306248 3528
rect 313372 3476 313424 3528
rect 314568 3476 314620 3528
rect 347780 3476 347832 3528
rect 349068 3476 349120 3528
rect 356060 3476 356112 3528
rect 357348 3476 357400 3528
rect 358728 3476 358780 3528
rect 450176 3476 450228 3528
rect 451188 3476 451240 3528
rect 582196 3476 582248 3528
rect 212448 3408 212500 3460
rect 239588 3408 239640 3460
rect 355968 3408 356020 3460
rect 446588 3408 446640 3460
rect 448428 3408 448480 3460
rect 578608 3408 578660 3460
rect 164056 3340 164108 3392
rect 169392 3340 169444 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 416780 3340 416832 3392
rect 417976 3340 418028 3392
rect 433340 3340 433392 3392
rect 434628 3340 434680 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 133788 3272 133840 3324
rect 138020 3272 138072 3324
rect 155868 3272 155920 3324
rect 157524 3272 157576 3324
rect 162768 3272 162820 3324
rect 167092 3272 167144 3324
rect 172336 3272 172388 3324
rect 180156 3272 180208 3324
rect 136088 3204 136140 3256
rect 139400 3204 139452 3256
rect 164148 3204 164200 3256
rect 168196 3204 168248 3256
rect 132592 3136 132644 3188
rect 138112 3136 138164 3188
rect 131396 3068 131448 3120
rect 136640 3068 136692 3120
rect 221740 3068 221792 3120
rect 157156 3000 157208 3052
rect 159916 3000 159968 3052
rect 143264 2864 143316 2916
rect 144920 2864 144972 2916
rect 165436 2864 165488 2916
rect 171784 2864 171836 2916
rect 502340 2728 502392 2780
rect 503628 2728 503680 2780
rect 563060 2728 563112 2780
rect 564348 2728 564400 2780
rect 571340 2728 571392 2780
rect 572628 2728 572680 2780
rect 364340 552 364392 604
rect 364524 552 364576 604
rect 367100 552 367152 604
rect 368020 552 368072 604
rect 368480 552 368532 604
rect 369216 552 369268 604
rect 369860 552 369912 604
rect 370412 552 370464 604
rect 372620 552 372672 604
rect 372804 552 372856 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 8128 679046 8156 685850
rect 8944 681760 8996 681766
rect 8944 681702 8996 681708
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 589286 8064 591926
rect 8024 589280 8076 589286
rect 8024 589222 8076 589228
rect 8024 579760 8076 579766
rect 7944 579708 8024 579714
rect 7944 579702 8076 579708
rect 7944 579686 8064 579702
rect 7944 579630 7972 579686
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 8116 579624 8168 579630
rect 8116 579566 8168 579572
rect 4066 567352 4122 567361
rect 4066 567287 4068 567296
rect 4120 567287 4122 567296
rect 4068 567258 4120 567264
rect 8128 562970 8156 579566
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 8116 562964 8168 562970
rect 8116 562906 8168 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 2870 509960 2926 509969
rect 2870 509895 2926 509904
rect 2884 509318 2912 509895
rect 2872 509312 2924 509318
rect 2872 509254 2924 509260
rect 3330 481128 3386 481137
rect 3330 481063 3386 481072
rect 3344 480282 3372 481063
rect 3332 480276 3384 480282
rect 3332 480218 3384 480224
rect 3436 455394 3464 553007
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8208 543788 8260 543794
rect 8208 543730 8260 543736
rect 8220 540977 8248 543730
rect 7930 540968 7986 540977
rect 7930 540903 7986 540912
rect 8206 540968 8262 540977
rect 8206 540903 8262 540912
rect 3698 538656 3754 538665
rect 3698 538591 3754 538600
rect 3712 538286 3740 538591
rect 3700 538280 3752 538286
rect 3700 538222 3752 538228
rect 7944 531350 7972 540903
rect 8036 531350 8064 531381
rect 7932 531344 7984 531350
rect 7932 531286 7984 531292
rect 8024 531344 8076 531350
rect 8114 531312 8170 531321
rect 8076 531292 8114 531298
rect 8024 531286 8114 531292
rect 8036 531270 8114 531286
rect 8114 531247 8170 531256
rect 8298 531312 8354 531321
rect 8298 531247 8354 531256
rect 8312 524346 8340 531247
rect 8116 524340 8168 524346
rect 8116 524282 8168 524288
rect 8300 524340 8352 524346
rect 8300 524282 8352 524288
rect 8128 515438 8156 524282
rect 8116 515432 8168 515438
rect 8116 515374 8168 515380
rect 8956 509250 8984 681702
rect 17224 667956 17276 667962
rect 17224 667898 17276 667904
rect 14464 652792 14516 652798
rect 14464 652734 14516 652740
rect 10324 623824 10376 623830
rect 10324 623766 10376 623772
rect 8944 509244 8996 509250
rect 8944 509186 8996 509192
rect 3514 495544 3570 495553
rect 3514 495479 3570 495488
rect 3424 455388 3476 455394
rect 3424 455330 3476 455336
rect 3146 452432 3202 452441
rect 3146 452367 3202 452376
rect 3160 451314 3188 452367
rect 3148 451308 3200 451314
rect 3148 451250 3200 451256
rect 3422 438016 3478 438025
rect 3422 437951 3478 437960
rect 3436 409834 3464 437951
rect 3528 433294 3556 495479
rect 10336 485790 10364 623766
rect 13084 594856 13136 594862
rect 13084 594798 13136 594804
rect 13096 567866 13124 594798
rect 13084 567860 13136 567866
rect 13084 567802 13136 567808
rect 11704 567316 11756 567322
rect 11704 567258 11756 567264
rect 10324 485784 10376 485790
rect 10324 485726 10376 485732
rect 8944 480276 8996 480282
rect 8944 480218 8996 480224
rect 3516 433288 3568 433294
rect 3516 433230 3568 433236
rect 8956 425066 8984 480218
rect 11716 463690 11744 567258
rect 13084 509312 13136 509318
rect 13084 509254 13136 509260
rect 11704 463684 11756 463690
rect 11704 463626 11756 463632
rect 13096 440230 13124 509254
rect 14476 494018 14504 652734
rect 15844 538280 15896 538286
rect 15844 538222 15896 538228
rect 14464 494012 14516 494018
rect 14464 493954 14516 493960
rect 15856 448526 15884 538222
rect 17236 502314 17264 667898
rect 19984 610020 20036 610026
rect 19984 609962 20036 609968
rect 17224 502308 17276 502314
rect 17224 502250 17276 502256
rect 19996 478854 20024 609962
rect 24780 515506 24808 699654
rect 41340 515574 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 72884 637560 72936 637566
rect 72884 637502 72936 637508
rect 72896 630578 72924 637502
rect 72896 630550 73108 630578
rect 73080 626550 73108 630550
rect 73068 626544 73120 626550
rect 73068 626486 73120 626492
rect 73068 616888 73120 616894
rect 73068 616830 73120 616836
rect 73080 611454 73108 616830
rect 73068 611448 73120 611454
rect 73068 611390 73120 611396
rect 72884 611312 72936 611318
rect 72884 611254 72936 611260
rect 72896 608546 72924 611254
rect 72974 608560 73030 608569
rect 72896 608518 72974 608546
rect 72974 608495 73030 608504
rect 73158 608560 73214 608569
rect 73158 608495 73214 608504
rect 73172 601594 73200 608495
rect 72976 601588 73028 601594
rect 72976 601530 73028 601536
rect 73160 601588 73212 601594
rect 73160 601530 73212 601536
rect 72988 598942 73016 601530
rect 72976 598936 73028 598942
rect 72976 598878 73028 598884
rect 72884 589348 72936 589354
rect 72884 589290 72936 589296
rect 72896 582418 72924 589290
rect 72700 582412 72752 582418
rect 72700 582354 72752 582360
rect 72884 582412 72936 582418
rect 72884 582354 72936 582360
rect 72712 579630 72740 582354
rect 72700 579624 72752 579630
rect 72700 579566 72752 579572
rect 72608 569968 72660 569974
rect 72608 569910 72660 569916
rect 72620 563106 72648 569910
rect 72608 563100 72660 563106
rect 72608 563042 72660 563048
rect 72700 562964 72752 562970
rect 72700 562906 72752 562912
rect 72712 560250 72740 562906
rect 72700 560244 72752 560250
rect 72700 560186 72752 560192
rect 72884 550656 72936 550662
rect 72884 550598 72936 550604
rect 72896 543658 72924 550598
rect 72700 543652 72752 543658
rect 72700 543594 72752 543600
rect 72884 543652 72936 543658
rect 72884 543594 72936 543600
rect 72712 534070 72740 543594
rect 72700 534064 72752 534070
rect 72700 534006 72752 534012
rect 72884 534064 72936 534070
rect 72884 534006 72936 534012
rect 72896 531298 72924 534006
rect 72804 531270 72924 531298
rect 72804 524482 72832 531270
rect 72792 524476 72844 524482
rect 72792 524418 72844 524424
rect 72792 521688 72844 521694
rect 72792 521630 72844 521636
rect 72804 515642 72832 521630
rect 89640 515710 89668 699654
rect 106200 515778 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 644450 137968 654094
rect 154500 644450 154528 654094
rect 137756 644422 137968 644450
rect 154316 644422 154528 644450
rect 137756 634846 137784 644422
rect 154316 634846 154344 644422
rect 137744 634840 137796 634846
rect 137744 634782 137796 634788
rect 137928 634840 137980 634846
rect 137928 634782 137980 634788
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 137940 625138 137968 634782
rect 154500 625138 154528 634782
rect 137756 625110 137968 625138
rect 154316 625110 154528 625138
rect 137756 615534 137784 625110
rect 154316 615534 154344 625110
rect 137744 615528 137796 615534
rect 137744 615470 137796 615476
rect 137928 615528 137980 615534
rect 137928 615470 137980 615476
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 137940 605826 137968 615470
rect 154500 605826 154528 615470
rect 137756 605798 137968 605826
rect 154316 605798 154528 605826
rect 137756 596222 137784 605798
rect 154316 596222 154344 605798
rect 137744 596216 137796 596222
rect 137928 596216 137980 596222
rect 137744 596158 137796 596164
rect 137848 596164 137928 596170
rect 137848 596158 137980 596164
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 137848 596142 137968 596158
rect 154408 596142 154528 596158
rect 137848 591954 137876 596142
rect 154408 591954 154436 596142
rect 137756 591926 137876 591954
rect 154316 591926 154436 591954
rect 137756 589286 137784 591926
rect 154316 589286 154344 591926
rect 137744 589280 137796 589286
rect 137744 589222 137796 589228
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 137744 579760 137796 579766
rect 137664 579708 137744 579714
rect 154304 579760 154356 579766
rect 137664 579702 137796 579708
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 137664 579686 137784 579702
rect 154224 579686 154344 579702
rect 137664 579630 137692 579686
rect 154224 579630 154252 579686
rect 137652 579624 137704 579630
rect 137652 579566 137704 579572
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 137560 569968 137612 569974
rect 137560 569910 137612 569916
rect 129004 567860 129056 567866
rect 129004 567802 129056 567808
rect 106188 515772 106240 515778
rect 106188 515714 106240 515720
rect 89628 515704 89680 515710
rect 89628 515646 89680 515652
rect 72792 515636 72844 515642
rect 72792 515578 72844 515584
rect 41328 515568 41380 515574
rect 41328 515510 41380 515516
rect 24768 515500 24820 515506
rect 24768 515442 24820 515448
rect 128360 509244 128412 509250
rect 128360 509186 128412 509192
rect 128372 508609 128400 509186
rect 128358 508600 128414 508609
rect 128358 508535 128414 508544
rect 128360 502308 128412 502314
rect 128360 502250 128412 502256
rect 128372 500993 128400 502250
rect 128358 500984 128414 500993
rect 128358 500919 128414 500928
rect 128360 494012 128412 494018
rect 128360 493954 128412 493960
rect 128372 493377 128400 493954
rect 128358 493368 128414 493377
rect 128358 493303 128414 493312
rect 128360 485784 128412 485790
rect 128358 485752 128360 485761
rect 128412 485752 128414 485761
rect 128358 485687 128414 485696
rect 19984 478848 20036 478854
rect 19984 478790 20036 478796
rect 128360 478848 128412 478854
rect 128360 478790 128412 478796
rect 128372 478145 128400 478790
rect 128358 478136 128414 478145
rect 128358 478071 128414 478080
rect 129016 470529 129044 567802
rect 137572 563106 137600 569910
rect 137560 563100 137612 563106
rect 137560 563042 137612 563048
rect 154408 562970 154436 579566
rect 137652 562964 137704 562970
rect 137652 562906 137704 562912
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 137664 560250 137692 562906
rect 137652 560244 137704 560250
rect 137652 560186 137704 560192
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 137836 550656 137888 550662
rect 137836 550598 137888 550604
rect 137848 543658 137876 550598
rect 154316 550594 154344 553302
rect 154304 550588 154356 550594
rect 154304 550530 154356 550536
rect 154488 543788 154540 543794
rect 154488 543730 154540 543736
rect 137652 543652 137704 543658
rect 137652 543594 137704 543600
rect 137836 543652 137888 543658
rect 137836 543594 137888 543600
rect 137664 534070 137692 543594
rect 154500 540977 154528 543730
rect 154210 540968 154266 540977
rect 154210 540903 154266 540912
rect 154486 540968 154542 540977
rect 154486 540903 154542 540912
rect 137652 534064 137704 534070
rect 137652 534006 137704 534012
rect 137836 534064 137888 534070
rect 137836 534006 137888 534012
rect 137848 531298 137876 534006
rect 154224 531350 154252 540903
rect 137756 531270 137876 531298
rect 154212 531344 154264 531350
rect 154212 531286 154264 531292
rect 154304 531344 154356 531350
rect 154304 531286 154356 531292
rect 137756 524482 137784 531270
rect 154316 524482 154344 531286
rect 137744 524476 137796 524482
rect 137744 524418 137796 524424
rect 154304 524476 154356 524482
rect 154304 524418 154356 524424
rect 154396 524340 154448 524346
rect 154396 524282 154448 524288
rect 137744 521688 137796 521694
rect 137744 521630 137796 521636
rect 137756 518922 137784 521630
rect 137756 518894 137968 518922
rect 137940 515522 137968 518894
rect 137940 515494 138060 515522
rect 154408 515506 154436 524282
rect 171060 515574 171088 700198
rect 196808 515772 196860 515778
rect 196808 515714 196860 515720
rect 185032 515704 185084 515710
rect 185032 515646 185084 515652
rect 173256 515636 173308 515642
rect 173256 515578 173308 515584
rect 161480 515568 161532 515574
rect 161480 515510 161532 515516
rect 171048 515568 171100 515574
rect 171048 515510 171100 515516
rect 138032 515438 138060 515494
rect 149704 515500 149756 515506
rect 149704 515442 149756 515448
rect 154396 515500 154448 515506
rect 154396 515442 154448 515448
rect 137928 515432 137980 515438
rect 137928 515374 137980 515380
rect 138020 515432 138072 515438
rect 138020 515374 138072 515380
rect 137940 512380 137968 515374
rect 149716 512380 149744 515442
rect 161492 512380 161520 515510
rect 173268 512380 173296 515578
rect 185044 512380 185072 515646
rect 196820 512380 196848 515714
rect 202800 515642 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 218992 579630 219020 582354
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 218992 560250 219020 562906
rect 218980 560244 219032 560250
rect 218980 560186 219032 560192
rect 219164 550656 219216 550662
rect 219164 550598 219216 550604
rect 219176 543658 219204 550598
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 219164 543652 219216 543658
rect 219164 543594 219216 543600
rect 218992 534070 219020 543594
rect 218980 534064 219032 534070
rect 218980 534006 219032 534012
rect 219164 534064 219216 534070
rect 219164 534006 219216 534012
rect 219176 531298 219204 534006
rect 219084 531270 219204 531298
rect 219084 524482 219112 531270
rect 219072 524476 219124 524482
rect 219072 524418 219124 524424
rect 219072 521688 219124 521694
rect 219072 521630 219124 521636
rect 202788 515636 202840 515642
rect 202788 515578 202840 515584
rect 219084 515438 219112 521630
rect 232228 515568 232280 515574
rect 232228 515510 232280 515516
rect 220452 515500 220504 515506
rect 220452 515442 220504 515448
rect 208584 515432 208636 515438
rect 208584 515374 208636 515380
rect 219072 515432 219124 515438
rect 219072 515374 219124 515380
rect 208596 512380 208624 515374
rect 220464 512380 220492 515442
rect 232240 512380 232268 515510
rect 235920 515506 235948 699654
rect 244004 515636 244056 515642
rect 244004 515578 244056 515584
rect 235908 515500 235960 515506
rect 235908 515442 235960 515448
rect 244016 512380 244044 515578
rect 267556 515500 267608 515506
rect 267556 515442 267608 515448
rect 255780 515432 255832 515438
rect 255780 515374 255832 515380
rect 255792 512380 255820 515374
rect 267568 512380 267596 515442
rect 267660 515438 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654158 284064 663734
rect 284024 654152 284076 654158
rect 284024 654094 284076 654100
rect 284208 654152 284260 654158
rect 284208 654094 284260 654100
rect 284220 644450 284248 654094
rect 284036 644422 284248 644450
rect 284036 634846 284064 644422
rect 284024 634840 284076 634846
rect 284024 634782 284076 634788
rect 284208 634840 284260 634846
rect 284208 634782 284260 634788
rect 284220 625138 284248 634782
rect 284036 625110 284248 625138
rect 284036 615534 284064 625110
rect 284024 615528 284076 615534
rect 284024 615470 284076 615476
rect 284208 615528 284260 615534
rect 284208 615470 284260 615476
rect 284220 605826 284248 615470
rect 284036 605798 284248 605826
rect 284036 596222 284064 605798
rect 284024 596216 284076 596222
rect 284208 596216 284260 596222
rect 284024 596158 284076 596164
rect 284128 596164 284208 596170
rect 284128 596158 284260 596164
rect 284128 596142 284248 596158
rect 284128 591954 284156 596142
rect 284036 591926 284156 591954
rect 284036 589286 284064 591926
rect 284024 589280 284076 589286
rect 284024 589222 284076 589228
rect 284024 579760 284076 579766
rect 283944 579708 284024 579714
rect 283944 579702 284076 579708
rect 283944 579686 284064 579702
rect 283944 579630 283972 579686
rect 283932 579624 283984 579630
rect 283932 579566 283984 579572
rect 284116 579624 284168 579630
rect 284116 579566 284168 579572
rect 284128 562970 284156 579566
rect 283932 562964 283984 562970
rect 283932 562906 283984 562912
rect 284116 562964 284168 562970
rect 284116 562906 284168 562912
rect 283944 553330 283972 562906
rect 283944 553302 284064 553330
rect 284036 550594 284064 553302
rect 284024 550588 284076 550594
rect 284024 550530 284076 550536
rect 284208 543788 284260 543794
rect 284208 543730 284260 543736
rect 284220 540977 284248 543730
rect 284206 540968 284262 540977
rect 284206 540903 284262 540912
rect 284390 540968 284446 540977
rect 284390 540903 284446 540912
rect 284404 533882 284432 540903
rect 284128 533854 284432 533882
rect 284128 531321 284156 533854
rect 284114 531312 284170 531321
rect 284114 531247 284170 531256
rect 284298 531312 284354 531321
rect 284298 531247 284354 531256
rect 284312 524346 284340 531247
rect 284116 524340 284168 524346
rect 284116 524282 284168 524288
rect 284300 524340 284352 524346
rect 284300 524282 284352 524288
rect 284128 516118 284156 524282
rect 284116 516112 284168 516118
rect 284116 516054 284168 516060
rect 291108 516112 291160 516118
rect 291108 516054 291160 516060
rect 267648 515432 267700 515438
rect 267648 515374 267700 515380
rect 279332 515432 279384 515438
rect 279332 515374 279384 515380
rect 279344 512380 279372 515374
rect 291120 512380 291148 516054
rect 300780 514894 300808 699654
rect 332520 697610 332548 703520
rect 348804 703474 348832 703520
rect 364996 703474 365024 703520
rect 348804 703446 348924 703474
rect 364996 703446 365116 703474
rect 331220 697604 331272 697610
rect 331220 697546 331272 697552
rect 332508 697604 332560 697610
rect 332508 697546 332560 697552
rect 326528 515500 326580 515506
rect 326528 515442 326580 515448
rect 314752 515432 314804 515438
rect 314752 515374 314804 515380
rect 300768 514888 300820 514894
rect 300768 514830 300820 514836
rect 302976 514888 303028 514894
rect 302976 514830 303028 514836
rect 302988 512380 303016 514830
rect 314764 512380 314792 515374
rect 326540 512380 326568 515442
rect 331232 515438 331260 697546
rect 348896 692850 348924 703446
rect 365088 692850 365116 703446
rect 347780 692844 347832 692850
rect 347780 692786 347832 692792
rect 348884 692844 348936 692850
rect 348884 692786 348936 692792
rect 364340 692844 364392 692850
rect 364340 692786 364392 692792
rect 365076 692844 365128 692850
rect 365076 692786 365128 692792
rect 347792 683074 347820 692786
rect 364352 683074 364380 692786
rect 347792 683046 348004 683074
rect 364352 683046 364564 683074
rect 347976 673538 348004 683046
rect 364536 673538 364564 683046
rect 347780 673532 347832 673538
rect 347780 673474 347832 673480
rect 347964 673532 348016 673538
rect 347964 673474 348016 673480
rect 364340 673532 364392 673538
rect 364340 673474 364392 673480
rect 364524 673532 364576 673538
rect 364524 673474 364576 673480
rect 347792 663762 347820 673474
rect 364352 663762 364380 673474
rect 347792 663734 348004 663762
rect 364352 663734 364564 663762
rect 347976 654158 348004 663734
rect 364536 654158 364564 663734
rect 347780 654152 347832 654158
rect 347780 654094 347832 654100
rect 347964 654152 348016 654158
rect 347964 654094 348016 654100
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 347792 644450 347820 654094
rect 364352 644450 364380 654094
rect 347792 644422 348004 644450
rect 364352 644422 364564 644450
rect 347976 634846 348004 644422
rect 364536 634846 364564 644422
rect 347780 634840 347832 634846
rect 347780 634782 347832 634788
rect 347964 634840 348016 634846
rect 347964 634782 348016 634788
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 347792 625138 347820 634782
rect 364352 625138 364380 634782
rect 347792 625110 348004 625138
rect 364352 625110 364564 625138
rect 347976 615534 348004 625110
rect 364536 615534 364564 625110
rect 347780 615528 347832 615534
rect 347780 615470 347832 615476
rect 347964 615528 348016 615534
rect 347964 615470 348016 615476
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 347792 605826 347820 615470
rect 364352 605826 364380 615470
rect 347792 605798 348004 605826
rect 364352 605798 364564 605826
rect 347976 596222 348004 605798
rect 364536 596222 364564 605798
rect 347780 596216 347832 596222
rect 347964 596216 348016 596222
rect 347832 596164 347912 596170
rect 347780 596158 347912 596164
rect 347964 596158 348016 596164
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 347792 596142 347912 596158
rect 364352 596142 364472 596158
rect 347884 596034 347912 596142
rect 364444 596034 364472 596142
rect 347884 596006 348004 596034
rect 364444 596006 364564 596034
rect 347976 591954 348004 596006
rect 364536 591954 364564 596006
rect 347884 591926 348004 591954
rect 364444 591926 364564 591954
rect 347884 589286 347912 591926
rect 364444 589286 364472 591926
rect 347872 589280 347924 589286
rect 347872 589222 347924 589228
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 347780 579692 347832 579698
rect 347780 579634 347832 579640
rect 364340 579692 364392 579698
rect 364340 579634 364392 579640
rect 347792 572642 347820 579634
rect 364352 572642 364380 579634
rect 347792 572614 347912 572642
rect 364352 572614 364472 572642
rect 347884 569906 347912 572614
rect 364444 569906 364472 572614
rect 347872 569900 347924 569906
rect 347872 569842 347924 569848
rect 364432 569900 364484 569906
rect 364432 569842 364484 569848
rect 348056 563100 348108 563106
rect 348056 563042 348108 563048
rect 364616 563100 364668 563106
rect 364616 563042 364668 563048
rect 348068 560289 348096 563042
rect 364628 560289 364656 563042
rect 347870 560280 347926 560289
rect 347870 560215 347926 560224
rect 348054 560280 348110 560289
rect 348054 560215 348110 560224
rect 364430 560280 364486 560289
rect 364430 560215 364486 560224
rect 364614 560280 364670 560289
rect 364614 560215 364670 560224
rect 347884 550662 347912 560215
rect 364444 550662 364472 560215
rect 347872 550656 347924 550662
rect 347872 550598 347924 550604
rect 348148 550656 348200 550662
rect 348148 550598 348200 550604
rect 364432 550656 364484 550662
rect 364432 550598 364484 550604
rect 364708 550656 364760 550662
rect 364708 550598 364760 550604
rect 348160 543862 348188 550598
rect 364720 543862 364748 550598
rect 348148 543856 348200 543862
rect 348148 543798 348200 543804
rect 364708 543856 364760 543862
rect 364708 543798 364760 543804
rect 348056 543720 348108 543726
rect 348056 543662 348108 543668
rect 364616 543720 364668 543726
rect 364616 543662 364668 543668
rect 348068 540977 348096 543662
rect 364628 540977 364656 543662
rect 347870 540968 347926 540977
rect 347870 540903 347926 540912
rect 348054 540968 348110 540977
rect 348054 540903 348110 540912
rect 364430 540968 364486 540977
rect 364430 540903 364486 540912
rect 364614 540968 364670 540977
rect 364614 540903 364670 540912
rect 347884 531350 347912 540903
rect 364444 531350 364472 540903
rect 347872 531344 347924 531350
rect 347872 531286 347924 531292
rect 348148 531344 348200 531350
rect 348148 531286 348200 531292
rect 364432 531344 364484 531350
rect 364432 531286 364484 531292
rect 364708 531344 364760 531350
rect 364708 531286 364760 531292
rect 348160 521694 348188 531286
rect 364720 521694 364748 531286
rect 347964 521688 348016 521694
rect 347964 521630 348016 521636
rect 348148 521688 348200 521694
rect 348148 521630 348200 521636
rect 364524 521688 364576 521694
rect 364524 521630 364576 521636
rect 364708 521688 364760 521694
rect 364708 521630 364760 521636
rect 347976 515506 348004 521630
rect 350080 515568 350132 515574
rect 350080 515510 350132 515516
rect 347964 515500 348016 515506
rect 347964 515442 348016 515448
rect 331220 515432 331272 515438
rect 331220 515374 331272 515380
rect 338304 515432 338356 515438
rect 338304 515374 338356 515380
rect 338316 512380 338344 515374
rect 350092 512380 350120 515510
rect 361856 515500 361908 515506
rect 361856 515442 361908 515448
rect 361868 512380 361896 515442
rect 364536 515438 364564 521630
rect 385500 515772 385552 515778
rect 385500 515714 385552 515720
rect 364524 515432 364576 515438
rect 364524 515374 364576 515380
rect 373632 515432 373684 515438
rect 373632 515374 373684 515380
rect 373644 512380 373672 515374
rect 385512 512380 385540 515714
rect 397276 515704 397328 515710
rect 397276 515646 397328 515652
rect 397288 512380 397316 515646
rect 397472 515574 397500 703520
rect 413664 703474 413692 703520
rect 413664 703446 413784 703474
rect 413756 698290 413784 703446
rect 413008 698284 413060 698290
rect 413008 698226 413060 698232
rect 413744 698284 413796 698290
rect 413744 698226 413796 698232
rect 413020 694142 413048 698226
rect 412824 694136 412876 694142
rect 412824 694078 412876 694084
rect 413008 694136 413060 694142
rect 413008 694078 413060 694084
rect 412836 692782 412864 694078
rect 412824 692776 412876 692782
rect 412824 692718 412876 692724
rect 429856 684486 429884 703520
rect 429200 684480 429252 684486
rect 429200 684422 429252 684428
rect 429844 684480 429896 684486
rect 429844 684422 429896 684428
rect 412640 683256 412692 683262
rect 412640 683198 412692 683204
rect 412652 683126 412680 683198
rect 429212 683126 429240 684422
rect 412640 683120 412692 683126
rect 412640 683062 412692 683068
rect 429200 683120 429252 683126
rect 429200 683062 429252 683068
rect 413100 666596 413152 666602
rect 413100 666538 413152 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 413112 659682 413140 666538
rect 429672 659682 429700 666538
rect 412928 659654 413140 659682
rect 429488 659654 429700 659682
rect 412928 647290 412956 659654
rect 429488 647290 429516 659654
rect 412824 647284 412876 647290
rect 412824 647226 412876 647232
rect 412916 647284 412968 647290
rect 412916 647226 412968 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 412836 640422 412864 647226
rect 429396 640422 429424 647226
rect 412824 640416 412876 640422
rect 412824 640358 412876 640364
rect 412916 640416 412968 640422
rect 412916 640358 412968 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 412928 630698 412956 640358
rect 429488 630698 429516 640358
rect 412732 630692 412784 630698
rect 412732 630634 412784 630640
rect 412916 630692 412968 630698
rect 412916 630634 412968 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 412744 630578 412772 630634
rect 429304 630578 429332 630634
rect 412744 630550 412864 630578
rect 429304 630550 429424 630578
rect 412836 621058 412864 630550
rect 429396 621058 429424 630550
rect 412836 621030 412956 621058
rect 429396 621030 429516 621058
rect 412928 611386 412956 621030
rect 429488 611386 429516 621030
rect 412732 611380 412784 611386
rect 412732 611322 412784 611328
rect 412916 611380 412968 611386
rect 412916 611322 412968 611328
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 412744 611266 412772 611322
rect 429304 611266 429332 611322
rect 412744 611238 412864 611266
rect 429304 611238 429424 611266
rect 412836 608598 412864 611238
rect 429396 608598 429424 611238
rect 412824 608592 412876 608598
rect 412824 608534 412876 608540
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 413008 601724 413060 601730
rect 413008 601666 413060 601672
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 413020 598942 413048 601666
rect 429580 598942 429608 601666
rect 413008 598936 413060 598942
rect 413008 598878 413060 598884
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 413100 589348 413152 589354
rect 413100 589290 413152 589296
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 413112 582486 413140 589290
rect 429672 582486 429700 589290
rect 413100 582480 413152 582486
rect 413100 582422 413152 582428
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 413008 582344 413060 582350
rect 413008 582286 413060 582292
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 413020 572642 413048 582286
rect 429580 572642 429608 582286
rect 412836 572614 413048 572642
rect 429396 572614 429608 572642
rect 412836 569922 412864 572614
rect 429396 569922 429424 572614
rect 412744 569894 412864 569922
rect 429304 569894 429424 569922
rect 412744 563174 412772 569894
rect 429304 563174 429332 569894
rect 412732 563168 412784 563174
rect 412732 563110 412784 563116
rect 429292 563168 429344 563174
rect 429292 563110 429344 563116
rect 412732 563032 412784 563038
rect 412732 562974 412784 562980
rect 429292 563032 429344 563038
rect 429292 562974 429344 562980
rect 412744 560250 412772 562974
rect 429304 560250 429332 562974
rect 412732 560244 412784 560250
rect 412732 560186 412784 560192
rect 429292 560244 429344 560250
rect 429292 560186 429344 560192
rect 412916 550656 412968 550662
rect 412916 550598 412968 550604
rect 429476 550656 429528 550662
rect 429476 550598 429528 550604
rect 412928 543658 412956 550598
rect 429488 543658 429516 550598
rect 412732 543652 412784 543658
rect 412732 543594 412784 543600
rect 412916 543652 412968 543658
rect 412916 543594 412968 543600
rect 429292 543652 429344 543658
rect 429292 543594 429344 543600
rect 429476 543652 429528 543658
rect 429476 543594 429528 543600
rect 412744 534018 412772 543594
rect 429304 534018 429332 543594
rect 412744 533990 412864 534018
rect 429304 533990 429424 534018
rect 412836 524498 412864 533990
rect 429396 524498 429424 533990
rect 412836 524470 412956 524498
rect 429396 524470 429516 524498
rect 409052 515636 409104 515642
rect 409052 515578 409104 515584
rect 397460 515568 397512 515574
rect 397460 515510 397512 515516
rect 409064 512380 409092 515578
rect 412928 515506 412956 524470
rect 420828 515568 420880 515574
rect 420828 515510 420880 515516
rect 412916 515500 412968 515506
rect 412916 515442 412968 515448
rect 420840 512380 420868 515510
rect 429488 515438 429516 524470
rect 462332 515778 462360 703520
rect 478524 703474 478552 703520
rect 494808 703474 494836 703520
rect 478524 703446 478644 703474
rect 494808 703446 494928 703474
rect 472624 696992 472676 696998
rect 472624 696934 472676 696940
rect 471244 650072 471296 650078
rect 471244 650014 471296 650020
rect 467104 603152 467156 603158
rect 467104 603094 467156 603100
rect 462320 515772 462372 515778
rect 462320 515714 462372 515720
rect 432604 515500 432656 515506
rect 432604 515442 432656 515448
rect 429476 515432 429528 515438
rect 429476 515374 429528 515380
rect 432616 512380 432644 515442
rect 444380 515432 444432 515438
rect 444380 515374 444432 515380
rect 444392 512380 444420 515374
rect 462964 509312 463016 509318
rect 462964 509254 463016 509260
rect 453212 509244 453264 509250
rect 453212 509186 453264 509192
rect 453224 508881 453252 509186
rect 453210 508872 453266 508881
rect 453210 508807 453266 508816
rect 453396 502308 453448 502314
rect 453396 502250 453448 502256
rect 453408 501809 453436 502250
rect 453394 501800 453450 501809
rect 453394 501735 453450 501744
rect 460204 498228 460256 498234
rect 460204 498170 460256 498176
rect 453948 495440 454000 495446
rect 453948 495382 454000 495388
rect 453960 494601 453988 495382
rect 453946 494592 454002 494601
rect 453946 494527 454002 494536
rect 453764 488504 453816 488510
rect 453764 488446 453816 488452
rect 453776 487529 453804 488446
rect 453762 487520 453818 487529
rect 453762 487455 453818 487464
rect 456064 485852 456116 485858
rect 456064 485794 456116 485800
rect 453764 481636 453816 481642
rect 453764 481578 453816 481584
rect 453776 480457 453804 481578
rect 453762 480448 453818 480457
rect 453762 480383 453818 480392
rect 453948 473340 454000 473346
rect 453948 473282 454000 473288
rect 453960 473249 453988 473282
rect 453946 473240 454002 473249
rect 453946 473175 454002 473184
rect 129002 470520 129058 470529
rect 129002 470455 129058 470464
rect 452752 466404 452804 466410
rect 452752 466346 452804 466352
rect 452764 466177 452792 466346
rect 452750 466168 452806 466177
rect 452750 466103 452806 466112
rect 128360 463684 128412 463690
rect 128360 463626 128412 463632
rect 128372 462913 128400 463626
rect 128358 462904 128414 462913
rect 128358 462839 128414 462848
rect 454684 462392 454736 462398
rect 454684 462334 454736 462340
rect 453396 459536 453448 459542
rect 453396 459478 453448 459484
rect 453408 459105 453436 459478
rect 453394 459096 453450 459105
rect 453394 459031 453450 459040
rect 128360 455388 128412 455394
rect 128360 455330 128412 455336
rect 128372 455297 128400 455330
rect 128358 455288 128414 455297
rect 128358 455223 128414 455232
rect 453948 452600 454000 452606
rect 453948 452542 454000 452548
rect 453960 451897 453988 452542
rect 453946 451888 454002 451897
rect 453946 451823 454002 451832
rect 58624 451308 58676 451314
rect 58624 451250 58676 451256
rect 15844 448520 15896 448526
rect 15844 448462 15896 448468
rect 13084 440224 13136 440230
rect 13084 440166 13136 440172
rect 8944 425060 8996 425066
rect 8944 425002 8996 425008
rect 3514 423736 3570 423745
rect 3514 423671 3570 423680
rect 3424 409828 3476 409834
rect 3424 409770 3476 409776
rect 3528 402966 3556 423671
rect 58636 418130 58664 451250
rect 128360 448520 128412 448526
rect 128360 448462 128412 448468
rect 128372 447681 128400 448462
rect 128358 447672 128414 447681
rect 128358 447607 128414 447616
rect 453672 445732 453724 445738
rect 453672 445674 453724 445680
rect 453684 444825 453712 445674
rect 453670 444816 453726 444825
rect 453670 444751 453726 444760
rect 128360 440224 128412 440230
rect 128360 440166 128412 440172
rect 128372 440065 128400 440166
rect 128358 440056 128414 440065
rect 128358 439991 128414 440000
rect 453304 438932 453356 438938
rect 453304 438874 453356 438880
rect 128360 433288 128412 433294
rect 128360 433230 128412 433236
rect 128372 432313 128400 433230
rect 128358 432304 128414 432313
rect 128358 432239 128414 432248
rect 128360 425060 128412 425066
rect 128360 425002 128412 425008
rect 128372 424697 128400 425002
rect 128358 424688 128414 424697
rect 128358 424623 128414 424632
rect 58624 418124 58676 418130
rect 58624 418066 58676 418072
rect 128360 418124 128412 418130
rect 128360 418066 128412 418072
rect 128372 417081 128400 418066
rect 128358 417072 128414 417081
rect 128358 417007 128414 417016
rect 128360 409828 128412 409834
rect 128360 409770 128412 409776
rect 128372 409465 128400 409770
rect 128358 409456 128414 409465
rect 128358 409391 128414 409400
rect 3516 402960 3568 402966
rect 3516 402902 3568 402908
rect 128360 402960 128412 402966
rect 128360 402902 128412 402908
rect 128372 401849 128400 402902
rect 452844 402552 452896 402558
rect 452844 402494 452896 402500
rect 452856 402121 452884 402494
rect 452842 402112 452898 402121
rect 452842 402047 452898 402056
rect 128358 401840 128414 401849
rect 128358 401775 128414 401784
rect 3422 395040 3478 395049
rect 3422 394975 3478 394984
rect 3436 394670 3464 394975
rect 3424 394664 3476 394670
rect 3424 394606 3476 394612
rect 128360 394664 128412 394670
rect 128360 394606 128412 394612
rect 128372 394233 128400 394606
rect 128358 394224 128414 394233
rect 128358 394159 128414 394168
rect 453316 387841 453344 438874
rect 453764 438864 453816 438870
rect 453764 438806 453816 438812
rect 453776 437753 453804 438806
rect 453762 437744 453818 437753
rect 453762 437679 453818 437688
rect 453948 430568 454000 430574
rect 453946 430536 453948 430545
rect 454000 430536 454002 430545
rect 453946 430471 454002 430480
rect 453948 423632 454000 423638
rect 453948 423574 454000 423580
rect 453960 423473 453988 423574
rect 453946 423464 454002 423473
rect 453946 423399 454002 423408
rect 453948 416424 454000 416430
rect 453946 416392 453948 416401
rect 454000 416392 454002 416401
rect 453946 416327 454002 416336
rect 453396 409420 453448 409426
rect 453396 409362 453448 409368
rect 453408 409193 453436 409362
rect 453394 409184 453450 409193
rect 453394 409119 453450 409128
rect 454696 402558 454724 462334
rect 456076 409426 456104 485794
rect 460216 416430 460244 498170
rect 462976 423638 463004 509254
rect 467116 466410 467144 603094
rect 471256 488510 471284 650014
rect 472636 509250 472664 696934
rect 478616 692850 478644 703446
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 477512 683074 477540 692786
rect 494900 685914 494928 703446
rect 494244 685908 494296 685914
rect 494244 685850 494296 685856
rect 494888 685908 494940 685914
rect 494888 685850 494940 685856
rect 477512 683046 477724 683074
rect 477696 673538 477724 683046
rect 494256 678994 494284 685850
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 490564 673532 490616 673538
rect 490564 673474 490616 673480
rect 477512 663762 477540 673474
rect 477512 663734 477724 663762
rect 477696 654158 477724 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 477512 644450 477540 654094
rect 477512 644422 477724 644450
rect 477696 634846 477724 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 477512 625138 477540 634782
rect 479524 626612 479576 626618
rect 479524 626554 479576 626560
rect 477512 625110 477724 625138
rect 477696 615534 477724 625110
rect 477500 615528 477552 615534
rect 477500 615470 477552 615476
rect 477684 615528 477736 615534
rect 477684 615470 477736 615476
rect 477512 605826 477540 615470
rect 477512 605798 477724 605826
rect 477696 596222 477724 605798
rect 477500 596216 477552 596222
rect 477684 596216 477736 596222
rect 477552 596164 477632 596170
rect 477500 596158 477632 596164
rect 477684 596158 477736 596164
rect 477512 596142 477632 596158
rect 477604 596034 477632 596142
rect 477604 596006 477724 596034
rect 476764 592068 476816 592074
rect 476764 592010 476816 592016
rect 475384 545148 475436 545154
rect 475384 545090 475436 545096
rect 472624 509244 472676 509250
rect 472624 509186 472676 509192
rect 471244 488504 471296 488510
rect 471244 488446 471296 488452
rect 467104 466404 467156 466410
rect 467104 466346 467156 466352
rect 475396 438870 475424 545090
rect 476776 459542 476804 592010
rect 477696 591954 477724 596006
rect 477604 591926 477724 591954
rect 477604 589286 477632 591926
rect 477592 589280 477644 589286
rect 477592 589222 477644 589228
rect 477500 579692 477552 579698
rect 477500 579634 477552 579640
rect 477512 572642 477540 579634
rect 477512 572614 477632 572642
rect 477604 569906 477632 572614
rect 477592 569900 477644 569906
rect 477592 569842 477644 569848
rect 477776 563100 477828 563106
rect 477776 563042 477828 563048
rect 477788 560289 477816 563042
rect 477590 560280 477646 560289
rect 477590 560215 477646 560224
rect 477774 560280 477830 560289
rect 477774 560215 477830 560224
rect 477604 550662 477632 560215
rect 477592 550656 477644 550662
rect 477592 550598 477644 550604
rect 477868 550656 477920 550662
rect 477868 550598 477920 550604
rect 477880 543862 477908 550598
rect 477868 543856 477920 543862
rect 477868 543798 477920 543804
rect 477776 543720 477828 543726
rect 477776 543662 477828 543668
rect 477788 540977 477816 543662
rect 477590 540968 477646 540977
rect 477590 540903 477646 540912
rect 477774 540968 477830 540977
rect 477774 540903 477830 540912
rect 477604 531350 477632 540903
rect 477592 531344 477644 531350
rect 477592 531286 477644 531292
rect 477868 531344 477920 531350
rect 477868 531286 477920 531292
rect 477880 521694 477908 531286
rect 477684 521688 477736 521694
rect 477684 521630 477736 521636
rect 477868 521688 477920 521694
rect 477868 521630 477920 521636
rect 477696 515710 477724 521630
rect 477684 515704 477736 515710
rect 477684 515646 477736 515652
rect 479536 473346 479564 626554
rect 489184 579692 489236 579698
rect 489184 579634 489236 579640
rect 483664 556232 483716 556238
rect 483664 556174 483716 556180
rect 479524 473340 479576 473346
rect 479524 473282 479576 473288
rect 476764 459536 476816 459542
rect 476764 459478 476816 459484
rect 483676 445738 483704 556174
rect 485044 532772 485096 532778
rect 485044 532714 485096 532720
rect 483664 445732 483716 445738
rect 483664 445674 483716 445680
rect 475384 438864 475436 438870
rect 475384 438806 475436 438812
rect 485056 430574 485084 532714
rect 489196 452606 489224 579634
rect 490576 495446 490604 673474
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 494164 659682 494192 666538
rect 494164 659654 494284 659682
rect 494256 654158 494284 659654
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 494072 644450 494100 654094
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 494072 625110 494284 625138
rect 494256 615534 494284 625110
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 494072 605826 494100 615470
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579737 493916 589222
rect 493874 579728 493930 579737
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 494072 572642 494100 579663
rect 494072 572614 494192 572642
rect 494164 569906 494192 572614
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 494348 560289 494376 563042
rect 494150 560280 494206 560289
rect 494150 560215 494206 560224
rect 494334 560280 494390 560289
rect 494334 560215 494390 560224
rect 494164 550662 494192 560215
rect 494152 550656 494204 550662
rect 494152 550598 494204 550604
rect 494428 550656 494480 550662
rect 494428 550598 494480 550604
rect 494440 543862 494468 550598
rect 494428 543856 494480 543862
rect 494428 543798 494480 543804
rect 494336 543720 494388 543726
rect 494336 543662 494388 543668
rect 494348 540977 494376 543662
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 494164 531350 494192 540903
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 494440 521694 494468 531286
rect 494244 521688 494296 521694
rect 494244 521630 494296 521636
rect 494428 521688 494480 521694
rect 494428 521630 494480 521636
rect 494256 515642 494284 521630
rect 494244 515636 494296 515642
rect 494244 515578 494296 515584
rect 527192 515574 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 694142 542768 698226
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 692782 542584 694078
rect 542544 692776 542596 692782
rect 542544 692718 542596 692724
rect 542728 692776 542780 692782
rect 542728 692718 542780 692724
rect 542740 683233 542768 692718
rect 559668 684486 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 558920 684480 558972 684486
rect 558920 684422 558972 684428
rect 559656 684480 559708 684486
rect 559656 684422 559708 684428
rect 542358 683224 542414 683233
rect 542358 683159 542414 683168
rect 542726 683224 542782 683233
rect 542726 683159 542782 683168
rect 542372 683126 542400 683159
rect 558932 683126 558960 684422
rect 542360 683120 542412 683126
rect 542360 683062 542412 683068
rect 558920 683120 558972 683126
rect 558920 683062 558972 683068
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 542832 659682 542860 666538
rect 559392 659682 559420 666538
rect 542648 659654 542860 659682
rect 559208 659654 559420 659682
rect 542648 647290 542676 659654
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 542556 640422 542584 647226
rect 559116 640422 559144 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 542648 630698 542676 640358
rect 559208 630698 559236 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 542464 630578 542492 630634
rect 559024 630578 559052 630634
rect 542464 630550 542584 630578
rect 559024 630550 559144 630578
rect 542556 621058 542584 630550
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 559116 621030 559236 621058
rect 542648 611386 542676 621030
rect 559208 611386 559236 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 542464 611266 542492 611322
rect 559024 611266 559052 611322
rect 542464 611238 542584 611266
rect 559024 611238 559144 611266
rect 542556 608598 542584 611238
rect 559116 608598 559144 611238
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 542740 598942 542768 601666
rect 559300 598942 559328 601666
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 579894 592512 579950 592521
rect 579894 592447 579950 592456
rect 579908 592074 579936 592447
rect 579896 592068 579948 592074
rect 579896 592010 579948 592016
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 542832 582486 542860 589290
rect 559392 582486 559420 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 542740 572642 542768 582286
rect 559300 572642 559328 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 542556 572614 542768 572642
rect 559116 572614 559328 572642
rect 542556 569922 542584 572614
rect 559116 569922 559144 572614
rect 542464 569894 542584 569922
rect 559024 569894 559144 569922
rect 542464 563174 542492 569894
rect 559024 563174 559052 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 542464 560250 542492 562974
rect 559024 560250 559052 562974
rect 542452 560244 542504 560250
rect 542452 560186 542504 560192
rect 559012 560244 559064 560250
rect 559012 560186 559064 560192
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 542636 550656 542688 550662
rect 542636 550598 542688 550604
rect 559196 550656 559248 550662
rect 559196 550598 559248 550604
rect 542648 543658 542676 550598
rect 559208 543658 559236 550598
rect 579894 545592 579950 545601
rect 579894 545527 579950 545536
rect 579908 545154 579936 545527
rect 579896 545148 579948 545154
rect 579896 545090 579948 545096
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542636 543652 542688 543658
rect 542636 543594 542688 543600
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559196 543652 559248 543658
rect 559196 543594 559248 543600
rect 542464 534018 542492 543594
rect 559024 534018 559052 543594
rect 542464 533990 542584 534018
rect 559024 533990 559144 534018
rect 542556 524498 542584 533990
rect 559116 524498 559144 533990
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 542556 524470 542676 524498
rect 559116 524470 559236 524498
rect 527180 515568 527232 515574
rect 527180 515510 527232 515516
rect 542648 515506 542676 524470
rect 542636 515500 542688 515506
rect 542636 515442 542688 515448
rect 559208 515438 559236 524470
rect 559196 515432 559248 515438
rect 559196 515374 559248 515380
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580276 502314 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580264 502308 580316 502314
rect 580264 502250 580316 502256
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 490564 495440 490616 495446
rect 490564 495382 490616 495388
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580368 481642 580396 639367
rect 580356 481636 580408 481642
rect 580356 481578 580408 481584
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 489184 452600 489236 452606
rect 489184 452542 489236 452548
rect 580262 451752 580318 451761
rect 580262 451687 580318 451696
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 579908 438938 579936 439855
rect 579896 438932 579948 438938
rect 579896 438874 579948 438880
rect 485044 430568 485096 430574
rect 485044 430510 485096 430516
rect 462964 423632 463016 423638
rect 462964 423574 463016 423580
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 460204 416424 460256 416430
rect 460204 416366 460256 416372
rect 580184 414730 580212 416463
rect 543004 414724 543056 414730
rect 543004 414666 543056 414672
rect 580172 414724 580224 414730
rect 580172 414666 580224 414672
rect 456064 409420 456116 409426
rect 456064 409362 456116 409368
rect 454684 402552 454736 402558
rect 454684 402494 454736 402500
rect 453764 396024 453816 396030
rect 453764 395966 453816 395972
rect 453776 394913 453804 395966
rect 453762 394904 453818 394913
rect 453762 394839 453818 394848
rect 454684 392012 454736 392018
rect 454684 391954 454736 391960
rect 453302 387832 453358 387841
rect 453302 387767 453358 387776
rect 129002 386608 129058 386617
rect 129002 386543 129058 386552
rect 129016 380866 129044 386543
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 129004 380860 129056 380866
rect 129004 380802 129056 380808
rect 453948 380860 454000 380866
rect 453948 380802 454000 380808
rect 3252 380633 3280 380802
rect 453960 380769 453988 380802
rect 453946 380760 454002 380769
rect 453946 380695 454002 380704
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 129002 378992 129058 379001
rect 129002 378927 129058 378936
rect 129016 367062 129044 378927
rect 453396 373992 453448 373998
rect 453396 373934 453448 373940
rect 453408 373561 453436 373934
rect 453394 373552 453450 373561
rect 453394 373487 453450 373496
rect 129278 371376 129334 371385
rect 129278 371311 129334 371320
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 129004 367056 129056 367062
rect 129004 366998 129056 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 129002 363760 129058 363769
rect 129002 363695 129058 363704
rect 128358 348392 128414 348401
rect 128358 348327 128414 348336
rect 128372 347818 128400 348327
rect 8944 347812 8996 347818
rect 8944 347754 8996 347760
rect 128360 347812 128412 347818
rect 128360 347754 128412 347760
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 8956 294914 8984 347754
rect 128358 333160 128414 333169
rect 128358 333095 128414 333104
rect 128372 332654 128400 333095
rect 13084 332648 13136 332654
rect 13084 332590 13136 332596
rect 128360 332648 128412 332654
rect 128360 332590 128412 332596
rect 11704 324352 11756 324358
rect 11704 324294 11756 324300
rect 10324 302252 10376 302258
rect 10324 302194 10376 302200
rect 3516 294908 3568 294914
rect 3516 294850 3568 294856
rect 8944 294908 8996 294914
rect 8944 294850 8996 294856
rect 3528 294409 3556 294850
rect 3514 294400 3570 294409
rect 3514 294335 3570 294344
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 3148 266348 3200 266354
rect 3148 266290 3200 266296
rect 3160 265713 3188 266290
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 8944 233300 8996 233306
rect 8944 233242 8996 233248
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 8956 79490 8984 233242
rect 10336 208350 10364 302194
rect 11716 252550 11744 324294
rect 13096 266354 13124 332590
rect 128358 325544 128414 325553
rect 128358 325479 128414 325488
rect 128372 324358 128400 325479
rect 128360 324352 128412 324358
rect 128360 324294 128412 324300
rect 129016 324290 129044 363695
rect 129186 356144 129242 356153
rect 129186 356079 129242 356088
rect 129094 340776 129150 340785
rect 129094 340711 129150 340720
rect 129004 324284 129056 324290
rect 129004 324226 129056 324232
rect 129002 317928 129058 317937
rect 129002 317863 129058 317872
rect 128358 310312 128414 310321
rect 128358 310247 128414 310256
rect 128372 309194 128400 310247
rect 15844 309188 15896 309194
rect 15844 309130 15896 309136
rect 128360 309188 128412 309194
rect 128360 309130 128412 309136
rect 13084 266348 13136 266354
rect 13084 266290 13136 266296
rect 13084 263628 13136 263634
rect 13084 263570 13136 263576
rect 11704 252544 11756 252550
rect 11704 252486 11756 252492
rect 11704 211200 11756 211206
rect 11704 211142 11756 211148
rect 10324 208344 10376 208350
rect 10324 208286 10376 208292
rect 10324 194608 10376 194614
rect 10324 194550 10376 194556
rect 3516 79484 3568 79490
rect 3516 79426 3568 79432
rect 8944 79484 8996 79490
rect 8944 79426 8996 79432
rect 3528 78985 3556 79426
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 10336 8294 10364 194550
rect 11716 35902 11744 211142
rect 13096 136610 13124 263570
rect 14464 256760 14516 256766
rect 14464 256702 14516 256708
rect 13084 136604 13136 136610
rect 13084 136546 13136 136552
rect 14476 122806 14504 256702
rect 15856 223582 15884 309130
rect 128358 302696 128414 302705
rect 128358 302631 128414 302640
rect 128372 302258 128400 302631
rect 128360 302252 128412 302258
rect 128360 302194 128412 302200
rect 128358 287464 128414 287473
rect 128358 287399 128414 287408
rect 128372 287094 128400 287399
rect 17224 287088 17276 287094
rect 17224 287030 17276 287036
rect 128360 287088 128412 287094
rect 128360 287030 128412 287036
rect 15844 223576 15896 223582
rect 15844 223518 15896 223524
rect 15844 218068 15896 218074
rect 15844 218010 15896 218016
rect 14464 122800 14516 122806
rect 14464 122742 14516 122748
rect 15856 51066 15884 218010
rect 17236 180810 17264 287030
rect 126244 278792 126296 278798
rect 126244 278734 126296 278740
rect 19984 241528 20036 241534
rect 19984 241470 20036 241476
rect 17224 180804 17276 180810
rect 17224 180746 17276 180752
rect 19996 93838 20024 241470
rect 126256 165578 126284 278734
rect 128358 264480 128414 264489
rect 128358 264415 128414 264424
rect 128372 263634 128400 264415
rect 128360 263628 128412 263634
rect 128360 263570 128412 263576
rect 128358 256864 128414 256873
rect 128358 256799 128414 256808
rect 128372 256766 128400 256799
rect 128360 256760 128412 256766
rect 128360 256702 128412 256708
rect 128358 241632 128414 241641
rect 128358 241567 128414 241576
rect 128372 241534 128400 241567
rect 128360 241528 128412 241534
rect 128360 241470 128412 241476
rect 129016 237386 129044 317863
rect 129108 280158 129136 340711
rect 129200 309126 129228 356079
rect 129292 338094 129320 371311
rect 454696 367062 454724 391954
rect 543016 380866 543044 414666
rect 580276 396030 580304 451687
rect 580354 404832 580410 404841
rect 580354 404767 580410 404776
rect 580264 396024 580316 396030
rect 580264 395966 580316 395972
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 543004 380860 543056 380866
rect 543004 380802 543056 380808
rect 580368 373998 580396 404767
rect 580356 373992 580408 373998
rect 580356 373934 580408 373940
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 452660 367056 452712 367062
rect 452660 366998 452712 367004
rect 454684 367056 454736 367062
rect 454684 366998 454736 367004
rect 452672 366489 452700 366998
rect 452658 366480 452714 366489
rect 452658 366415 452714 366424
rect 580276 360194 580304 369543
rect 453948 360188 454000 360194
rect 453948 360130 454000 360136
rect 580264 360188 580316 360194
rect 580264 360130 580316 360136
rect 453960 359417 453988 360130
rect 453946 359408 454002 359417
rect 453946 359343 454002 359352
rect 580262 357912 580318 357921
rect 580262 357847 580318 357856
rect 580276 353258 580304 357847
rect 453764 353252 453816 353258
rect 453764 353194 453816 353200
rect 580264 353252 580316 353258
rect 580264 353194 580316 353200
rect 453776 352209 453804 353194
rect 453762 352200 453818 352209
rect 453762 352135 453818 352144
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345710 580212 346015
rect 453948 345704 454000 345710
rect 453948 345646 454000 345652
rect 580172 345704 580224 345710
rect 580172 345646 580224 345652
rect 453960 345137 453988 345646
rect 453946 345128 454002 345137
rect 453946 345063 454002 345072
rect 129280 338088 129332 338094
rect 129280 338030 129332 338036
rect 453486 338056 453542 338065
rect 453486 337991 453542 338000
rect 453394 330848 453450 330857
rect 453394 330783 453450 330792
rect 453302 323776 453358 323785
rect 453302 323711 453358 323720
rect 129188 309120 129240 309126
rect 129188 309062 129240 309068
rect 452934 302424 452990 302433
rect 452934 302359 452936 302368
rect 452988 302359 452990 302368
rect 452936 302330 452988 302336
rect 453316 299470 453344 323711
rect 453408 311846 453436 330783
rect 453500 322930 453528 337991
rect 453488 322924 453540 322930
rect 453488 322866 453540 322872
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 453578 316704 453634 316713
rect 453578 316639 453634 316648
rect 453396 311840 453448 311846
rect 453396 311782 453448 311788
rect 453486 309496 453542 309505
rect 453486 309431 453542 309440
rect 453304 299464 453356 299470
rect 453304 299406 453356 299412
rect 453394 295216 453450 295225
rect 453394 295151 453450 295160
rect 129370 295080 129426 295089
rect 129370 295015 129426 295024
rect 129096 280152 129148 280158
rect 129096 280094 129148 280100
rect 129094 279848 129150 279857
rect 129094 279783 129150 279792
rect 129108 278798 129136 279783
rect 129096 278792 129148 278798
rect 129096 278734 129148 278740
rect 129278 272096 129334 272105
rect 129278 272031 129334 272040
rect 129186 249248 129242 249257
rect 129186 249183 129242 249192
rect 129004 237380 129056 237386
rect 129004 237322 129056 237328
rect 128358 234016 128414 234025
rect 128358 233951 128414 233960
rect 128372 233306 128400 233951
rect 128360 233300 128412 233306
rect 128360 233242 128412 233248
rect 129094 226400 129150 226409
rect 129094 226335 129150 226344
rect 128358 218784 128414 218793
rect 128358 218719 128414 218728
rect 128372 218074 128400 218719
rect 128360 218068 128412 218074
rect 128360 218010 128412 218016
rect 128360 211200 128412 211206
rect 128358 211168 128360 211177
rect 128412 211168 128414 211177
rect 128358 211103 128414 211112
rect 129002 203552 129058 203561
rect 129002 203487 129058 203496
rect 128634 195936 128690 195945
rect 128634 195871 128690 195880
rect 128648 194614 128676 195871
rect 128636 194608 128688 194614
rect 128636 194550 128688 194556
rect 126244 165572 126296 165578
rect 126244 165514 126296 165520
rect 19984 93832 20036 93838
rect 19984 93774 20036 93780
rect 15844 51060 15896 51066
rect 15844 51002 15896 51008
rect 11704 35896 11756 35902
rect 11704 35838 11756 35844
rect 129016 22098 129044 203487
rect 129108 64870 129136 226335
rect 129200 109002 129228 249183
rect 129292 151774 129320 272031
rect 129384 194546 129412 295015
rect 453302 288144 453358 288153
rect 453302 288079 453358 288088
rect 453026 281072 453082 281081
rect 453026 281007 453082 281016
rect 453040 280226 453068 281007
rect 453028 280220 453080 280226
rect 453028 280162 453080 280168
rect 452842 252512 452898 252521
rect 452842 252447 452898 252456
rect 452856 250510 452884 252447
rect 452844 250504 452896 250510
rect 452844 250446 452896 250452
rect 453118 231160 453174 231169
rect 453118 231095 453174 231104
rect 453132 230518 453160 231095
rect 453120 230512 453172 230518
rect 453120 230454 453172 230460
rect 453316 218006 453344 288079
rect 453408 229090 453436 295151
rect 453500 264926 453528 309431
rect 453592 276010 453620 316639
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 454684 302388 454736 302394
rect 454684 302330 454736 302336
rect 453580 276004 453632 276010
rect 453580 275946 453632 275952
rect 453670 273864 453726 273873
rect 453670 273799 453726 273808
rect 453578 266792 453634 266801
rect 453578 266727 453634 266736
rect 453488 264920 453540 264926
rect 453488 264862 453540 264868
rect 453486 245440 453542 245449
rect 453486 245375 453542 245384
rect 453396 229084 453448 229090
rect 453396 229026 453448 229032
rect 453394 224088 453450 224097
rect 453394 224023 453450 224032
rect 453304 218000 453356 218006
rect 453304 217942 453356 217948
rect 452934 217016 452990 217025
rect 452934 216951 452990 216960
rect 452948 216850 452976 216951
rect 452936 216844 452988 216850
rect 452936 216786 452988 216792
rect 453302 202736 453358 202745
rect 453302 202671 453358 202680
rect 129372 194540 129424 194546
rect 129372 194482 129424 194488
rect 135732 192222 136482 192250
rect 131132 192086 132434 192114
rect 132512 192086 133170 192114
rect 129280 151768 129332 151774
rect 129280 151710 129332 151716
rect 129188 108996 129240 109002
rect 129188 108938 129240 108944
rect 129096 64864 129148 64870
rect 129096 64806 129148 64812
rect 129004 22092 129056 22098
rect 129004 22034 129056 22040
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 127808 4140 127860 4146
rect 127808 4082 127860 4088
rect 126612 3732 126664 3738
rect 126612 3674 126664 3680
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 126624 480 126652 3674
rect 127820 480 127848 4082
rect 130200 4072 130252 4078
rect 130200 4014 130252 4020
rect 129004 4004 129056 4010
rect 129004 3946 129056 3952
rect 129016 480 129044 3946
rect 130212 480 130240 4014
rect 131132 3534 131160 192086
rect 131120 3528 131172 3534
rect 131120 3470 131172 3476
rect 132512 3466 132540 192086
rect 133880 181484 133932 181490
rect 133880 181426 133932 181432
rect 133892 4146 133920 181426
rect 133880 4140 133932 4146
rect 133880 4082 133932 4088
rect 133984 3738 134012 192100
rect 134536 192086 134826 192114
rect 135272 192086 135654 192114
rect 134536 181490 134564 192086
rect 134524 181484 134576 181490
rect 134524 181426 134576 181432
rect 135272 4010 135300 192086
rect 135732 189258 135760 192222
rect 135640 189230 135760 189258
rect 136652 192086 137310 192114
rect 135640 186266 135668 189230
rect 135548 186238 135668 186266
rect 135548 183569 135576 186238
rect 135350 183560 135406 183569
rect 135350 183495 135406 183504
rect 135534 183560 135590 183569
rect 135534 183495 135590 183504
rect 135364 173942 135392 183495
rect 135352 173936 135404 173942
rect 135352 173878 135404 173884
rect 135628 173936 135680 173942
rect 135628 173878 135680 173884
rect 135640 166954 135668 173878
rect 135548 166926 135668 166954
rect 135548 164218 135576 166926
rect 135352 164212 135404 164218
rect 135352 164154 135404 164160
rect 135536 164212 135588 164218
rect 135536 164154 135588 164160
rect 135364 154601 135392 164154
rect 135350 154592 135406 154601
rect 135350 154527 135406 154536
rect 135626 154592 135682 154601
rect 135626 154527 135682 154536
rect 135640 147642 135668 154527
rect 135548 147614 135668 147642
rect 135548 140026 135576 147614
rect 135364 139998 135576 140026
rect 135364 135289 135392 139998
rect 135350 135280 135406 135289
rect 135350 135215 135406 135224
rect 135626 135280 135682 135289
rect 135626 135215 135682 135224
rect 135640 128330 135668 135215
rect 135548 128302 135668 128330
rect 135548 120714 135576 128302
rect 135364 120686 135576 120714
rect 135364 115977 135392 120686
rect 135350 115968 135406 115977
rect 135350 115903 135406 115912
rect 135626 115968 135682 115977
rect 135626 115903 135682 115912
rect 135640 109018 135668 115903
rect 135548 108990 135668 109018
rect 135548 101402 135576 108990
rect 135364 101374 135576 101402
rect 135364 96665 135392 101374
rect 135350 96656 135406 96665
rect 135350 96591 135406 96600
rect 135626 96656 135682 96665
rect 135626 96591 135682 96600
rect 135640 89706 135668 96591
rect 135456 89678 135668 89706
rect 135456 86970 135484 89678
rect 135444 86964 135496 86970
rect 135444 86906 135496 86912
rect 135352 77308 135404 77314
rect 135352 77250 135404 77256
rect 135364 77178 135392 77250
rect 135352 77172 135404 77178
rect 135352 77114 135404 77120
rect 135444 70304 135496 70310
rect 135444 70246 135496 70252
rect 135456 60722 135484 70246
rect 135444 60716 135496 60722
rect 135444 60658 135496 60664
rect 135628 60716 135680 60722
rect 135628 60658 135680 60664
rect 135640 57934 135668 60658
rect 135628 57928 135680 57934
rect 135628 57870 135680 57876
rect 135536 48340 135588 48346
rect 135536 48282 135588 48288
rect 135548 41426 135576 48282
rect 135456 41410 135576 41426
rect 135444 41404 135576 41410
rect 135496 41398 135576 41404
rect 135628 41404 135680 41410
rect 135444 41346 135496 41352
rect 135628 41346 135680 41352
rect 135640 38622 135668 41346
rect 135628 38616 135680 38622
rect 135628 38558 135680 38564
rect 135536 29028 135588 29034
rect 135536 28970 135588 28976
rect 135548 22114 135576 28970
rect 135456 22098 135576 22114
rect 135444 22092 135576 22098
rect 135496 22086 135576 22092
rect 135628 22092 135680 22098
rect 135444 22034 135496 22040
rect 135628 22034 135680 22040
rect 135640 19310 135668 22034
rect 135628 19304 135680 19310
rect 135628 19246 135680 19252
rect 135628 12300 135680 12306
rect 135628 12242 135680 12248
rect 135640 4078 135668 12242
rect 135628 4072 135680 4078
rect 135628 4014 135680 4020
rect 135260 4004 135312 4010
rect 135260 3946 135312 3952
rect 133972 3732 134024 3738
rect 133972 3674 134024 3680
rect 132500 3460 132552 3466
rect 132500 3402 132552 3408
rect 134892 3460 134944 3466
rect 134892 3402 134944 3408
rect 133788 3324 133840 3330
rect 133788 3266 133840 3272
rect 132592 3188 132644 3194
rect 132592 3130 132644 3136
rect 131396 3120 131448 3126
rect 131396 3062 131448 3068
rect 131408 480 131436 3062
rect 132604 480 132632 3130
rect 133800 480 133828 3266
rect 134904 480 134932 3402
rect 136088 3256 136140 3262
rect 136088 3198 136140 3204
rect 136100 480 136128 3198
rect 136652 3126 136680 192086
rect 138020 185632 138072 185638
rect 138020 185574 138072 185580
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 136640 3120 136692 3126
rect 136640 3062 136692 3068
rect 137296 480 137324 3470
rect 138032 3330 138060 185574
rect 138020 3324 138072 3330
rect 138020 3266 138072 3272
rect 138124 3194 138152 192100
rect 138584 192086 138966 192114
rect 139504 192086 139794 192114
rect 140240 192086 140622 192114
rect 140792 192086 141450 192114
rect 142172 192086 142278 192114
rect 142448 192086 143106 192114
rect 143644 192086 143934 192114
rect 144472 192086 144762 192114
rect 144932 192086 145590 192114
rect 138584 185638 138612 192086
rect 138572 185632 138624 185638
rect 138572 185574 138624 185580
rect 139400 185632 139452 185638
rect 139400 185574 139452 185580
rect 138480 3936 138532 3942
rect 138480 3878 138532 3884
rect 138112 3188 138164 3194
rect 138112 3130 138164 3136
rect 138492 480 138520 3878
rect 139412 3262 139440 185574
rect 139504 3466 139532 192086
rect 140240 185638 140268 192086
rect 140228 185632 140280 185638
rect 140228 185574 140280 185580
rect 139676 4072 139728 4078
rect 139676 4014 139728 4020
rect 139492 3460 139544 3466
rect 139492 3402 139544 3408
rect 139400 3256 139452 3262
rect 139400 3198 139452 3204
rect 139688 480 139716 4014
rect 140792 3534 140820 192086
rect 142068 4140 142120 4146
rect 142068 4082 142120 4088
rect 140872 4004 140924 4010
rect 140872 3946 140924 3952
rect 140780 3528 140832 3534
rect 140780 3470 140832 3476
rect 140884 480 140912 3946
rect 142080 480 142108 4082
rect 142172 3942 142200 192086
rect 142448 4078 142476 192086
rect 143540 185632 143592 185638
rect 143540 185574 143592 185580
rect 143552 4146 143580 185574
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 142436 4072 142488 4078
rect 142436 4014 142488 4020
rect 143644 4010 143672 192086
rect 144472 185638 144500 192086
rect 144460 185632 144512 185638
rect 144460 185574 144512 185580
rect 143632 4004 143684 4010
rect 143632 3946 143684 3952
rect 142160 3936 142212 3942
rect 142160 3878 142212 3884
rect 144460 3460 144512 3466
rect 144460 3402 144512 3408
rect 143264 2916 143316 2922
rect 143264 2858 143316 2864
rect 143276 480 143304 2858
rect 144472 480 144500 3402
rect 144932 2922 144960 192086
rect 146300 185632 146352 185638
rect 146300 185574 146352 185580
rect 146312 3534 146340 185574
rect 145656 3528 145708 3534
rect 145656 3470 145708 3476
rect 146300 3528 146352 3534
rect 146300 3470 146352 3476
rect 144920 2916 144972 2922
rect 144920 2858 144972 2864
rect 145668 480 145696 3470
rect 146404 3466 146432 192100
rect 146864 192086 147246 192114
rect 147784 192086 148074 192114
rect 148520 192086 148902 192114
rect 149072 192086 149730 192114
rect 150452 192086 150558 192114
rect 150636 192086 151386 192114
rect 151832 192086 152214 192114
rect 153042 192086 153148 192114
rect 153870 192086 154528 192114
rect 146864 185638 146892 192086
rect 146852 185632 146904 185638
rect 146852 185574 146904 185580
rect 147680 185632 147732 185638
rect 147680 185574 147732 185580
rect 146852 3596 146904 3602
rect 146852 3538 146904 3544
rect 146392 3460 146444 3466
rect 146392 3402 146444 3408
rect 146864 480 146892 3538
rect 147692 3482 147720 185574
rect 147784 3602 147812 192086
rect 148520 185638 148548 192086
rect 148508 185632 148560 185638
rect 148508 185574 148560 185580
rect 147772 3596 147824 3602
rect 147772 3538 147824 3544
rect 147692 3454 148088 3482
rect 148060 480 148088 3454
rect 149072 3346 149100 192086
rect 149072 3318 149284 3346
rect 149256 480 149284 3318
rect 150452 480 150480 192086
rect 150636 3534 150664 192086
rect 151832 3534 151860 192086
rect 153120 3534 153148 192086
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151544 3528 151596 3534
rect 151544 3470 151596 3476
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 152740 3528 152792 3534
rect 152740 3470 152792 3476
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 153936 3528 153988 3534
rect 153936 3470 153988 3476
rect 151556 480 151584 3470
rect 152752 480 152780 3470
rect 153948 480 153976 3470
rect 154500 3466 154528 192086
rect 154684 190126 154712 192100
rect 155434 192086 155908 192114
rect 154672 190120 154724 190126
rect 154672 190062 154724 190068
rect 155776 190120 155828 190126
rect 155776 190062 155828 190068
rect 155788 3534 155816 190062
rect 155776 3528 155828 3534
rect 155776 3470 155828 3476
rect 154488 3460 154540 3466
rect 154488 3402 154540 3408
rect 155132 3460 155184 3466
rect 155132 3402 155184 3408
rect 155144 480 155172 3402
rect 155880 3330 155908 192086
rect 156248 189378 156276 192100
rect 157090 192086 157196 192114
rect 156236 189372 156288 189378
rect 156236 189314 156288 189320
rect 156328 3528 156380 3534
rect 156328 3470 156380 3476
rect 155868 3324 155920 3330
rect 155868 3266 155920 3272
rect 156340 480 156368 3470
rect 157168 3058 157196 192086
rect 157248 189372 157300 189378
rect 157248 189314 157300 189320
rect 157260 3534 157288 189314
rect 157904 189106 157932 192100
rect 158732 189854 158760 192100
rect 159574 192086 160048 192114
rect 158720 189848 158772 189854
rect 158720 189790 158772 189796
rect 159916 189848 159968 189854
rect 159916 189790 159968 189796
rect 157892 189100 157944 189106
rect 157892 189042 157944 189048
rect 158628 189100 158680 189106
rect 158628 189042 158680 189048
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 158640 3466 158668 189042
rect 159928 4078 159956 189790
rect 160020 4146 160048 192086
rect 160388 189174 160416 192100
rect 161230 192086 161336 192114
rect 162058 192086 162808 192114
rect 160376 189168 160428 189174
rect 160376 189110 160428 189116
rect 160008 4140 160060 4146
rect 160008 4082 160060 4088
rect 159916 4072 159968 4078
rect 159916 4014 159968 4020
rect 158720 3528 158772 3534
rect 158720 3470 158772 3476
rect 158628 3460 158680 3466
rect 158628 3402 158680 3408
rect 157524 3324 157576 3330
rect 157524 3266 157576 3272
rect 157156 3052 157208 3058
rect 157156 2994 157208 3000
rect 157536 480 157564 3266
rect 158732 480 158760 3470
rect 161308 3466 161336 192086
rect 161388 189168 161440 189174
rect 161388 189110 161440 189116
rect 161400 3602 161428 189110
rect 162308 4072 162360 4078
rect 162308 4014 162360 4020
rect 161388 3596 161440 3602
rect 161388 3538 161440 3544
rect 161112 3460 161164 3466
rect 161112 3402 161164 3408
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 159916 3052 159968 3058
rect 159916 2994 159968 3000
rect 159928 480 159956 2994
rect 161124 480 161152 3402
rect 162320 480 162348 4014
rect 162780 3330 162808 192086
rect 162872 189106 162900 192100
rect 163714 192086 164096 192114
rect 162860 189100 162912 189106
rect 162860 189042 162912 189048
rect 163504 4140 163556 4146
rect 163504 4082 163556 4088
rect 162768 3324 162820 3330
rect 162768 3266 162820 3272
rect 163516 480 163544 4082
rect 164068 3398 164096 192086
rect 164528 189378 164556 192100
rect 165370 192086 165476 192114
rect 164516 189372 164568 189378
rect 164516 189314 164568 189320
rect 164148 189100 164200 189106
rect 164148 189042 164200 189048
rect 164056 3392 164108 3398
rect 164056 3334 164108 3340
rect 164160 3262 164188 189042
rect 164700 3596 164752 3602
rect 164700 3538 164752 3544
rect 164148 3256 164200 3262
rect 164148 3198 164200 3204
rect 164712 480 164740 3538
rect 165448 2922 165476 192086
rect 165528 189372 165580 189378
rect 165528 189314 165580 189320
rect 165540 3534 165568 189314
rect 166184 189106 166212 192100
rect 167012 189106 167040 192100
rect 167854 192086 168328 192114
rect 166172 189100 166224 189106
rect 166172 189042 166224 189048
rect 166908 189100 166960 189106
rect 166908 189042 166960 189048
rect 167000 189100 167052 189106
rect 167000 189042 167052 189048
rect 168196 189100 168248 189106
rect 168196 189042 168248 189048
rect 166920 4146 166948 189042
rect 166908 4140 166960 4146
rect 166908 4082 166960 4088
rect 168208 3874 168236 189042
rect 168196 3868 168248 3874
rect 168196 3810 168248 3816
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 168300 3466 168328 192086
rect 168668 190330 168696 192100
rect 169510 192086 169708 192114
rect 170338 192086 171088 192114
rect 168656 190324 168708 190330
rect 168656 190266 168708 190272
rect 169576 190324 169628 190330
rect 169576 190266 169628 190272
rect 169588 3942 169616 190266
rect 169576 3936 169628 3942
rect 169576 3878 169628 3884
rect 169680 3806 169708 192086
rect 169668 3800 169720 3806
rect 169668 3742 169720 3748
rect 171060 3534 171088 192086
rect 171152 189106 171180 192100
rect 171994 192086 172468 192114
rect 171140 189100 171192 189106
rect 171140 189042 171192 189048
rect 172336 189100 172388 189106
rect 172336 189042 172388 189048
rect 170588 3528 170640 3534
rect 170588 3470 170640 3476
rect 171048 3528 171100 3534
rect 171048 3470 171100 3476
rect 165896 3460 165948 3466
rect 165896 3402 165948 3408
rect 168288 3460 168340 3466
rect 168288 3402 168340 3408
rect 165436 2916 165488 2922
rect 165436 2858 165488 2864
rect 165908 480 165936 3402
rect 169392 3392 169444 3398
rect 169392 3334 169444 3340
rect 167092 3324 167144 3330
rect 167092 3266 167144 3272
rect 167104 480 167132 3266
rect 168196 3256 168248 3262
rect 168196 3198 168248 3204
rect 168208 480 168236 3198
rect 169404 480 169432 3334
rect 170600 480 170628 3470
rect 172348 3330 172376 189042
rect 172440 3670 172468 192086
rect 172808 189378 172836 192100
rect 173650 192086 173756 192114
rect 172796 189372 172848 189378
rect 172796 189314 172848 189320
rect 173728 4826 173756 192086
rect 173808 189372 173860 189378
rect 173808 189314 173860 189320
rect 173716 4820 173768 4826
rect 173716 4762 173768 4768
rect 172980 4140 173032 4146
rect 172980 4082 173032 4088
rect 172428 3664 172480 3670
rect 172428 3606 172480 3612
rect 172336 3324 172388 3330
rect 172336 3266 172388 3272
rect 171784 2916 171836 2922
rect 171784 2858 171836 2864
rect 171796 480 171824 2858
rect 172992 480 173020 4082
rect 173820 3602 173848 189314
rect 174464 189106 174492 192100
rect 175292 189446 175320 192100
rect 176120 189854 176148 192100
rect 176108 189848 176160 189854
rect 176108 189790 176160 189796
rect 175280 189440 175332 189446
rect 175280 189382 175332 189388
rect 176568 189440 176620 189446
rect 176568 189382 176620 189388
rect 174452 189100 174504 189106
rect 174452 189042 174504 189048
rect 175188 189100 175240 189106
rect 175188 189042 175240 189048
rect 175200 4010 175228 189042
rect 176580 4078 176608 189382
rect 176948 189106 176976 192100
rect 177790 192086 177988 192114
rect 176936 189100 176988 189106
rect 176936 189042 176988 189048
rect 177856 189100 177908 189106
rect 177856 189042 177908 189048
rect 176568 4072 176620 4078
rect 176568 4014 176620 4020
rect 175188 4004 175240 4010
rect 175188 3946 175240 3952
rect 177868 3942 177896 189042
rect 176568 3936 176620 3942
rect 176568 3878 176620 3884
rect 177856 3936 177908 3942
rect 177856 3878 177908 3884
rect 174176 3868 174228 3874
rect 174176 3810 174228 3816
rect 173808 3596 173860 3602
rect 173808 3538 173860 3544
rect 174188 480 174216 3810
rect 175372 3460 175424 3466
rect 175372 3402 175424 3408
rect 175384 480 175412 3402
rect 176580 480 176608 3878
rect 177764 3800 177816 3806
rect 177764 3742 177816 3748
rect 177776 480 177804 3742
rect 177960 3466 177988 192086
rect 178512 189106 178540 192100
rect 178500 189100 178552 189106
rect 178500 189042 178552 189048
rect 179236 189100 179288 189106
rect 179236 189042 179288 189048
rect 179248 6186 179276 189042
rect 179236 6180 179288 6186
rect 179236 6122 179288 6128
rect 179340 3534 179368 192100
rect 180182 192086 180748 192114
rect 180720 3738 180748 192086
rect 180996 189786 181024 192100
rect 181838 192086 182128 192114
rect 180984 189780 181036 189786
rect 180984 189722 181036 189728
rect 182100 3874 182128 192086
rect 182652 189446 182680 192100
rect 183388 192086 183494 192114
rect 184322 192086 184888 192114
rect 182640 189440 182692 189446
rect 182640 189382 182692 189388
rect 183388 7614 183416 192086
rect 184204 189848 184256 189854
rect 184204 189790 184256 189796
rect 183468 189440 183520 189446
rect 183468 189382 183520 189388
rect 183376 7608 183428 7614
rect 183376 7550 183428 7556
rect 182088 3868 182140 3874
rect 182088 3810 182140 3816
rect 183480 3806 183508 189382
rect 183744 4820 183796 4826
rect 183744 4762 183796 4768
rect 183468 3800 183520 3806
rect 183468 3742 183520 3748
rect 180708 3732 180760 3738
rect 180708 3674 180760 3680
rect 181352 3664 181404 3670
rect 181352 3606 181404 3612
rect 178960 3528 179012 3534
rect 178960 3470 179012 3476
rect 179328 3528 179380 3534
rect 179328 3470 179380 3476
rect 177948 3460 178000 3466
rect 177948 3402 178000 3408
rect 178972 480 179000 3470
rect 180156 3324 180208 3330
rect 180156 3266 180208 3272
rect 180168 480 180196 3266
rect 181364 480 181392 3606
rect 182548 3596 182600 3602
rect 182548 3538 182600 3544
rect 182560 480 182588 3538
rect 183756 480 183784 4762
rect 184216 4214 184244 189790
rect 184860 11762 184888 192086
rect 185136 189310 185164 192100
rect 185978 192086 186176 192114
rect 185124 189304 185176 189310
rect 185124 189246 185176 189252
rect 184848 11756 184900 11762
rect 184848 11698 184900 11704
rect 186148 9042 186176 192086
rect 186228 189304 186280 189310
rect 186228 189246 186280 189252
rect 186136 9036 186188 9042
rect 186136 8978 186188 8984
rect 184204 4208 184256 4214
rect 184204 4150 184256 4156
rect 186044 4072 186096 4078
rect 186044 4014 186096 4020
rect 184848 4004 184900 4010
rect 184848 3946 184900 3952
rect 184860 480 184888 3946
rect 186056 480 186084 4014
rect 186240 3670 186268 189246
rect 186792 189106 186820 192100
rect 186780 189100 186832 189106
rect 186780 189042 186832 189048
rect 187516 189100 187568 189106
rect 187516 189042 187568 189048
rect 187528 13122 187556 189042
rect 187516 13116 187568 13122
rect 187516 13058 187568 13064
rect 187240 4208 187292 4214
rect 187240 4150 187292 4156
rect 186228 3664 186280 3670
rect 186228 3606 186280 3612
rect 187252 480 187280 4150
rect 187620 3602 187648 192100
rect 188462 192086 189028 192114
rect 189000 10334 189028 192086
rect 189276 189106 189304 192100
rect 190118 192086 190408 192114
rect 189264 189100 189316 189106
rect 189264 189042 189316 189048
rect 190276 189100 190328 189106
rect 190276 189042 190328 189048
rect 190288 14482 190316 189042
rect 190276 14476 190328 14482
rect 190276 14418 190328 14424
rect 188988 10328 189040 10334
rect 188988 10270 189040 10276
rect 188436 3936 188488 3942
rect 188436 3878 188488 3884
rect 187608 3596 187660 3602
rect 187608 3538 187660 3544
rect 188448 480 188476 3878
rect 190380 3466 190408 192086
rect 190932 189106 190960 192100
rect 191668 192086 191774 192114
rect 192602 192086 193168 192114
rect 190920 189100 190972 189106
rect 190920 189042 190972 189048
rect 191668 15910 191696 192086
rect 192484 189780 192536 189786
rect 192484 189722 192536 189728
rect 191748 189100 191800 189106
rect 191748 189042 191800 189048
rect 191656 15904 191708 15910
rect 191656 15846 191708 15852
rect 191760 6186 191788 189042
rect 190828 6180 190880 6186
rect 190828 6122 190880 6128
rect 191748 6180 191800 6186
rect 191748 6122 191800 6128
rect 189632 3460 189684 3466
rect 189632 3402 189684 3408
rect 190368 3460 190420 3466
rect 190368 3402 190420 3408
rect 189644 480 189672 3402
rect 190840 480 190868 6122
rect 192496 4214 192524 189722
rect 192484 4208 192536 4214
rect 192484 4150 192536 4156
rect 193140 3534 193168 192086
rect 193416 189310 193444 192100
rect 194258 192086 194456 192114
rect 193404 189304 193456 189310
rect 193404 189246 193456 189252
rect 194428 17338 194456 192086
rect 194508 189304 194560 189310
rect 194508 189246 194560 189252
rect 194416 17332 194468 17338
rect 194416 17274 194468 17280
rect 194520 4826 194548 189246
rect 195072 189106 195100 192100
rect 195900 189786 195928 192100
rect 196742 192086 197308 192114
rect 195888 189780 195940 189786
rect 195888 189722 195940 189728
rect 195060 189100 195112 189106
rect 195060 189042 195112 189048
rect 195888 189100 195940 189106
rect 195888 189042 195940 189048
rect 194508 4820 194560 4826
rect 194508 4762 194560 4768
rect 194416 4208 194468 4214
rect 194416 4150 194468 4156
rect 193220 3732 193272 3738
rect 193220 3674 193272 3680
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 192036 480 192064 3470
rect 193232 480 193260 3674
rect 194428 480 194456 4150
rect 195900 3942 195928 189042
rect 197280 18698 197308 192086
rect 197556 189378 197584 192100
rect 198398 192086 198596 192114
rect 197544 189372 197596 189378
rect 197544 189314 197596 189320
rect 197268 18692 197320 18698
rect 197268 18634 197320 18640
rect 198568 7614 198596 192086
rect 198648 189372 198700 189378
rect 198648 189314 198700 189320
rect 198004 7608 198056 7614
rect 198004 7550 198056 7556
rect 198556 7608 198608 7614
rect 198556 7550 198608 7556
rect 195888 3936 195940 3942
rect 195888 3878 195940 3884
rect 195612 3868 195664 3874
rect 195612 3810 195664 3816
rect 195624 480 195652 3810
rect 196808 3800 196860 3806
rect 196808 3742 196860 3748
rect 196820 480 196848 3742
rect 198016 480 198044 7550
rect 198660 3874 198688 189314
rect 199212 189106 199240 192100
rect 199200 189100 199252 189106
rect 199200 189042 199252 189048
rect 198740 11756 198792 11762
rect 198740 11698 198792 11704
rect 198648 3868 198700 3874
rect 198648 3810 198700 3816
rect 198752 3346 198780 11698
rect 200040 3806 200068 192100
rect 200790 192086 201448 192114
rect 200764 189100 200816 189106
rect 200764 189042 200816 189048
rect 200776 20058 200804 189042
rect 200764 20052 200816 20058
rect 200764 19994 200816 20000
rect 201420 8974 201448 192086
rect 201604 190194 201632 192100
rect 202446 192086 202828 192114
rect 201592 190188 201644 190194
rect 201592 190130 201644 190136
rect 202696 190188 202748 190194
rect 202696 190130 202748 190136
rect 202708 21486 202736 190130
rect 202696 21480 202748 21486
rect 202696 21422 202748 21428
rect 201500 13116 201552 13122
rect 201500 13058 201552 13064
rect 201408 8968 201460 8974
rect 201408 8910 201460 8916
rect 200028 3800 200080 3806
rect 200028 3742 200080 3748
rect 200396 3664 200448 3670
rect 200396 3606 200448 3612
rect 198752 3318 199240 3346
rect 199212 480 199240 3318
rect 200408 480 200436 3606
rect 201512 3602 201540 13058
rect 201592 9036 201644 9042
rect 201592 8978 201644 8984
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 201604 3482 201632 8978
rect 202800 3738 202828 192086
rect 203260 189446 203288 192100
rect 203248 189440 203300 189446
rect 203248 189382 203300 189388
rect 204088 22778 204116 192100
rect 204930 192086 205588 192114
rect 204168 189440 204220 189446
rect 204168 189382 204220 189388
rect 204076 22772 204128 22778
rect 204076 22714 204128 22720
rect 204180 11762 204208 189382
rect 204168 11756 204220 11762
rect 204168 11698 204220 11704
rect 204260 10328 204312 10334
rect 204260 10270 204312 10276
rect 202788 3732 202840 3738
rect 202788 3674 202840 3680
rect 203892 3664 203944 3670
rect 203892 3606 203944 3612
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202708 480 202736 3538
rect 203904 480 203932 3606
rect 204272 3346 204300 10270
rect 205560 4010 205588 192086
rect 205744 189310 205772 192100
rect 206586 192086 206876 192114
rect 205732 189304 205784 189310
rect 205732 189246 205784 189252
rect 206848 24138 206876 192086
rect 206928 189304 206980 189310
rect 206928 189246 206980 189252
rect 206836 24132 206888 24138
rect 206836 24074 206888 24080
rect 205640 14476 205692 14482
rect 205640 14418 205692 14424
rect 205548 4004 205600 4010
rect 205548 3946 205600 3952
rect 205652 3346 205680 14418
rect 206940 10334 206968 189246
rect 207400 189106 207428 192100
rect 207388 189100 207440 189106
rect 207388 189042 207440 189048
rect 208228 13190 208256 192100
rect 209070 192086 209728 192114
rect 208308 189100 208360 189106
rect 208308 189042 208360 189048
rect 208216 13184 208268 13190
rect 208216 13126 208268 13132
rect 206928 10328 206980 10334
rect 206928 10270 206980 10276
rect 208320 3738 208348 189042
rect 209700 17270 209728 192086
rect 209884 189310 209912 192100
rect 210726 192086 211016 192114
rect 209872 189304 209924 189310
rect 209872 189246 209924 189252
rect 209688 17264 209740 17270
rect 209688 17206 209740 17212
rect 209872 15904 209924 15910
rect 209872 15846 209924 15852
rect 208676 6180 208728 6186
rect 208676 6122 208728 6128
rect 208308 3732 208360 3738
rect 208308 3674 208360 3680
rect 207480 3460 207532 3466
rect 207480 3402 207532 3408
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3402
rect 208688 480 208716 6122
rect 209884 480 209912 15846
rect 210988 6186 211016 192086
rect 211068 189304 211120 189310
rect 211068 189246 211120 189252
rect 210976 6180 211028 6186
rect 210976 6122 211028 6128
rect 211080 5250 211108 189246
rect 211540 189106 211568 192100
rect 212382 192086 212488 192114
rect 213210 192086 213592 192114
rect 211528 189100 211580 189106
rect 211528 189042 211580 189048
rect 212356 189100 212408 189106
rect 212356 189042 212408 189048
rect 212368 25634 212396 189042
rect 212356 25628 212408 25634
rect 212356 25570 212408 25576
rect 210988 5222 211108 5250
rect 210988 3466 211016 5222
rect 212264 4820 212316 4826
rect 212264 4762 212316 4768
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 210976 3460 211028 3466
rect 210976 3402 211028 3408
rect 211080 480 211108 3470
rect 212276 480 212304 4762
rect 212460 3466 212488 192086
rect 213184 189780 213236 189786
rect 213184 189722 213236 189728
rect 212540 17332 212592 17338
rect 212540 17274 212592 17280
rect 212448 3460 212500 3466
rect 212448 3402 212500 3408
rect 212552 3346 212580 17274
rect 213196 4214 213224 189722
rect 213564 189174 213592 192086
rect 214024 189378 214052 192100
rect 214866 192086 215156 192114
rect 214012 189372 214064 189378
rect 214012 189314 214064 189320
rect 213552 189168 213604 189174
rect 213552 189110 213604 189116
rect 215128 35222 215156 192086
rect 215208 189372 215260 189378
rect 215208 189314 215260 189320
rect 215116 35216 215168 35222
rect 215116 35158 215168 35164
rect 215220 18630 215248 189314
rect 215680 189106 215708 192100
rect 215668 189100 215720 189106
rect 215668 189042 215720 189048
rect 216508 26926 216536 192100
rect 217350 192086 218008 192114
rect 216588 189100 216640 189106
rect 216588 189042 216640 189048
rect 216496 26920 216548 26926
rect 216496 26862 216548 26868
rect 215208 18624 215260 18630
rect 215208 18566 215260 18572
rect 216600 14482 216628 189042
rect 217980 36582 218008 192086
rect 218164 189106 218192 192100
rect 219006 192086 219296 192114
rect 218152 189100 218204 189106
rect 218152 189042 218204 189048
rect 217968 36576 218020 36582
rect 217968 36518 218020 36524
rect 219268 19990 219296 192086
rect 219820 190262 219848 192100
rect 220662 192086 220768 192114
rect 219808 190256 219860 190262
rect 219808 190198 219860 190204
rect 220636 190256 220688 190262
rect 220636 190198 220688 190204
rect 219348 189100 219400 189106
rect 219348 189042 219400 189048
rect 219256 19984 219308 19990
rect 219256 19926 219308 19932
rect 216680 18692 216732 18698
rect 216680 18634 216732 18640
rect 216588 14476 216640 14482
rect 216588 14418 216640 14424
rect 213184 4208 213236 4214
rect 213184 4150 213236 4156
rect 215852 4208 215904 4214
rect 215852 4150 215904 4156
rect 214656 3936 214708 3942
rect 214656 3878 214708 3884
rect 212552 3318 213500 3346
rect 213472 480 213500 3318
rect 214668 480 214696 3878
rect 215864 480 215892 4150
rect 216692 3346 216720 18634
rect 219360 7614 219388 189042
rect 220648 37942 220676 190198
rect 220636 37936 220688 37942
rect 220636 37878 220688 37884
rect 219440 20052 219492 20058
rect 219440 19994 219492 20000
rect 219348 7608 219400 7614
rect 219348 7550 219400 7556
rect 219348 7404 219400 7410
rect 219348 7346 219400 7352
rect 218152 3868 218204 3874
rect 218152 3810 218204 3816
rect 216692 3318 217088 3346
rect 217060 480 217088 3318
rect 218164 480 218192 3810
rect 219360 480 219388 7346
rect 219452 3482 219480 19994
rect 220740 15910 220768 192086
rect 221280 189168 221332 189174
rect 221280 189110 221332 189116
rect 221292 188986 221320 189110
rect 221476 189106 221504 192100
rect 222304 189514 222332 192100
rect 223132 189786 223160 192100
rect 223120 189780 223172 189786
rect 223120 189722 223172 189728
rect 222292 189508 222344 189514
rect 222292 189450 222344 189456
rect 223488 189508 223540 189514
rect 223488 189450 223540 189456
rect 221464 189100 221516 189106
rect 221464 189042 221516 189048
rect 222844 189100 222896 189106
rect 222844 189042 222896 189048
rect 221292 188958 221504 188986
rect 220728 15904 220780 15910
rect 220728 15846 220780 15852
rect 221476 4826 221504 188958
rect 222856 21418 222884 189042
rect 223500 39370 223528 189450
rect 223868 189310 223896 192100
rect 224710 192086 224816 192114
rect 225538 192086 226288 192114
rect 223856 189304 223908 189310
rect 223856 189246 223908 189252
rect 224788 40730 224816 192086
rect 224868 189304 224920 189310
rect 224868 189246 224920 189252
rect 224776 40724 224828 40730
rect 224776 40666 224828 40672
rect 223488 39364 223540 39370
rect 223488 39306 223540 39312
rect 224880 28286 224908 189246
rect 224868 28280 224920 28286
rect 224868 28222 224920 28228
rect 223580 21480 223632 21486
rect 223580 21422 223632 21428
rect 222844 21412 222896 21418
rect 222844 21354 222896 21360
rect 222936 8968 222988 8974
rect 222936 8910 222988 8916
rect 221464 4820 221516 4826
rect 221464 4762 221516 4768
rect 219452 3454 220584 3482
rect 220556 480 220584 3454
rect 221740 3120 221792 3126
rect 221740 3062 221792 3068
rect 221752 480 221780 3062
rect 222948 480 222976 8910
rect 223592 3482 223620 21422
rect 226260 8974 226288 192086
rect 226352 189106 226380 192100
rect 227194 192086 227576 192114
rect 226340 189100 226392 189106
rect 226340 189042 226392 189048
rect 227548 42090 227576 192086
rect 228008 189106 228036 192100
rect 228850 192086 228956 192114
rect 227628 189100 227680 189106
rect 227628 189042 227680 189048
rect 227996 189100 228048 189106
rect 227996 189042 228048 189048
rect 227536 42084 227588 42090
rect 227536 42026 227588 42032
rect 227640 29714 227668 189042
rect 227628 29708 227680 29714
rect 227628 29650 227680 29656
rect 228928 22778 228956 192086
rect 229664 189718 229692 192100
rect 229652 189712 229704 189718
rect 229652 189654 229704 189660
rect 230388 189712 230440 189718
rect 230388 189654 230440 189660
rect 229008 189100 229060 189106
rect 229008 189042 229060 189048
rect 227812 22772 227864 22778
rect 227812 22714 227864 22720
rect 228916 22772 228968 22778
rect 228916 22714 228968 22720
rect 226340 11756 226392 11762
rect 226340 11698 226392 11704
rect 226248 8968 226300 8974
rect 226248 8910 226300 8916
rect 225328 3664 225380 3670
rect 225328 3606 225380 3612
rect 223592 3454 224172 3482
rect 224144 480 224172 3454
rect 225340 480 225368 3606
rect 226352 3482 226380 11698
rect 226352 3454 226564 3482
rect 226536 480 226564 3454
rect 227824 1442 227852 22714
rect 229020 11762 229048 189042
rect 230400 43450 230428 189654
rect 230492 189310 230520 192100
rect 231334 192086 231716 192114
rect 230480 189304 230532 189310
rect 230480 189246 230532 189252
rect 230388 43444 230440 43450
rect 230388 43386 230440 43392
rect 231688 24138 231716 192086
rect 231768 189304 231820 189310
rect 231768 189246 231820 189252
rect 230480 24132 230532 24138
rect 230480 24074 230532 24080
rect 231676 24132 231728 24138
rect 231676 24074 231728 24080
rect 229008 11756 229060 11762
rect 229008 11698 229060 11704
rect 229100 10328 229152 10334
rect 229100 10270 229152 10276
rect 228916 3732 228968 3738
rect 228916 3674 228968 3680
rect 227732 1414 227852 1442
rect 227732 480 227760 1414
rect 228928 480 228956 3674
rect 229112 3482 229140 10270
rect 230492 3482 230520 24074
rect 231780 10334 231808 189246
rect 232148 189106 232176 192100
rect 232990 192086 233188 192114
rect 233818 192086 234568 192114
rect 232136 189100 232188 189106
rect 232136 189042 232188 189048
rect 233056 189100 233108 189106
rect 233056 189042 233108 189048
rect 233068 49026 233096 189042
rect 233056 49020 233108 49026
rect 233056 48962 233108 48968
rect 233160 13122 233188 192086
rect 234540 25566 234568 192086
rect 234632 189582 234660 192100
rect 234620 189576 234672 189582
rect 234620 189518 234672 189524
rect 235460 188358 235488 192100
rect 235816 189576 235868 189582
rect 235816 189518 235868 189524
rect 235448 188352 235500 188358
rect 235448 188294 235500 188300
rect 235828 44878 235856 189518
rect 236288 189378 236316 192100
rect 237130 192086 237236 192114
rect 236276 189372 236328 189378
rect 236276 189314 236328 189320
rect 237208 47598 237236 192086
rect 237944 189990 237972 192100
rect 237932 189984 237984 189990
rect 237932 189926 237984 189932
rect 238668 189984 238720 189990
rect 238668 189926 238720 189932
rect 237288 189372 237340 189378
rect 237288 189314 237340 189320
rect 237196 47592 237248 47598
rect 237196 47534 237248 47540
rect 235816 44872 235868 44878
rect 235816 44814 235868 44820
rect 237300 31142 237328 189314
rect 237288 31136 237340 31142
rect 237288 31078 237340 31084
rect 237380 25628 237432 25634
rect 237380 25570 237432 25576
rect 234528 25560 234580 25566
rect 234528 25502 234580 25508
rect 234620 17264 234672 17270
rect 234620 17206 234672 17212
rect 233240 13184 233292 13190
rect 233240 13126 233292 13132
rect 233148 13116 233200 13122
rect 233148 13058 233200 13064
rect 231768 10328 231820 10334
rect 231768 10270 231820 10276
rect 232504 3596 232556 3602
rect 232504 3538 232556 3544
rect 229112 3454 230152 3482
rect 230492 3454 231348 3482
rect 230124 480 230152 3454
rect 231320 480 231348 3454
rect 232516 480 232544 3538
rect 233252 3482 233280 13126
rect 234632 3482 234660 17206
rect 237196 6180 237248 6186
rect 237196 6122 237248 6128
rect 236000 3528 236052 3534
rect 233252 3454 233740 3482
rect 234632 3454 234844 3482
rect 236000 3470 236052 3476
rect 233712 480 233740 3454
rect 234816 480 234844 3454
rect 236012 480 236040 3470
rect 237208 480 237236 6122
rect 237392 3482 237420 25570
rect 238680 6186 238708 189926
rect 238772 189310 238800 192100
rect 239614 192086 239996 192114
rect 238760 189304 238812 189310
rect 238760 189246 238812 189252
rect 239968 50386 239996 192086
rect 240428 189854 240456 192100
rect 241270 192086 241468 192114
rect 242098 192086 242848 192114
rect 240416 189848 240468 189854
rect 240416 189790 240468 189796
rect 240048 189304 240100 189310
rect 240048 189246 240100 189252
rect 239956 50380 240008 50386
rect 239956 50322 240008 50328
rect 240060 32502 240088 189246
rect 241440 33794 241468 192086
rect 242164 189780 242216 189786
rect 242164 189722 242216 189728
rect 241428 33788 241480 33794
rect 241428 33730 241480 33736
rect 240048 32496 240100 32502
rect 240048 32438 240100 32444
rect 241520 18624 241572 18630
rect 241520 18566 241572 18572
rect 238668 6180 238720 6186
rect 238668 6122 238720 6128
rect 240784 4820 240836 4826
rect 240784 4762 240836 4768
rect 237392 3454 238432 3482
rect 238404 480 238432 3454
rect 239588 3460 239640 3466
rect 239588 3402 239640 3408
rect 239600 480 239628 3402
rect 240796 480 240824 4762
rect 241532 3482 241560 18566
rect 242176 4826 242204 189722
rect 242820 51746 242848 192086
rect 242912 189106 242940 192100
rect 243754 192086 244136 192114
rect 242900 189100 242952 189106
rect 242900 189042 242952 189048
rect 242808 51740 242860 51746
rect 242808 51682 242860 51688
rect 244108 46238 244136 192086
rect 244568 190126 244596 192100
rect 245410 192086 245608 192114
rect 244556 190120 244608 190126
rect 244556 190062 244608 190068
rect 245476 190120 245528 190126
rect 245476 190062 245528 190068
rect 244188 189100 244240 189106
rect 244188 189042 244240 189048
rect 244096 46232 244148 46238
rect 244096 46174 244148 46180
rect 242900 35216 242952 35222
rect 242900 35158 242952 35164
rect 242164 4820 242216 4826
rect 242164 4762 242216 4768
rect 242912 3482 242940 35158
rect 244200 17270 244228 189042
rect 245488 53106 245516 190062
rect 245476 53100 245528 53106
rect 245476 53042 245528 53048
rect 244280 26920 244332 26926
rect 244280 26862 244332 26868
rect 244188 17264 244240 17270
rect 244188 17206 244240 17212
rect 244292 3534 244320 26862
rect 245580 14482 245608 192086
rect 246132 189106 246160 192100
rect 246868 192086 246974 192114
rect 247802 192086 248368 192114
rect 246120 189100 246172 189106
rect 246120 189042 246172 189048
rect 246868 54534 246896 192086
rect 246948 189100 247000 189106
rect 246948 189042 247000 189048
rect 246856 54528 246908 54534
rect 246856 54470 246908 54476
rect 245660 36576 245712 36582
rect 245660 36518 245712 36524
rect 244372 14476 244424 14482
rect 244372 14418 244424 14424
rect 245568 14476 245620 14482
rect 245568 14418 245620 14424
rect 244280 3528 244332 3534
rect 241532 3454 242020 3482
rect 242912 3454 243216 3482
rect 244280 3470 244332 3476
rect 241992 480 242020 3454
rect 243188 480 243216 3454
rect 244384 480 244412 14418
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245672 3482 245700 36518
rect 246960 26926 246988 189042
rect 246948 26920 247000 26926
rect 246948 26862 247000 26868
rect 248340 7614 248368 192086
rect 248616 189310 248644 192100
rect 249458 192086 249656 192114
rect 248604 189304 248656 189310
rect 248604 189246 248656 189252
rect 249628 57254 249656 192086
rect 250272 189514 250300 192100
rect 251008 192086 251114 192114
rect 251942 192086 252508 192114
rect 250260 189508 250312 189514
rect 250260 189450 250312 189456
rect 249708 189304 249760 189310
rect 249708 189246 249760 189252
rect 249616 57248 249668 57254
rect 249616 57190 249668 57196
rect 249720 35222 249748 189246
rect 249800 37936 249852 37942
rect 249800 37878 249852 37884
rect 249708 35216 249760 35222
rect 249708 35158 249760 35164
rect 248420 19984 248472 19990
rect 248420 19926 248472 19932
rect 247960 7608 248012 7614
rect 247960 7550 248012 7556
rect 248328 7608 248380 7614
rect 248328 7550 248380 7556
rect 245580 480 245608 3470
rect 245672 3454 246804 3482
rect 246776 480 246804 3454
rect 247972 480 248000 7550
rect 248432 3482 248460 19926
rect 249812 3482 249840 37878
rect 251008 36650 251036 192086
rect 251088 189508 251140 189514
rect 251088 189450 251140 189456
rect 250996 36644 251048 36650
rect 250996 36586 251048 36592
rect 251100 18630 251128 189450
rect 252480 29646 252508 192086
rect 252756 186998 252784 192100
rect 253584 190126 253612 192100
rect 254426 192086 255176 192114
rect 253572 190120 253624 190126
rect 253572 190062 253624 190068
rect 252744 186992 252796 186998
rect 252744 186934 252796 186940
rect 255148 58682 255176 192086
rect 255136 58676 255188 58682
rect 255136 58618 255188 58624
rect 252560 39364 252612 39370
rect 252560 39306 252612 39312
rect 252468 29640 252520 29646
rect 252468 29582 252520 29588
rect 251088 18624 251140 18630
rect 251088 18566 251140 18572
rect 251180 15904 251232 15910
rect 251180 15846 251232 15852
rect 251192 3482 251220 15846
rect 252572 3534 252600 39306
rect 252652 21412 252704 21418
rect 252652 21354 252704 21360
rect 252560 3528 252612 3534
rect 248432 3454 249196 3482
rect 249812 3454 250392 3482
rect 251192 3454 251496 3482
rect 252560 3470 252612 3476
rect 249168 480 249196 3454
rect 250364 480 250392 3454
rect 251468 480 251496 3454
rect 252664 480 252692 21354
rect 255240 15978 255268 192100
rect 256082 192086 256648 192114
rect 255964 189848 256016 189854
rect 255964 189790 256016 189796
rect 255320 28280 255372 28286
rect 255320 28222 255372 28228
rect 255228 15972 255280 15978
rect 255228 15914 255280 15920
rect 255044 4820 255096 4826
rect 255044 4762 255096 4768
rect 253848 3528 253900 3534
rect 253848 3470 253900 3476
rect 253860 480 253888 3470
rect 255056 480 255084 4762
rect 255332 3618 255360 28222
rect 255976 4826 256004 189790
rect 256620 37942 256648 192086
rect 256896 189106 256924 192100
rect 257344 190120 257396 190126
rect 257344 190062 257396 190068
rect 256884 189100 256936 189106
rect 256884 189042 256936 189048
rect 256700 40724 256752 40730
rect 256700 40666 256752 40672
rect 256608 37936 256660 37942
rect 256608 37878 256660 37884
rect 255964 4820 256016 4826
rect 255964 4762 256016 4768
rect 255332 3590 256280 3618
rect 256252 480 256280 3590
rect 256712 3482 256740 40666
rect 257356 28286 257384 190062
rect 257724 189854 257752 192100
rect 257712 189848 257764 189854
rect 257712 189790 257764 189796
rect 258552 189106 258580 192100
rect 257988 189100 258040 189106
rect 257988 189042 258040 189048
rect 258540 189100 258592 189106
rect 258540 189042 258592 189048
rect 259276 189100 259328 189106
rect 259276 189042 259328 189048
rect 258000 60042 258028 189042
rect 259288 177342 259316 189042
rect 259276 177336 259328 177342
rect 259276 177278 259328 177284
rect 259380 62830 259408 192100
rect 260222 192086 260788 192114
rect 259368 62824 259420 62830
rect 259368 62766 259420 62772
rect 257988 60036 258040 60042
rect 257988 59978 258040 59984
rect 259460 29708 259512 29714
rect 259460 29650 259512 29656
rect 257344 28280 257396 28286
rect 257344 28222 257396 28228
rect 258632 8968 258684 8974
rect 258632 8910 258684 8916
rect 256712 3454 257476 3482
rect 257448 480 257476 3454
rect 258644 480 258672 8910
rect 259472 3482 259500 29650
rect 260760 8974 260788 192086
rect 261036 189378 261064 192100
rect 261878 192086 262076 192114
rect 261024 189372 261076 189378
rect 261024 189314 261076 189320
rect 262048 64190 262076 192086
rect 262128 189372 262180 189378
rect 262128 189314 262180 189320
rect 262036 64184 262088 64190
rect 262036 64126 262088 64132
rect 260840 42084 260892 42090
rect 260840 42026 260892 42032
rect 260748 8968 260800 8974
rect 260748 8910 260800 8916
rect 260852 3482 260880 42026
rect 262140 39370 262168 189314
rect 262692 189106 262720 192100
rect 263428 192086 263534 192114
rect 264362 192086 264928 192114
rect 262680 189100 262732 189106
rect 262680 189042 262732 189048
rect 263428 40730 263456 192086
rect 263508 189100 263560 189106
rect 263508 189042 263560 189048
rect 263416 40724 263468 40730
rect 263416 40666 263468 40672
rect 262128 39364 262180 39370
rect 262128 39306 262180 39312
rect 262220 22772 262272 22778
rect 262220 22714 262272 22720
rect 262232 3602 262260 22714
rect 263520 11762 263548 189042
rect 263600 43444 263652 43450
rect 263600 43386 263652 43392
rect 262312 11756 262364 11762
rect 262312 11698 262364 11704
rect 263508 11756 263560 11762
rect 263508 11698 263560 11704
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 262324 3482 262352 11698
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 259472 3454 259868 3482
rect 260852 3454 261064 3482
rect 259840 480 259868 3454
rect 261036 480 261064 3454
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3538
rect 263612 3482 263640 43386
rect 264900 32434 264928 192086
rect 265176 189310 265204 192100
rect 266018 192086 266216 192114
rect 265164 189304 265216 189310
rect 265164 189246 265216 189252
rect 266188 42158 266216 192086
rect 266268 189304 266320 189310
rect 266268 189246 266320 189252
rect 266176 42152 266228 42158
rect 266176 42094 266228 42100
rect 264888 32428 264940 32434
rect 264888 32370 264940 32376
rect 266280 19990 266308 189246
rect 266832 189106 266860 192100
rect 266820 189100 266872 189106
rect 266820 189042 266872 189048
rect 267556 189100 267608 189106
rect 267556 189042 267608 189048
rect 267568 65550 267596 189042
rect 267556 65544 267608 65550
rect 267556 65486 267608 65492
rect 266360 24132 266412 24138
rect 266360 24074 266412 24080
rect 266268 19984 266320 19990
rect 266268 19926 266320 19932
rect 264980 10328 265032 10334
rect 264980 10270 265032 10276
rect 264992 3482 265020 10270
rect 266372 3482 266400 24074
rect 267660 10334 267688 192100
rect 268502 192086 269068 192114
rect 267740 49020 267792 49026
rect 267740 48962 267792 48968
rect 267648 10328 267700 10334
rect 267648 10270 267700 10276
rect 263612 3454 264652 3482
rect 264992 3454 265848 3482
rect 266372 3454 267044 3482
rect 264624 480 264652 3454
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 267752 3346 267780 48962
rect 269040 31074 269068 192086
rect 269224 189990 269252 192100
rect 270066 192086 270448 192114
rect 269212 189984 269264 189990
rect 269212 189926 269264 189932
rect 270316 189984 270368 189990
rect 270316 189926 270368 189932
rect 270328 66910 270356 189926
rect 270316 66904 270368 66910
rect 270316 66846 270368 66852
rect 269028 31068 269080 31074
rect 269028 31010 269080 31016
rect 270420 13122 270448 192086
rect 270880 189990 270908 192100
rect 271722 192086 271828 192114
rect 272550 192086 273208 192114
rect 270868 189984 270920 189990
rect 270868 189926 270920 189932
rect 271800 68338 271828 192086
rect 271972 189984 272024 189990
rect 271972 189926 272024 189932
rect 271984 188358 272012 189926
rect 271880 188352 271932 188358
rect 271880 188294 271932 188300
rect 271972 188352 272024 188358
rect 271972 188294 272024 188300
rect 271788 68332 271840 68338
rect 271788 68274 271840 68280
rect 270500 44872 270552 44878
rect 270500 44814 270552 44820
rect 269120 13116 269172 13122
rect 269120 13058 269172 13064
rect 270408 13116 270460 13122
rect 270408 13058 270460 13064
rect 269132 3346 269160 13058
rect 270512 3602 270540 44814
rect 270592 25560 270644 25566
rect 270592 25502 270644 25508
rect 270500 3596 270552 3602
rect 270500 3538 270552 3544
rect 270604 3482 270632 25502
rect 271696 3596 271748 3602
rect 271696 3538 271748 3544
rect 270512 3454 270632 3482
rect 267752 3318 268148 3346
rect 269132 3318 269344 3346
rect 268120 480 268148 3318
rect 269316 480 269344 3318
rect 270512 480 270540 3454
rect 271708 480 271736 3538
rect 271892 3346 271920 188294
rect 273180 6254 273208 192086
rect 273364 189106 273392 192100
rect 274192 189786 274220 192100
rect 274180 189780 274232 189786
rect 274180 189722 274232 189728
rect 275020 189446 275048 192100
rect 275008 189440 275060 189446
rect 275008 189382 275060 189388
rect 273352 189100 273404 189106
rect 273352 189042 273404 189048
rect 274548 189100 274600 189106
rect 274548 189042 274600 189048
rect 274560 43450 274588 189042
rect 275848 178702 275876 192100
rect 276690 192086 277348 192114
rect 275928 189440 275980 189446
rect 275928 189382 275980 189388
rect 275836 178696 275888 178702
rect 275836 178638 275888 178644
rect 274640 47592 274692 47598
rect 274640 47534 274692 47540
rect 274548 43444 274600 43450
rect 274548 43386 274600 43392
rect 273260 31136 273312 31142
rect 273260 31078 273312 31084
rect 273168 6248 273220 6254
rect 273168 6190 273220 6196
rect 273272 3346 273300 31078
rect 274652 3346 274680 47534
rect 275940 4894 275968 189382
rect 277320 35290 277348 192086
rect 277504 189378 277532 192100
rect 278346 192086 278636 192114
rect 277492 189372 277544 189378
rect 277492 189314 277544 189320
rect 278608 44878 278636 192086
rect 278688 189372 278740 189378
rect 278688 189314 278740 189320
rect 278596 44872 278648 44878
rect 278596 44814 278648 44820
rect 277308 35284 277360 35290
rect 277308 35226 277360 35232
rect 277400 32496 277452 32502
rect 277400 32438 277452 32444
rect 276480 6180 276532 6186
rect 276480 6122 276532 6128
rect 275928 4888 275980 4894
rect 275928 4830 275980 4836
rect 271892 3318 272932 3346
rect 273272 3318 274128 3346
rect 274652 3318 275324 3346
rect 272904 480 272932 3318
rect 274100 480 274128 3318
rect 275296 480 275324 3318
rect 276492 480 276520 6122
rect 277412 3482 277440 32438
rect 278700 21486 278728 189314
rect 279160 189106 279188 192100
rect 280002 192086 280108 192114
rect 280830 192086 281488 192114
rect 279148 189100 279200 189106
rect 279148 189042 279200 189048
rect 279976 189100 280028 189106
rect 279976 189042 280028 189048
rect 279988 71058 280016 189042
rect 279976 71052 280028 71058
rect 279976 70994 280028 71000
rect 278780 50380 278832 50386
rect 278780 50322 278832 50328
rect 278688 21480 278740 21486
rect 278688 21422 278740 21428
rect 278792 3482 278820 50322
rect 280080 22778 280108 192086
rect 280804 189780 280856 189786
rect 280804 189722 280856 189728
rect 280816 33794 280844 189722
rect 281460 47598 281488 192086
rect 281644 190194 281672 192100
rect 282486 192086 282868 192114
rect 281632 190188 281684 190194
rect 281632 190130 281684 190136
rect 282736 190188 282788 190194
rect 282736 190130 282788 190136
rect 282748 73846 282776 190130
rect 282736 73840 282788 73846
rect 282736 73782 282788 73788
rect 281540 51740 281592 51746
rect 281540 51682 281592 51688
rect 281448 47592 281500 47598
rect 281448 47534 281500 47540
rect 280160 33788 280212 33794
rect 280160 33730 280212 33736
rect 280804 33788 280856 33794
rect 280804 33730 280856 33736
rect 280068 22772 280120 22778
rect 280068 22714 280120 22720
rect 280068 4820 280120 4826
rect 280068 4762 280120 4768
rect 277412 3454 277716 3482
rect 278792 3454 278912 3482
rect 277688 480 277716 3454
rect 278884 480 278912 3454
rect 280080 480 280108 4762
rect 280172 3482 280200 33730
rect 281552 3482 281580 51682
rect 282840 24138 282868 192086
rect 283300 189174 283328 192100
rect 284142 192086 284248 192114
rect 284970 192086 285628 192114
rect 283288 189168 283340 189174
rect 283288 189110 283340 189116
rect 284116 189168 284168 189174
rect 284116 189110 284168 189116
rect 284128 49026 284156 189110
rect 284116 49020 284168 49026
rect 284116 48962 284168 48968
rect 284220 36582 284248 192086
rect 284300 46232 284352 46238
rect 284300 46174 284352 46180
rect 284208 36576 284260 36582
rect 284208 36518 284260 36524
rect 282828 24132 282880 24138
rect 282828 24074 282880 24080
rect 282920 17264 282972 17270
rect 282920 17206 282972 17212
rect 282932 3482 282960 17206
rect 284312 3482 284340 46174
rect 285600 17270 285628 192086
rect 285784 189514 285812 192100
rect 286626 192086 286916 192114
rect 285772 189508 285824 189514
rect 285772 189450 285824 189456
rect 286888 76566 286916 192086
rect 286968 189508 287020 189514
rect 286968 189450 287020 189456
rect 286876 76560 286928 76566
rect 286876 76502 286928 76508
rect 285680 53100 285732 53106
rect 285680 53042 285732 53048
rect 285588 17264 285640 17270
rect 285588 17206 285640 17212
rect 285692 3482 285720 53042
rect 286980 46238 287008 189450
rect 287440 189106 287468 192100
rect 287428 189100 287480 189106
rect 287428 189042 287480 189048
rect 288268 50386 288296 192100
rect 289110 192086 289768 192114
rect 288348 189100 288400 189106
rect 288348 189042 288400 189048
rect 288256 50380 288308 50386
rect 288256 50322 288308 50328
rect 286968 46232 287020 46238
rect 286968 46174 287020 46180
rect 287060 26920 287112 26926
rect 287060 26862 287112 26868
rect 287072 3534 287100 26862
rect 288360 14482 288388 189042
rect 289740 77994 289768 192086
rect 289924 189106 289952 192100
rect 290766 192086 291056 192114
rect 289912 189100 289964 189106
rect 289912 189042 289964 189048
rect 289728 77988 289780 77994
rect 289728 77930 289780 77936
rect 288440 54528 288492 54534
rect 288440 54470 288492 54476
rect 287152 14476 287204 14482
rect 287152 14418 287204 14424
rect 288348 14476 288400 14482
rect 288348 14418 288400 14424
rect 287060 3528 287112 3534
rect 280172 3454 281304 3482
rect 281552 3454 282500 3482
rect 282932 3454 283696 3482
rect 284312 3454 284800 3482
rect 285692 3454 285996 3482
rect 287060 3470 287112 3476
rect 281276 480 281304 3454
rect 282472 480 282500 3454
rect 283668 480 283696 3454
rect 284772 480 284800 3454
rect 285968 480 285996 3454
rect 287164 480 287192 14418
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288452 3482 288480 54470
rect 291028 51746 291056 192086
rect 291580 189106 291608 192100
rect 292330 192086 292528 192114
rect 291108 189100 291160 189106
rect 291108 189042 291160 189048
rect 291568 189100 291620 189106
rect 291568 189042 291620 189048
rect 292396 189100 292448 189106
rect 292396 189042 292448 189048
rect 291016 51740 291068 51746
rect 291016 51682 291068 51688
rect 291120 7614 291148 189042
rect 292408 79354 292436 189042
rect 292396 79348 292448 79354
rect 292396 79290 292448 79296
rect 291200 35216 291252 35222
rect 291200 35158 291252 35164
rect 290740 7608 290792 7614
rect 290740 7550 290792 7556
rect 291108 7608 291160 7614
rect 291108 7550 291160 7556
rect 288360 480 288388 3470
rect 288452 3454 289584 3482
rect 289556 480 289584 3454
rect 290752 480 290780 7550
rect 291212 3482 291240 35158
rect 292500 25566 292528 192086
rect 293144 189106 293172 192100
rect 293972 189446 294000 192100
rect 294800 189786 294828 192100
rect 295628 190398 295656 192100
rect 296470 192086 296668 192114
rect 297298 192086 298048 192114
rect 295616 190392 295668 190398
rect 295616 190334 295668 190340
rect 296536 190392 296588 190398
rect 296536 190334 296588 190340
rect 294788 189780 294840 189786
rect 294788 189722 294840 189728
rect 293960 189440 294012 189446
rect 293960 189382 294012 189388
rect 295248 189440 295300 189446
rect 295248 189382 295300 189388
rect 293132 189100 293184 189106
rect 293132 189042 293184 189048
rect 293868 189100 293920 189106
rect 293868 189042 293920 189048
rect 292580 57248 292632 57254
rect 292580 57190 292632 57196
rect 292488 25560 292540 25566
rect 292488 25502 292540 25508
rect 292592 3482 292620 57190
rect 293880 53106 293908 189042
rect 295260 80714 295288 189382
rect 295248 80708 295300 80714
rect 295248 80650 295300 80656
rect 296548 54534 296576 190334
rect 296536 54528 296588 54534
rect 296536 54470 296588 54476
rect 293868 53100 293920 53106
rect 293868 53042 293920 53048
rect 296640 39438 296668 192086
rect 296720 186992 296772 186998
rect 296720 186934 296772 186940
rect 296628 39432 296680 39438
rect 296628 39374 296680 39380
rect 295340 36644 295392 36650
rect 295340 36586 295392 36592
rect 293960 18624 294012 18630
rect 293960 18566 294012 18572
rect 293972 3482 294000 18566
rect 295352 3482 295380 36586
rect 296732 3534 296760 186934
rect 296812 29640 296864 29646
rect 296812 29582 296864 29588
rect 296720 3528 296772 3534
rect 291212 3454 291976 3482
rect 292592 3454 293172 3482
rect 293972 3454 294368 3482
rect 295352 3454 295564 3482
rect 296720 3470 296772 3476
rect 291948 480 291976 3454
rect 293144 480 293172 3454
rect 294340 480 294368 3454
rect 295536 480 295564 3454
rect 296824 1442 296852 29582
rect 298020 26926 298048 192086
rect 298112 189106 298140 192100
rect 298954 192086 299336 192114
rect 298100 189100 298152 189106
rect 298100 189042 298152 189048
rect 299308 82142 299336 192086
rect 299768 189378 299796 192100
rect 300610 192086 300716 192114
rect 299756 189372 299808 189378
rect 299756 189314 299808 189320
rect 299388 189100 299440 189106
rect 299388 189042 299440 189048
rect 299296 82136 299348 82142
rect 299296 82078 299348 82084
rect 299400 55962 299428 189042
rect 299480 58676 299532 58682
rect 299480 58618 299532 58624
rect 299388 55956 299440 55962
rect 299388 55898 299440 55904
rect 298100 28280 298152 28286
rect 298100 28222 298152 28228
rect 298008 26920 298060 26926
rect 298008 26862 298060 26868
rect 297916 3528 297968 3534
rect 297916 3470 297968 3476
rect 298112 3482 298140 28222
rect 299492 3482 299520 58618
rect 300688 57254 300716 192086
rect 300768 189372 300820 189378
rect 300768 189314 300820 189320
rect 300676 57248 300728 57254
rect 300676 57190 300728 57196
rect 300780 15910 300808 189314
rect 301424 189106 301452 192100
rect 301504 189848 301556 189854
rect 301504 189790 301556 189796
rect 301412 189100 301464 189106
rect 301412 189042 301464 189048
rect 301516 19310 301544 189790
rect 302252 189310 302280 192100
rect 303094 192086 303476 192114
rect 302240 189304 302292 189310
rect 302240 189246 302292 189252
rect 302148 189100 302200 189106
rect 302148 189042 302200 189048
rect 302160 83502 302188 189042
rect 302148 83496 302200 83502
rect 302148 83438 302200 83444
rect 303448 58682 303476 192086
rect 303908 190398 303936 192100
rect 304750 192086 304948 192114
rect 305578 192086 306328 192114
rect 303896 190392 303948 190398
rect 303896 190334 303948 190340
rect 304816 190392 304868 190398
rect 304816 190334 304868 190340
rect 303528 189304 303580 189310
rect 303528 189246 303580 189252
rect 303436 58676 303488 58682
rect 303436 58618 303488 58624
rect 302240 37936 302292 37942
rect 302240 37878 302292 37884
rect 301504 19304 301556 19310
rect 301504 19246 301556 19252
rect 300860 15972 300912 15978
rect 300860 15914 300912 15920
rect 300768 15904 300820 15910
rect 300768 15846 300820 15852
rect 300872 3482 300900 15914
rect 302252 3482 302280 37878
rect 303540 28286 303568 189246
rect 304828 84862 304856 190334
rect 304816 84856 304868 84862
rect 304816 84798 304868 84804
rect 303620 60036 303672 60042
rect 303620 59978 303672 59984
rect 303528 28280 303580 28286
rect 303528 28222 303580 28228
rect 303632 3482 303660 59978
rect 304920 29646 304948 192086
rect 305000 177336 305052 177342
rect 305000 177278 305052 177284
rect 304908 29640 304960 29646
rect 304908 29582 304960 29588
rect 305012 3534 305040 177278
rect 306300 61402 306328 192086
rect 306392 189310 306420 192100
rect 306380 189304 306432 189310
rect 306380 189246 306432 189252
rect 307220 189174 307248 192100
rect 307668 189304 307720 189310
rect 307668 189246 307720 189252
rect 307208 189168 307260 189174
rect 307208 189110 307260 189116
rect 307680 113830 307708 189246
rect 308048 189106 308076 192100
rect 308890 192086 309088 192114
rect 308036 189100 308088 189106
rect 308036 189042 308088 189048
rect 308956 189100 309008 189106
rect 308956 189042 309008 189048
rect 307668 113824 307720 113830
rect 307668 113766 307720 113772
rect 306380 62824 306432 62830
rect 306380 62766 306432 62772
rect 306288 61396 306340 61402
rect 306288 61338 306340 61344
rect 305092 19304 305144 19310
rect 305092 19246 305144 19252
rect 305000 3528 305052 3534
rect 296732 1414 296852 1442
rect 296732 480 296760 1414
rect 297928 480 297956 3470
rect 298112 3454 299152 3482
rect 299492 3454 300348 3482
rect 300872 3454 301452 3482
rect 302252 3454 302648 3482
rect 303632 3454 303844 3482
rect 305000 3470 305052 3476
rect 299124 480 299152 3454
rect 300320 480 300348 3454
rect 301424 480 301452 3454
rect 302620 480 302648 3454
rect 303816 480 303844 3454
rect 305104 1442 305132 19246
rect 306196 3528 306248 3534
rect 306196 3470 306248 3476
rect 305012 1414 305132 1442
rect 305012 480 305040 1414
rect 306208 480 306236 3470
rect 306392 3346 306420 62766
rect 308968 60042 308996 189042
rect 308956 60036 309008 60042
rect 308956 59978 309008 59984
rect 308588 8968 308640 8974
rect 308588 8910 308640 8916
rect 306392 3318 307432 3346
rect 307404 480 307432 3318
rect 308600 480 308628 8910
rect 309060 4826 309088 192086
rect 309704 189718 309732 192100
rect 309692 189712 309744 189718
rect 309692 189654 309744 189660
rect 310428 189712 310480 189718
rect 310428 189654 310480 189660
rect 309784 189168 309836 189174
rect 309784 189110 309836 189116
rect 309140 39364 309192 39370
rect 309140 39306 309192 39312
rect 309048 4820 309100 4826
rect 309048 4762 309100 4768
rect 309152 3346 309180 39306
rect 309796 8974 309824 189110
rect 310440 18630 310468 189654
rect 310532 189310 310560 192100
rect 311374 192086 311756 192114
rect 310520 189304 310572 189310
rect 310520 189246 310572 189252
rect 311728 117978 311756 192086
rect 312188 189310 312216 192100
rect 313030 192086 313136 192114
rect 313858 192086 314516 192114
rect 311808 189304 311860 189310
rect 311808 189246 311860 189252
rect 312176 189304 312228 189310
rect 312176 189246 312228 189252
rect 311716 117972 311768 117978
rect 311716 117914 311768 117920
rect 310520 64184 310572 64190
rect 310520 64126 310572 64132
rect 310428 18624 310480 18630
rect 310428 18566 310480 18572
rect 309784 8968 309836 8974
rect 309784 8910 309836 8916
rect 310532 3346 310560 64126
rect 311820 6186 311848 189246
rect 313108 134570 313136 192086
rect 313188 189304 313240 189310
rect 313188 189246 313240 189252
rect 313096 134564 313148 134570
rect 313096 134506 313148 134512
rect 313200 11762 313228 189246
rect 314488 177342 314516 192086
rect 314476 177336 314528 177342
rect 314476 177278 314528 177284
rect 313280 40724 313332 40730
rect 313280 40666 313332 40672
rect 311900 11756 311952 11762
rect 311900 11698 311952 11704
rect 313188 11756 313240 11762
rect 313188 11698 313240 11704
rect 311808 6180 311860 6186
rect 311808 6122 311860 6128
rect 311912 3346 311940 11698
rect 309152 3318 309824 3346
rect 310532 3318 311020 3346
rect 311912 3318 312216 3346
rect 309796 480 309824 3318
rect 310992 480 311020 3318
rect 312188 480 312216 3318
rect 313292 1578 313320 40666
rect 314580 32434 314608 192100
rect 315422 192086 315988 192114
rect 315960 42090 315988 192086
rect 316236 190126 316264 192100
rect 317078 192086 317368 192114
rect 316224 190120 316276 190126
rect 316224 190062 316276 190068
rect 317236 190120 317288 190126
rect 317236 190062 317288 190068
rect 317248 86290 317276 190062
rect 317236 86284 317288 86290
rect 317236 86226 317288 86232
rect 316040 42152 316092 42158
rect 316040 42094 316092 42100
rect 315948 42084 316000 42090
rect 315948 42026 316000 42032
rect 313372 32428 313424 32434
rect 313372 32370 313424 32376
rect 314568 32428 314620 32434
rect 314568 32370 314620 32376
rect 313384 3534 313412 32370
rect 314660 19984 314712 19990
rect 314660 19926 314712 19932
rect 313372 3528 313424 3534
rect 313372 3470 313424 3476
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 313292 1550 313412 1578
rect 313384 480 313412 1550
rect 314580 480 314608 3470
rect 314672 3346 314700 19926
rect 316052 3482 316080 42094
rect 317340 19990 317368 192086
rect 317892 189446 317920 192100
rect 318628 192086 318734 192114
rect 319562 192086 320128 192114
rect 317880 189440 317932 189446
rect 317880 189382 317932 189388
rect 318628 89010 318656 192086
rect 318708 189440 318760 189446
rect 318708 189382 318760 189388
rect 318616 89004 318668 89010
rect 318616 88946 318668 88952
rect 317420 65544 317472 65550
rect 317420 65486 317472 65492
rect 317328 19984 317380 19990
rect 317328 19926 317380 19932
rect 317432 3482 317460 65486
rect 318720 62830 318748 189382
rect 318708 62824 318760 62830
rect 318708 62766 318760 62772
rect 320100 10334 320128 192086
rect 320376 190330 320404 192100
rect 321218 192086 321508 192114
rect 320364 190324 320416 190330
rect 320364 190266 320416 190272
rect 321376 190324 321428 190330
rect 321376 190266 321428 190272
rect 321388 108322 321416 190266
rect 321376 108316 321428 108322
rect 321376 108258 321428 108264
rect 321480 90370 321508 192086
rect 322032 189514 322060 192100
rect 322768 192086 322874 192114
rect 323702 192086 324268 192114
rect 322020 189508 322072 189514
rect 322020 189450 322072 189456
rect 321468 90364 321520 90370
rect 321468 90306 321520 90312
rect 321560 66904 321612 66910
rect 321560 66846 321612 66852
rect 320180 31068 320232 31074
rect 320180 31010 320232 31016
rect 318800 10328 318852 10334
rect 318800 10270 318852 10276
rect 320088 10328 320140 10334
rect 320088 10270 320140 10276
rect 318812 3482 318840 10270
rect 320192 3482 320220 31010
rect 321572 3482 321600 66846
rect 322768 65550 322796 192086
rect 322848 189508 322900 189514
rect 322848 189450 322900 189456
rect 322756 65544 322808 65550
rect 322756 65486 322808 65492
rect 322860 13122 322888 189450
rect 322940 188352 322992 188358
rect 322940 188294 322992 188300
rect 321652 13116 321704 13122
rect 321652 13058 321704 13064
rect 322848 13116 322900 13122
rect 322848 13058 322900 13064
rect 321664 3602 321692 13058
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 316052 3454 317000 3482
rect 317432 3454 318104 3482
rect 318812 3454 319300 3482
rect 320192 3454 320496 3482
rect 321572 3454 321692 3482
rect 314672 3318 315804 3346
rect 315776 480 315804 3318
rect 316972 480 317000 3454
rect 318076 480 318104 3454
rect 319272 480 319300 3454
rect 320468 480 320496 3454
rect 321664 480 321692 3454
rect 322860 480 322888 3538
rect 322952 3482 322980 188294
rect 324240 91798 324268 192086
rect 324516 189106 324544 192100
rect 325358 192086 325648 192114
rect 326186 192086 326936 192114
rect 324504 189100 324556 189106
rect 324504 189042 324556 189048
rect 324228 91792 324280 91798
rect 324228 91734 324280 91740
rect 324320 68332 324372 68338
rect 324320 68274 324372 68280
rect 324332 3482 324360 68274
rect 325620 66910 325648 192086
rect 326908 104174 326936 192086
rect 326896 104168 326948 104174
rect 326896 104110 326948 104116
rect 325608 66904 325660 66910
rect 325608 66846 325660 66852
rect 327000 31074 327028 192100
rect 327842 192086 328408 192114
rect 327724 189100 327776 189106
rect 327724 189042 327776 189048
rect 327080 43444 327132 43450
rect 327080 43386 327132 43392
rect 326988 31068 327040 31074
rect 326988 31010 327040 31016
rect 326436 6248 326488 6254
rect 326436 6190 326488 6196
rect 322952 3454 324084 3482
rect 324332 3454 325280 3482
rect 324056 480 324084 3454
rect 325252 480 325280 3454
rect 326448 480 326476 6190
rect 327092 3482 327120 43386
rect 327736 35222 327764 189042
rect 328380 68338 328408 192086
rect 328656 190330 328684 192100
rect 329498 192086 329788 192114
rect 328644 190324 328696 190330
rect 328644 190266 328696 190272
rect 329656 190324 329708 190330
rect 329656 190266 329708 190272
rect 329668 93158 329696 190266
rect 329656 93152 329708 93158
rect 329656 93094 329708 93100
rect 328368 68332 328420 68338
rect 328368 68274 328420 68280
rect 327724 35216 327776 35222
rect 327724 35158 327776 35164
rect 329760 33794 329788 192086
rect 330312 189514 330340 192100
rect 331048 192086 331154 192114
rect 331982 192086 332548 192114
rect 330300 189508 330352 189514
rect 330300 189450 330352 189456
rect 331048 109750 331076 192086
rect 331128 189508 331180 189514
rect 331128 189450 331180 189456
rect 331036 109744 331088 109750
rect 331036 109686 331088 109692
rect 331140 69698 331168 189450
rect 331220 178696 331272 178702
rect 331220 178638 331272 178644
rect 331128 69692 331180 69698
rect 331128 69634 331180 69640
rect 328460 33788 328512 33794
rect 328460 33730 328512 33736
rect 329748 33788 329800 33794
rect 329748 33730 329800 33736
rect 328472 3482 328500 33730
rect 330024 4888 330076 4894
rect 330024 4830 330076 4836
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330036 480 330064 4830
rect 331232 480 331260 178638
rect 331312 35284 331364 35290
rect 331312 35226 331364 35232
rect 331324 3482 331352 35226
rect 332520 21418 332548 192086
rect 332796 190262 332824 192100
rect 333638 192086 333836 192114
rect 332784 190256 332836 190262
rect 332784 190198 332836 190204
rect 333808 94518 333836 192086
rect 333888 190256 333940 190262
rect 333888 190198 333940 190204
rect 333796 94512 333848 94518
rect 333796 94454 333848 94460
rect 333900 72486 333928 190198
rect 334452 189718 334480 192100
rect 335188 192086 335294 192114
rect 336122 192086 336688 192114
rect 334440 189712 334492 189718
rect 334440 189654 334492 189660
rect 335188 75206 335216 192086
rect 335268 189712 335320 189718
rect 335268 189654 335320 189660
rect 335176 75200 335228 75206
rect 335176 75142 335228 75148
rect 333888 72480 333940 72486
rect 333888 72422 333940 72428
rect 333980 44872 334032 44878
rect 333980 44814 334032 44820
rect 332600 21480 332652 21486
rect 332600 21422 332652 21428
rect 332508 21412 332560 21418
rect 332508 21354 332560 21360
rect 332612 3482 332640 21422
rect 333992 3482 334020 44814
rect 335280 37942 335308 189654
rect 336660 95946 336688 192086
rect 336936 189310 336964 192100
rect 337686 192086 337976 192114
rect 336924 189304 336976 189310
rect 336924 189246 336976 189252
rect 336648 95940 336700 95946
rect 336648 95882 336700 95888
rect 335360 71052 335412 71058
rect 335360 70994 335412 71000
rect 335268 37936 335320 37942
rect 335268 37878 335320 37884
rect 335372 3482 335400 70994
rect 337948 44878 337976 192086
rect 338028 189304 338080 189310
rect 338028 189246 338080 189252
rect 337936 44872 337988 44878
rect 337936 44814 337988 44820
rect 338040 22778 338068 189246
rect 338500 189106 338528 192100
rect 339342 192086 339448 192114
rect 340170 192086 340828 192114
rect 338488 189100 338540 189106
rect 338488 189042 338540 189048
rect 339316 189100 339368 189106
rect 339316 189042 339368 189048
rect 339328 101454 339356 189042
rect 339316 101448 339368 101454
rect 339316 101390 339368 101396
rect 338120 47592 338172 47598
rect 338120 47534 338172 47540
rect 336740 22772 336792 22778
rect 336740 22714 336792 22720
rect 338028 22772 338080 22778
rect 338028 22714 338080 22720
rect 336752 3482 336780 22714
rect 338132 3482 338160 47534
rect 339420 40730 339448 192086
rect 339500 73840 339552 73846
rect 339500 73782 339552 73788
rect 339408 40724 339460 40730
rect 339408 40666 339460 40672
rect 331324 3454 332456 3482
rect 332612 3454 333652 3482
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 332428 480 332456 3454
rect 333624 480 333652 3454
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339512 480 339540 73782
rect 340800 47598 340828 192086
rect 340984 189990 341012 192100
rect 341826 192086 342208 192114
rect 340972 189984 341024 189990
rect 340972 189926 341024 189932
rect 342076 189984 342128 189990
rect 342076 189926 342128 189932
rect 342088 97306 342116 189926
rect 342076 97300 342128 97306
rect 342076 97242 342128 97248
rect 340880 49020 340932 49026
rect 340880 48962 340932 48968
rect 340788 47592 340840 47598
rect 340788 47534 340840 47540
rect 339592 24132 339644 24138
rect 339592 24074 339644 24080
rect 339604 3482 339632 24074
rect 340892 3482 340920 48962
rect 342180 24138 342208 192086
rect 342640 189106 342668 192100
rect 343482 192086 343588 192114
rect 344310 192086 344968 192114
rect 342628 189100 342680 189106
rect 342628 189042 342680 189048
rect 343560 98666 343588 192086
rect 344284 189100 344336 189106
rect 344284 189042 344336 189048
rect 343548 98660 343600 98666
rect 343548 98602 343600 98608
rect 344296 49026 344324 189042
rect 344284 49020 344336 49026
rect 344284 48962 344336 48968
rect 342260 36576 342312 36582
rect 342260 36518 342312 36524
rect 342168 24132 342220 24138
rect 342168 24074 342220 24080
rect 342272 3482 342300 36518
rect 344940 17270 344968 192086
rect 345124 189310 345152 192100
rect 345966 192086 346256 192114
rect 345112 189304 345164 189310
rect 345112 189246 345164 189252
rect 346228 100026 346256 192086
rect 346780 189446 346808 192100
rect 346768 189440 346820 189446
rect 346768 189382 346820 189388
rect 346308 189304 346360 189310
rect 346308 189246 346360 189252
rect 346216 100020 346268 100026
rect 346216 99962 346268 99968
rect 346320 46238 346348 189246
rect 346400 76560 346452 76566
rect 346400 76502 346452 76508
rect 345020 46232 345072 46238
rect 345020 46174 345072 46180
rect 346308 46232 346360 46238
rect 346308 46174 346360 46180
rect 343640 17264 343692 17270
rect 343640 17206 343692 17212
rect 344928 17264 344980 17270
rect 344928 17206 344980 17212
rect 343652 3482 343680 17206
rect 345032 3482 345060 46174
rect 346412 3482 346440 76502
rect 347608 71058 347636 192100
rect 348450 192086 349108 192114
rect 347688 189440 347740 189446
rect 347688 189382 347740 189388
rect 347596 71052 347648 71058
rect 347596 70994 347648 71000
rect 347700 43450 347728 189382
rect 349080 76566 349108 192086
rect 349264 189378 349292 192100
rect 350106 192086 350396 192114
rect 349252 189372 349304 189378
rect 349252 189314 349304 189320
rect 349160 77988 349212 77994
rect 349160 77930 349212 77936
rect 349068 76560 349120 76566
rect 349068 76502 349120 76508
rect 347780 50380 347832 50386
rect 347780 50322 347832 50328
rect 347688 43444 347740 43450
rect 347688 43386 347740 43392
rect 347792 3534 347820 50322
rect 347872 14476 347924 14482
rect 347872 14418 347924 14424
rect 347780 3528 347832 3534
rect 339604 3454 340736 3482
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 343652 3454 344324 3482
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 347780 3470 347832 3476
rect 340708 480 340736 3454
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 3454
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 14418
rect 349068 3528 349120 3534
rect 349068 3470 349120 3476
rect 349172 3482 349200 77930
rect 350368 50386 350396 192086
rect 350448 189372 350500 189378
rect 350448 189314 350500 189320
rect 350356 50380 350408 50386
rect 350356 50322 350408 50328
rect 350460 14482 350488 189314
rect 350920 189106 350948 192100
rect 351762 192086 351868 192114
rect 352590 192086 353248 192114
rect 350908 189100 350960 189106
rect 350908 189042 350960 189048
rect 351736 189100 351788 189106
rect 351736 189042 351788 189048
rect 351748 102814 351776 189042
rect 351736 102808 351788 102814
rect 351736 102750 351788 102756
rect 351840 36582 351868 192086
rect 352564 189780 352616 189786
rect 352564 189722 352616 189728
rect 351920 51740 351972 51746
rect 351920 51682 351972 51688
rect 351828 36576 351880 36582
rect 351828 36518 351880 36524
rect 350448 14476 350500 14482
rect 350448 14418 350500 14424
rect 351368 7608 351420 7614
rect 351368 7550 351420 7556
rect 349080 480 349108 3470
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 7550
rect 351932 3618 351960 51682
rect 352576 4894 352604 189722
rect 353220 51746 353248 192086
rect 353404 190126 353432 192100
rect 354246 192086 354628 192114
rect 353392 190120 353444 190126
rect 353392 190062 353444 190068
rect 354496 190120 354548 190126
rect 354496 190062 354548 190068
rect 354508 105602 354536 190062
rect 354496 105596 354548 105602
rect 354496 105538 354548 105544
rect 353300 79348 353352 79354
rect 353300 79290 353352 79296
rect 353208 51740 353260 51746
rect 353208 51682 353260 51688
rect 352564 4888 352616 4894
rect 352564 4830 352616 4836
rect 351932 3590 352604 3618
rect 352576 480 352604 3590
rect 353312 3482 353340 79290
rect 354600 7614 354628 192086
rect 355060 190262 355088 192100
rect 355902 192086 356008 192114
rect 356730 192086 357388 192114
rect 355048 190256 355100 190262
rect 355048 190198 355100 190204
rect 355876 190256 355928 190262
rect 355876 190198 355928 190204
rect 355888 73846 355916 190198
rect 355876 73840 355928 73846
rect 355876 73782 355928 73788
rect 354680 25560 354732 25566
rect 354680 25502 354732 25508
rect 354588 7608 354640 7614
rect 354588 7550 354640 7556
rect 353312 3454 353800 3482
rect 353772 480 353800 3454
rect 354692 3346 354720 25502
rect 355980 3466 356008 192086
rect 356060 80708 356112 80714
rect 356060 80650 356112 80656
rect 356072 3534 356100 80650
rect 356152 53100 356204 53106
rect 356152 53042 356204 53048
rect 356060 3528 356112 3534
rect 356060 3470 356112 3476
rect 355968 3460 356020 3466
rect 355968 3402 356020 3408
rect 354692 3318 354996 3346
rect 354968 480 354996 3318
rect 356164 480 356192 53042
rect 357360 39370 357388 192086
rect 357544 189106 357572 192100
rect 358386 192086 358768 192114
rect 357532 189100 357584 189106
rect 357532 189042 357584 189048
rect 358636 189100 358688 189106
rect 358636 189042 358688 189048
rect 358648 53106 358676 189042
rect 358636 53100 358688 53106
rect 358636 53042 358688 53048
rect 357348 39364 357400 39370
rect 357348 39306 357400 39312
rect 358544 4888 358596 4894
rect 358544 4830 358596 4836
rect 357348 3528 357400 3534
rect 357348 3470 357400 3476
rect 357360 480 357388 3470
rect 358556 480 358584 4830
rect 358740 3534 358768 192086
rect 359200 189786 359228 192100
rect 359950 192086 360148 192114
rect 360778 192086 361528 192114
rect 359188 189780 359240 189786
rect 359188 189722 359240 189728
rect 360120 54534 360148 192086
rect 358820 54528 358872 54534
rect 358820 54470 358872 54476
rect 360108 54528 360160 54534
rect 360108 54470 360160 54476
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358832 3346 358860 54470
rect 360200 39432 360252 39438
rect 360200 39374 360252 39380
rect 360212 3346 360240 39374
rect 361500 4146 361528 192086
rect 361592 190058 361620 192100
rect 362434 192086 362908 192114
rect 361580 190052 361632 190058
rect 361580 189994 361632 190000
rect 362776 190052 362828 190058
rect 362776 189994 362828 190000
rect 362788 64190 362816 189994
rect 362776 64184 362828 64190
rect 362776 64126 362828 64132
rect 362880 55894 362908 192086
rect 363248 189106 363276 192100
rect 364090 192086 364196 192114
rect 363236 189100 363288 189106
rect 363236 189042 363288 189048
rect 364168 159390 364196 192086
rect 364904 189718 364932 192100
rect 364892 189712 364944 189718
rect 364892 189654 364944 189660
rect 365628 189712 365680 189718
rect 365628 189654 365680 189660
rect 364248 189100 364300 189106
rect 364248 189042 364300 189048
rect 364156 159384 364208 159390
rect 364156 159326 364208 159332
rect 362960 55956 363012 55962
rect 362960 55898 363012 55904
rect 362868 55888 362920 55894
rect 362868 55830 362920 55836
rect 361580 26920 361632 26926
rect 361580 26862 361632 26868
rect 361488 4140 361540 4146
rect 361488 4082 361540 4088
rect 361592 3346 361620 26862
rect 362972 3346 363000 55898
rect 364260 4010 364288 189042
rect 364340 82136 364392 82142
rect 364340 82078 364392 82084
rect 364248 4004 364300 4010
rect 364248 3946 364300 3952
rect 358832 3318 359780 3346
rect 360212 3318 360976 3346
rect 361592 3318 362172 3346
rect 362972 3318 363368 3346
rect 359752 480 359780 3318
rect 360948 480 360976 3318
rect 362144 480 362172 3318
rect 363340 480 363368 3318
rect 364352 610 364380 82078
rect 365640 80714 365668 189654
rect 365732 189310 365760 192100
rect 366574 192086 366956 192114
rect 365720 189304 365772 189310
rect 365720 189246 365772 189252
rect 366928 158030 366956 192086
rect 367008 189304 367060 189310
rect 367008 189246 367060 189252
rect 366916 158024 366968 158030
rect 366916 157966 366968 157972
rect 365628 80708 365680 80714
rect 365628 80650 365680 80656
rect 365720 57248 365772 57254
rect 365720 57190 365772 57196
rect 365732 3602 365760 57190
rect 365812 15904 365864 15910
rect 365812 15846 365864 15852
rect 365720 3596 365772 3602
rect 365720 3538 365772 3544
rect 365824 3482 365852 15846
rect 367020 4078 367048 189246
rect 367388 181490 367416 192100
rect 368230 192086 368428 192114
rect 369058 192086 369808 192114
rect 367376 181484 367428 181490
rect 367376 181426 367428 181432
rect 367100 83496 367152 83502
rect 367100 83438 367152 83444
rect 367008 4072 367060 4078
rect 367008 4014 367060 4020
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 365732 3454 365852 3482
rect 364340 604 364392 610
rect 364340 546 364392 552
rect 364524 604 364576 610
rect 364524 546 364576 552
rect 364536 480 364564 546
rect 365732 480 365760 3454
rect 366928 480 366956 3538
rect 367112 610 367140 83438
rect 368400 3942 368428 192086
rect 369780 28286 369808 192086
rect 369872 190058 369900 192100
rect 370714 192086 371188 192114
rect 369860 190052 369912 190058
rect 369860 189994 369912 190000
rect 371056 190052 371108 190058
rect 371056 189994 371108 190000
rect 371068 140078 371096 189994
rect 371056 140072 371108 140078
rect 371056 140014 371108 140020
rect 369860 58676 369912 58682
rect 369860 58618 369912 58624
rect 368480 28280 368532 28286
rect 368480 28222 368532 28228
rect 369768 28280 369820 28286
rect 369768 28222 369820 28228
rect 368388 3936 368440 3942
rect 368388 3878 368440 3884
rect 368492 610 368520 28222
rect 369872 610 369900 58618
rect 371160 3874 371188 192086
rect 371528 189378 371556 192100
rect 372370 192086 372476 192114
rect 371516 189372 371568 189378
rect 371516 189314 371568 189320
rect 372448 111110 372476 192086
rect 373184 189990 373212 192100
rect 373172 189984 373224 189990
rect 373172 189926 373224 189932
rect 373908 189984 373960 189990
rect 373908 189926 373960 189932
rect 372528 189372 372580 189378
rect 372528 189314 372580 189320
rect 372436 111104 372488 111110
rect 372436 111046 372488 111052
rect 371240 84856 371292 84862
rect 371240 84798 371292 84804
rect 371148 3868 371200 3874
rect 371148 3810 371200 3816
rect 371252 626 371280 84798
rect 372540 26926 372568 189314
rect 372620 29640 372672 29646
rect 372620 29582 372672 29588
rect 372528 26920 372580 26926
rect 372528 26862 372580 26868
rect 367100 604 367152 610
rect 367100 546 367152 552
rect 368020 604 368072 610
rect 368020 546 368072 552
rect 368480 604 368532 610
rect 368480 546 368532 552
rect 369216 604 369268 610
rect 369216 546 369268 552
rect 369860 604 369912 610
rect 369860 546 369912 552
rect 370412 604 370464 610
rect 371252 598 371648 626
rect 372632 610 372660 29582
rect 373920 3806 373948 189926
rect 374012 189310 374040 192100
rect 374854 192086 375236 192114
rect 374000 189304 374052 189310
rect 374000 189246 374052 189252
rect 375208 138718 375236 192086
rect 375668 189310 375696 192100
rect 376510 192086 376616 192114
rect 377338 192086 378088 192114
rect 375288 189304 375340 189310
rect 375288 189246 375340 189252
rect 375656 189304 375708 189310
rect 375656 189246 375708 189252
rect 375196 138712 375248 138718
rect 375196 138654 375248 138660
rect 374000 113824 374052 113830
rect 374000 113766 374052 113772
rect 373908 3800 373960 3806
rect 373908 3742 373960 3748
rect 374012 3602 374040 113766
rect 375300 87650 375328 189246
rect 376588 156670 376616 192086
rect 376668 189304 376720 189310
rect 376668 189246 376720 189252
rect 376576 156664 376628 156670
rect 376576 156606 376628 156612
rect 375288 87644 375340 87650
rect 375288 87586 375340 87592
rect 374092 61396 374144 61402
rect 374092 61338 374144 61344
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 374104 1578 374132 61338
rect 376392 8968 376444 8974
rect 376392 8910 376444 8916
rect 375196 3596 375248 3602
rect 375196 3538 375248 3544
rect 374012 1550 374132 1578
rect 370412 546 370464 552
rect 368032 480 368060 546
rect 369228 480 369256 546
rect 370424 480 370452 546
rect 371620 480 371648 598
rect 372620 604 372672 610
rect 372620 546 372672 552
rect 372804 604 372856 610
rect 372804 546 372856 552
rect 372816 480 372844 546
rect 374012 480 374040 1550
rect 375208 480 375236 3538
rect 376404 480 376432 8910
rect 376680 3738 376708 189246
rect 376760 60036 376812 60042
rect 376760 59978 376812 59984
rect 376668 3732 376720 3738
rect 376668 3674 376720 3680
rect 376772 3346 376800 59978
rect 378060 57254 378088 192086
rect 378152 189310 378180 192100
rect 378140 189304 378192 189310
rect 378140 189246 378192 189252
rect 378980 189174 379008 192100
rect 379808 190126 379836 192100
rect 380650 192086 380848 192114
rect 379796 190120 379848 190126
rect 379796 190062 379848 190068
rect 380716 190120 380768 190126
rect 380716 190062 380768 190068
rect 379428 189304 379480 189310
rect 379428 189246 379480 189252
rect 378968 189168 379020 189174
rect 378968 189110 379020 189116
rect 378048 57248 378100 57254
rect 378048 57190 378100 57196
rect 378784 4820 378836 4826
rect 378784 4762 378836 4768
rect 376772 3318 377628 3346
rect 377600 480 377628 3318
rect 378796 480 378824 4762
rect 379440 3670 379468 189246
rect 380728 137290 380756 190062
rect 380716 137284 380768 137290
rect 380716 137226 380768 137232
rect 379520 18624 379572 18630
rect 379520 18566 379572 18572
rect 379428 3664 379480 3670
rect 379428 3606 379480 3612
rect 379532 3346 379560 18566
rect 380820 3602 380848 192086
rect 381464 189106 381492 192100
rect 381544 189780 381596 189786
rect 381544 189722 381596 189728
rect 381452 189100 381504 189106
rect 381452 189042 381504 189048
rect 381556 8974 381584 189722
rect 382292 189106 382320 192100
rect 383042 192086 383608 192114
rect 382188 189100 382240 189106
rect 382188 189042 382240 189048
rect 382280 189100 382332 189106
rect 382280 189042 382332 189048
rect 383476 189100 383528 189106
rect 383476 189042 383528 189048
rect 381544 8968 381596 8974
rect 381544 8910 381596 8916
rect 381176 6180 381228 6186
rect 381176 6122 381228 6128
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 379532 3318 380020 3346
rect 379992 480 380020 3318
rect 381188 480 381216 6122
rect 382200 4826 382228 189042
rect 383488 155242 383516 189042
rect 383476 155236 383528 155242
rect 383476 155178 383528 155184
rect 382280 117972 382332 117978
rect 382280 117914 382332 117920
rect 382188 4820 382240 4826
rect 382188 4762 382240 4768
rect 382292 1578 382320 117914
rect 383580 58682 383608 192086
rect 383856 189786 383884 192100
rect 384698 192086 384988 192114
rect 383844 189780 383896 189786
rect 383844 189722 383896 189728
rect 384304 189168 384356 189174
rect 384304 189110 384356 189116
rect 384316 134570 384344 189110
rect 384960 153882 384988 192086
rect 385512 189106 385540 192100
rect 385500 189100 385552 189106
rect 385500 189042 385552 189048
rect 386236 189100 386288 189106
rect 386236 189042 386288 189048
rect 385040 177336 385092 177342
rect 385040 177278 385092 177284
rect 384948 153876 385000 153882
rect 384948 153818 385000 153824
rect 383660 134564 383712 134570
rect 383660 134506 383712 134512
rect 384304 134564 384356 134570
rect 384304 134506 384356 134512
rect 383568 58676 383620 58682
rect 383568 58618 383620 58624
rect 382372 11756 382424 11762
rect 382372 11698 382424 11704
rect 382384 3398 382412 11698
rect 383672 3482 383700 134506
rect 385052 3482 385080 177278
rect 386248 60042 386276 189042
rect 386340 188358 386368 192100
rect 387182 192086 387748 192114
rect 386328 188352 386380 188358
rect 386328 188294 386380 188300
rect 386236 60036 386288 60042
rect 386236 59978 386288 59984
rect 387720 32434 387748 192086
rect 387996 189514 388024 192100
rect 387984 189508 388036 189514
rect 387984 189450 388036 189456
rect 388824 186998 388852 192100
rect 389088 189508 389140 189514
rect 389088 189450 389140 189456
rect 388812 186992 388864 186998
rect 388812 186934 388864 186940
rect 389100 61402 389128 189450
rect 389652 189106 389680 192100
rect 390388 192086 390494 192114
rect 391322 192086 391888 192114
rect 389640 189100 389692 189106
rect 389640 189042 389692 189048
rect 390388 135930 390416 192086
rect 390468 189100 390520 189106
rect 390468 189042 390520 189048
rect 390376 135924 390428 135930
rect 390376 135866 390428 135872
rect 389180 86284 389232 86290
rect 389180 86226 389232 86232
rect 389088 61396 389140 61402
rect 389088 61338 389140 61344
rect 387800 42084 387852 42090
rect 387800 42026 387852 42032
rect 386420 32428 386472 32434
rect 386420 32370 386472 32376
rect 387708 32428 387760 32434
rect 387708 32370 387760 32376
rect 386432 3482 386460 32370
rect 387812 3482 387840 42026
rect 389192 3482 389220 86226
rect 390480 15910 390508 189042
rect 390560 62824 390612 62830
rect 390560 62766 390612 62772
rect 390468 15904 390520 15910
rect 390468 15846 390520 15852
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 386432 3454 387104 3482
rect 387812 3454 388300 3482
rect 389192 3454 389496 3482
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 1550 382412 1578
rect 382384 480 382412 1550
rect 383580 480 383608 3334
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 3454
rect 388272 480 388300 3454
rect 389468 480 389496 3454
rect 390572 3398 390600 62766
rect 390652 19984 390704 19990
rect 390652 19926 390704 19932
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 19926
rect 391860 6186 391888 192086
rect 392136 189106 392164 192100
rect 392978 192086 393268 192114
rect 392124 189100 392176 189106
rect 392124 189042 392176 189048
rect 393136 189100 393188 189106
rect 393136 189042 393188 189048
rect 393148 152522 393176 189042
rect 393136 152516 393188 152522
rect 393136 152458 393188 152464
rect 391940 89004 391992 89010
rect 391940 88946 391992 88952
rect 391848 6180 391900 6186
rect 391848 6122 391900 6128
rect 391952 3482 391980 88946
rect 393240 62830 393268 192086
rect 393792 185638 393820 192100
rect 393780 185632 393832 185638
rect 393780 185574 393832 185580
rect 393228 62824 393280 62830
rect 393228 62766 393280 62772
rect 394620 10334 394648 192100
rect 395462 192086 396028 192114
rect 396000 108322 396028 192086
rect 396276 184210 396304 192100
rect 397118 192086 397408 192114
rect 396264 184204 396316 184210
rect 396264 184146 396316 184152
rect 397380 151094 397408 192086
rect 397932 189582 397960 192100
rect 398668 192086 398774 192114
rect 399602 192086 400168 192114
rect 397920 189576 397972 189582
rect 397920 189518 397972 189524
rect 398668 182850 398696 192086
rect 398748 189576 398800 189582
rect 398748 189518 398800 189524
rect 398656 182844 398708 182850
rect 398656 182786 398708 182792
rect 397368 151088 397420 151094
rect 397368 151030 397420 151036
rect 394700 108316 394752 108322
rect 394700 108258 394752 108264
rect 395988 108316 396040 108322
rect 395988 108258 396040 108264
rect 393320 10328 393372 10334
rect 393320 10270 393372 10276
rect 394608 10328 394660 10334
rect 394608 10270 394660 10276
rect 393332 3482 393360 10270
rect 394712 3482 394740 108258
rect 396080 90364 396132 90370
rect 396080 90306 396132 90312
rect 396092 3482 396120 90306
rect 398760 82142 398788 189518
rect 398748 82136 398800 82142
rect 398748 82078 398800 82084
rect 398840 65544 398892 65550
rect 398840 65486 398892 65492
rect 397460 13116 397512 13122
rect 397460 13058 397512 13064
rect 397472 3482 397500 13058
rect 398852 3482 398880 65486
rect 400140 18630 400168 192086
rect 400416 189310 400444 192100
rect 401258 192086 401456 192114
rect 400404 189304 400456 189310
rect 400404 189246 400456 189252
rect 401428 180130 401456 192086
rect 401508 189304 401560 189310
rect 401508 189246 401560 189252
rect 401416 180124 401468 180130
rect 401416 180066 401468 180072
rect 400220 91792 400272 91798
rect 400220 91734 400272 91740
rect 400128 18624 400180 18630
rect 400128 18566 400180 18572
rect 391952 3454 393084 3482
rect 393332 3454 394280 3482
rect 394712 3454 395476 3482
rect 396092 3454 396672 3482
rect 397472 3454 397868 3482
rect 398852 3454 399064 3482
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 393056 480 393084 3454
rect 394252 480 394280 3454
rect 395448 480 395476 3454
rect 396644 480 396672 3454
rect 397840 480 397868 3454
rect 399036 480 399064 3454
rect 400232 480 400260 91734
rect 401520 79354 401548 189246
rect 402072 189106 402100 192100
rect 402808 192086 402914 192114
rect 403742 192086 404308 192114
rect 402060 189100 402112 189106
rect 402060 189042 402112 189048
rect 402808 133210 402836 192086
rect 402888 189100 402940 189106
rect 402888 189042 402940 189048
rect 402796 133204 402848 133210
rect 402796 133146 402848 133152
rect 401508 79348 401560 79354
rect 401508 79290 401560 79296
rect 401600 66904 401652 66910
rect 401600 66846 401652 66852
rect 400312 35216 400364 35222
rect 400312 35158 400364 35164
rect 400324 3482 400352 35158
rect 401612 3482 401640 66846
rect 402900 35222 402928 189042
rect 402980 104168 403032 104174
rect 402980 104110 403032 104116
rect 402888 35216 402940 35222
rect 402888 35158 402940 35164
rect 402992 3482 403020 104110
rect 404280 11762 404308 192086
rect 404556 189106 404584 192100
rect 405306 192086 405688 192114
rect 404544 189100 404596 189106
rect 404544 189042 404596 189048
rect 405556 189100 405608 189106
rect 405556 189042 405608 189048
rect 405568 149734 405596 189042
rect 405556 149728 405608 149734
rect 405556 149670 405608 149676
rect 405660 65550 405688 192086
rect 406120 189106 406148 192100
rect 406962 192086 407068 192114
rect 407790 192086 408448 192114
rect 406108 189100 406160 189106
rect 406108 189042 406160 189048
rect 406936 189100 406988 189106
rect 406936 189042 406988 189048
rect 406948 178702 406976 189042
rect 406936 178696 406988 178702
rect 406936 178638 406988 178644
rect 405740 68332 405792 68338
rect 405740 68274 405792 68280
rect 405648 65544 405700 65550
rect 405648 65486 405700 65492
rect 404360 31068 404412 31074
rect 404360 31010 404412 31016
rect 404268 11756 404320 11762
rect 404268 11698 404320 11704
rect 404372 3482 404400 31010
rect 405752 3482 405780 68274
rect 407040 31074 407068 192086
rect 407120 93152 407172 93158
rect 407120 93094 407172 93100
rect 407028 31068 407080 31074
rect 407028 31010 407080 31016
rect 407132 3482 407160 93094
rect 408420 68338 408448 192086
rect 408604 190194 408632 192100
rect 409446 192086 409828 192114
rect 408592 190188 408644 190194
rect 408592 190130 408644 190136
rect 409696 190188 409748 190194
rect 409696 190130 409748 190136
rect 409708 177342 409736 190130
rect 409696 177336 409748 177342
rect 409696 177278 409748 177284
rect 408500 69692 408552 69698
rect 408500 69634 408552 69640
rect 408408 68332 408460 68338
rect 408408 68274 408460 68280
rect 408512 4214 408540 69634
rect 409800 33794 409828 192086
rect 410260 189446 410288 192100
rect 410248 189440 410300 189446
rect 410248 189382 410300 189388
rect 411088 175982 411116 192100
rect 411930 192086 412588 192114
rect 411168 189440 411220 189446
rect 411168 189382 411220 189388
rect 411076 175976 411128 175982
rect 411076 175918 411128 175924
rect 409880 109744 409932 109750
rect 409880 109686 409932 109692
rect 408592 33788 408644 33794
rect 408592 33730 408644 33736
rect 409788 33788 409840 33794
rect 409788 33730 409840 33736
rect 408500 4208 408552 4214
rect 408500 4150 408552 4156
rect 408604 3482 408632 33730
rect 409696 4208 409748 4214
rect 409696 4150 409748 4156
rect 400324 3454 401364 3482
rect 401612 3454 402560 3482
rect 402992 3454 403756 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 407132 3454 407344 3482
rect 401336 480 401364 3454
rect 402532 480 402560 3454
rect 403728 480 403756 3454
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407316 480 407344 3454
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 4150
rect 409892 3482 409920 109686
rect 411180 69698 411208 189382
rect 411168 69692 411220 69698
rect 411168 69634 411220 69640
rect 412560 21418 412588 192086
rect 412744 189378 412772 192100
rect 413586 192086 413876 192114
rect 412732 189372 412784 189378
rect 412732 189314 412784 189320
rect 413848 174554 413876 192086
rect 413928 189372 413980 189378
rect 413928 189314 413980 189320
rect 413836 174548 413888 174554
rect 413836 174490 413888 174496
rect 412640 72480 412692 72486
rect 412640 72422 412692 72428
rect 411260 21412 411312 21418
rect 411260 21354 411312 21360
rect 412548 21412 412600 21418
rect 412548 21354 412600 21360
rect 411272 3482 411300 21354
rect 412652 3482 412680 72422
rect 413940 66910 413968 189314
rect 414400 189106 414428 192100
rect 415242 192086 415348 192114
rect 416070 192086 416728 192114
rect 414388 189100 414440 189106
rect 414388 189042 414440 189048
rect 415320 131782 415348 192086
rect 416044 189100 416096 189106
rect 416044 189042 416096 189048
rect 416056 148374 416084 189042
rect 416044 148368 416096 148374
rect 416044 148310 416096 148316
rect 415308 131776 415360 131782
rect 415308 131718 415360 131724
rect 414020 94512 414072 94518
rect 414020 94454 414072 94460
rect 413928 66904 413980 66910
rect 413928 66846 413980 66852
rect 414032 3482 414060 94454
rect 415400 37936 415452 37942
rect 415400 37878 415452 37884
rect 415412 3482 415440 37878
rect 416700 13122 416728 192086
rect 416884 190194 416912 192100
rect 417726 192086 418108 192114
rect 416872 190188 416924 190194
rect 416872 190130 416924 190136
rect 417976 190188 418028 190194
rect 417976 190130 418028 190136
rect 417988 146946 418016 190130
rect 417976 146940 418028 146946
rect 417976 146882 418028 146888
rect 416780 95940 416832 95946
rect 416780 95882 416832 95888
rect 416688 13116 416740 13122
rect 416688 13058 416740 13064
rect 409892 3454 410932 3482
rect 411272 3454 412128 3482
rect 412652 3454 413324 3482
rect 414032 3454 414520 3482
rect 415412 3454 415716 3482
rect 410904 480 410932 3454
rect 412100 480 412128 3454
rect 413296 480 413324 3454
rect 414492 480 414520 3454
rect 415688 480 415716 3454
rect 416792 3398 416820 95882
rect 418080 77994 418108 192086
rect 418540 189174 418568 192100
rect 419382 192086 419488 192114
rect 420210 192086 420868 192114
rect 418528 189168 418580 189174
rect 418528 189110 418580 189116
rect 419356 189168 419408 189174
rect 419356 189110 419408 189116
rect 419368 173194 419396 189110
rect 419356 173188 419408 173194
rect 419356 173130 419408 173136
rect 418068 77988 418120 77994
rect 418068 77930 418120 77936
rect 416872 75200 416924 75206
rect 416872 75142 416924 75148
rect 416780 3392 416832 3398
rect 416780 3334 416832 3340
rect 416884 480 416912 75142
rect 419460 22778 419488 192086
rect 420840 72486 420868 192086
rect 421024 189990 421052 192100
rect 421866 192086 422248 192114
rect 421012 189984 421064 189990
rect 421012 189926 421064 189932
rect 422116 189984 422168 189990
rect 422116 189926 422168 189932
rect 422128 171834 422156 189926
rect 422116 171828 422168 171834
rect 422116 171770 422168 171776
rect 420920 101448 420972 101454
rect 420920 101390 420972 101396
rect 420828 72480 420880 72486
rect 420828 72422 420880 72428
rect 419540 44872 419592 44878
rect 419540 44814 419592 44820
rect 418160 22772 418212 22778
rect 418160 22714 418212 22720
rect 419448 22772 419500 22778
rect 419448 22714 419500 22720
rect 418172 3482 418200 22714
rect 419552 3482 419580 44814
rect 420932 3482 420960 101390
rect 422220 37942 422248 192086
rect 422680 189106 422708 192100
rect 422668 189100 422720 189106
rect 422668 189042 422720 189048
rect 423508 169046 423536 192100
rect 424350 192086 425008 192114
rect 423588 189100 423640 189106
rect 423588 189042 423640 189048
rect 423496 169040 423548 169046
rect 423496 168982 423548 168988
rect 423600 75206 423628 189042
rect 423588 75200 423640 75206
rect 423588 75142 423640 75148
rect 423680 47592 423732 47598
rect 423680 47534 423732 47540
rect 422300 40724 422352 40730
rect 422300 40666 422352 40672
rect 422208 37936 422260 37942
rect 422208 37878 422260 37884
rect 422312 3482 422340 40666
rect 423692 3482 423720 47534
rect 424980 42090 425008 192086
rect 425164 189106 425192 192100
rect 426006 192086 426296 192114
rect 425152 189100 425204 189106
rect 425152 189042 425204 189048
rect 426268 167686 426296 192086
rect 426820 189106 426848 192100
rect 427662 192086 427768 192114
rect 426348 189100 426400 189106
rect 426348 189042 426400 189048
rect 426808 189100 426860 189106
rect 426808 189042 426860 189048
rect 427636 189100 427688 189106
rect 427636 189042 427688 189048
rect 426256 167680 426308 167686
rect 426256 167622 426308 167628
rect 425060 97300 425112 97306
rect 425060 97242 425112 97248
rect 424968 42084 425020 42090
rect 424968 42026 425020 42032
rect 425072 3482 425100 97242
rect 426360 44878 426388 189042
rect 427648 145586 427676 189042
rect 427636 145580 427688 145586
rect 427636 145522 427688 145528
rect 427740 49026 427768 192086
rect 428384 189718 428412 192100
rect 428372 189712 428424 189718
rect 428372 189654 428424 189660
rect 429108 189712 429160 189718
rect 429108 189654 429160 189660
rect 427820 98660 427872 98666
rect 427820 98602 427872 98608
rect 426440 49020 426492 49026
rect 426440 48962 426492 48968
rect 427728 49020 427780 49026
rect 427728 48962 427780 48968
rect 426348 44872 426400 44878
rect 426348 44814 426400 44820
rect 425152 24132 425204 24138
rect 425152 24074 425204 24080
rect 425164 4214 425192 24074
rect 425152 4208 425204 4214
rect 425152 4150 425204 4156
rect 426348 4208 426400 4214
rect 426348 4150 426400 4156
rect 418172 3454 419212 3482
rect 419552 3454 420408 3482
rect 420932 3454 421604 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 425072 3454 425192 3482
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 417988 480 418016 3334
rect 419184 480 419212 3454
rect 420380 480 420408 3454
rect 421576 480 421604 3454
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425164 480 425192 3454
rect 426360 480 426388 4150
rect 426452 3482 426480 48962
rect 427832 3482 427860 98602
rect 429120 19990 429148 189654
rect 429212 189106 429240 192100
rect 430054 192086 430528 192114
rect 429200 189100 429252 189106
rect 429200 189042 429252 189048
rect 430396 189100 430448 189106
rect 430396 189042 430448 189048
rect 430408 144226 430436 189042
rect 430396 144220 430448 144226
rect 430396 144162 430448 144168
rect 430500 83502 430528 192086
rect 430868 189106 430896 192100
rect 431710 192086 431908 192114
rect 432538 192086 433288 192114
rect 430856 189100 430908 189106
rect 430856 189042 430908 189048
rect 431776 189100 431828 189106
rect 431776 189042 431828 189048
rect 431788 166326 431816 189042
rect 431776 166320 431828 166326
rect 431776 166262 431828 166268
rect 430488 83496 430540 83502
rect 430488 83438 430540 83444
rect 430580 46232 430632 46238
rect 430580 46174 430632 46180
rect 429108 19984 429160 19990
rect 429108 19926 429160 19932
rect 429200 17264 429252 17270
rect 429200 17206 429252 17212
rect 429212 3482 429240 17206
rect 430592 3482 430620 46174
rect 431880 24138 431908 192086
rect 433260 130422 433288 192086
rect 433352 190058 433380 192100
rect 434194 192086 434668 192114
rect 433340 190052 433392 190058
rect 433340 189994 433392 190000
rect 434536 190052 434588 190058
rect 434536 189994 434588 190000
rect 434548 164898 434576 189994
rect 434536 164892 434588 164898
rect 434536 164834 434588 164840
rect 433248 130416 433300 130422
rect 433248 130358 433300 130364
rect 431960 100020 432012 100026
rect 431960 99962 432012 99968
rect 431868 24132 431920 24138
rect 431868 24074 431920 24080
rect 431972 3482 432000 99962
rect 433340 71052 433392 71058
rect 433340 70994 433392 71000
rect 426452 3454 427584 3482
rect 427832 3454 428780 3482
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 431972 3454 432368 3482
rect 427556 480 427584 3454
rect 428752 480 428780 3454
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3454
rect 433352 3398 433380 70994
rect 434640 43450 434668 192086
rect 435008 189378 435036 192100
rect 435850 192086 435956 192114
rect 434996 189372 435048 189378
rect 434996 189314 435048 189320
rect 435928 163538 435956 192086
rect 436008 189372 436060 189378
rect 436008 189314 436060 189320
rect 435916 163532 435968 163538
rect 435916 163474 435968 163480
rect 434720 76560 434772 76566
rect 434720 76502 434772 76508
rect 433432 43444 433484 43450
rect 433432 43386 433484 43392
rect 434628 43444 434680 43450
rect 434628 43386 434680 43392
rect 433444 3482 433472 43386
rect 434732 3482 434760 76502
rect 436020 71058 436048 189314
rect 436664 189106 436692 192100
rect 437492 189310 437520 192100
rect 438334 192086 438716 192114
rect 437480 189304 437532 189310
rect 437480 189246 437532 189252
rect 436652 189100 436704 189106
rect 436652 189042 436704 189048
rect 437388 189100 437440 189106
rect 437388 189042 437440 189048
rect 436008 71052 436060 71058
rect 436008 70994 436060 71000
rect 437400 14482 437428 189042
rect 438688 162178 438716 192086
rect 439148 190398 439176 192100
rect 439990 192086 440188 192114
rect 440818 192086 441568 192114
rect 439136 190392 439188 190398
rect 439136 190334 439188 190340
rect 440056 190392 440108 190398
rect 440056 190334 440108 190340
rect 438768 189304 438820 189310
rect 438768 189246 438820 189252
rect 438676 162172 438728 162178
rect 438676 162114 438728 162120
rect 438780 86290 438808 189246
rect 440068 142866 440096 190334
rect 440056 142860 440108 142866
rect 440056 142802 440108 142808
rect 438860 102808 438912 102814
rect 438860 102750 438912 102756
rect 438768 86284 438820 86290
rect 438768 86226 438820 86232
rect 437480 50380 437532 50386
rect 437480 50322 437532 50328
rect 436100 14476 436152 14482
rect 436100 14418 436152 14424
rect 437388 14476 437440 14482
rect 437388 14418 437440 14424
rect 436112 3482 436140 14418
rect 437492 3482 437520 50322
rect 438872 3482 438900 102750
rect 440160 46238 440188 192086
rect 440148 46232 440200 46238
rect 440148 46174 440200 46180
rect 440240 36576 440292 36582
rect 440240 36518 440292 36524
rect 440252 3482 440280 36518
rect 441540 25566 441568 192086
rect 441632 190126 441660 192100
rect 442474 192086 442948 192114
rect 441620 190120 441672 190126
rect 441620 190062 441672 190068
rect 442816 190120 442868 190126
rect 442816 190062 442868 190068
rect 442828 141438 442856 190062
rect 442816 141432 442868 141438
rect 442816 141374 442868 141380
rect 441620 51740 441672 51746
rect 441620 51682 441672 51688
rect 441528 25560 441580 25566
rect 441528 25502 441580 25508
rect 441632 3482 441660 51682
rect 442920 50386 442948 192086
rect 443288 190262 443316 192100
rect 444130 192086 444328 192114
rect 443276 190256 443328 190262
rect 443276 190198 443328 190204
rect 444196 190256 444248 190262
rect 444196 190198 444248 190204
rect 444208 160750 444236 190198
rect 444196 160744 444248 160750
rect 444196 160686 444248 160692
rect 443000 105596 443052 105602
rect 443000 105538 443052 105544
rect 442908 50380 442960 50386
rect 442908 50322 442960 50328
rect 433444 3454 433564 3482
rect 434732 3454 435864 3482
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433536 480 433564 3454
rect 434628 3392 434680 3398
rect 434628 3334 434680 3340
rect 434640 480 434668 3334
rect 435836 480 435864 3454
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 105538
rect 444300 36582 444328 192086
rect 444944 189106 444972 192100
rect 445772 189174 445800 192100
rect 446614 192086 447088 192114
rect 445760 189168 445812 189174
rect 445760 189110 445812 189116
rect 444932 189100 444984 189106
rect 444932 189042 444984 189048
rect 445668 189100 445720 189106
rect 445668 189042 445720 189048
rect 445680 73846 445708 189042
rect 444380 73840 444432 73846
rect 444380 73782 444432 73788
rect 445668 73840 445720 73846
rect 445668 73782 445720 73788
rect 444288 36576 444340 36582
rect 444288 36518 444340 36524
rect 444196 7608 444248 7614
rect 444196 7550 444248 7556
rect 444208 480 444236 7550
rect 444392 3482 444420 73782
rect 447060 47598 447088 192086
rect 447428 189446 447456 192100
rect 448256 189854 448284 192100
rect 449098 192086 449848 192114
rect 448244 189848 448296 189854
rect 448244 189790 448296 189796
rect 447416 189440 447468 189446
rect 447416 189382 447468 189388
rect 448428 189440 448480 189446
rect 448428 189382 448480 189388
rect 447048 47592 447100 47598
rect 447048 47534 447100 47540
rect 447140 39364 447192 39370
rect 447140 39306 447192 39312
rect 447152 3482 447180 39306
rect 444392 3454 445432 3482
rect 445404 480 445432 3454
rect 446588 3460 446640 3466
rect 447152 3454 447824 3482
rect 448440 3466 448468 189382
rect 448520 53100 448572 53106
rect 448520 53042 448572 53048
rect 448532 3482 448560 53042
rect 449820 39370 449848 192086
rect 449912 189582 449940 192100
rect 449900 189576 449952 189582
rect 449900 189518 449952 189524
rect 451188 189576 451240 189582
rect 451188 189518 451240 189524
rect 449808 39364 449860 39370
rect 449808 39306 449860 39312
rect 451200 3534 451228 189518
rect 451924 189168 451976 189174
rect 451924 189110 451976 189116
rect 451280 54528 451332 54534
rect 451280 54470 451332 54476
rect 451292 4214 451320 54470
rect 451372 8968 451424 8974
rect 451372 8910 451424 8916
rect 451280 4208 451332 4214
rect 451280 4150 451332 4156
rect 450176 3528 450228 3534
rect 446588 3402 446640 3408
rect 446600 480 446628 3402
rect 447796 480 447824 3454
rect 448428 3460 448480 3466
rect 448532 3454 449020 3482
rect 450176 3470 450228 3476
rect 451188 3528 451240 3534
rect 451384 3482 451412 8910
rect 451936 7614 451964 189110
rect 453316 30326 453344 202671
rect 453408 77246 453436 224023
rect 453500 124166 453528 245375
rect 453592 171086 453620 266727
rect 453684 182170 453712 273799
rect 453946 259720 454002 259729
rect 453946 259655 454002 259664
rect 453960 259486 453988 259655
rect 453948 259480 454000 259486
rect 453948 259422 454000 259428
rect 454696 252550 454724 302330
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 456064 280220 456116 280226
rect 456064 280162 456116 280168
rect 454684 252544 454736 252550
rect 454684 252486 454736 252492
rect 453946 238368 454002 238377
rect 453946 238303 454002 238312
rect 453960 237454 453988 238303
rect 453948 237448 454000 237454
rect 453948 237390 454000 237396
rect 454684 216844 454736 216850
rect 454684 216786 454736 216792
rect 453948 209840 454000 209846
rect 453946 209808 453948 209817
rect 454000 209808 454002 209817
rect 453946 209743 454002 209752
rect 453946 195664 454002 195673
rect 453946 195599 454002 195608
rect 453960 194614 453988 195599
rect 453948 194608 454000 194614
rect 453948 194550 454000 194556
rect 453672 182164 453724 182170
rect 453672 182106 453724 182112
rect 453580 171080 453632 171086
rect 453580 171022 453632 171028
rect 453488 124160 453540 124166
rect 453488 124102 453540 124108
rect 453396 77240 453448 77246
rect 453396 77182 453448 77188
rect 454696 64870 454724 216786
rect 456076 205630 456104 280162
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 471244 259480 471296 259486
rect 471244 259422 471296 259428
rect 469864 237448 469916 237454
rect 469864 237390 469916 237396
rect 456064 205624 456116 205630
rect 456064 205566 456116 205572
rect 456064 189848 456116 189854
rect 456064 189790 456116 189796
rect 454684 64864 454736 64870
rect 454684 64806 454736 64812
rect 454040 64184 454092 64190
rect 454040 64126 454092 64132
rect 453304 30320 453356 30326
rect 453304 30262 453356 30268
rect 451924 7608 451976 7614
rect 451924 7550 451976 7556
rect 452476 4208 452528 4214
rect 452476 4150 452528 4156
rect 451188 3470 451240 3476
rect 448428 3402 448480 3408
rect 448992 480 449020 3454
rect 450188 480 450216 3470
rect 451292 3454 451412 3482
rect 451292 480 451320 3454
rect 452488 480 452516 4150
rect 453672 4140 453724 4146
rect 453672 4082 453724 4088
rect 453684 480 453712 4082
rect 454052 3482 454080 64126
rect 455420 55888 455472 55894
rect 455420 55830 455472 55836
rect 455432 3482 455460 55830
rect 456076 8974 456104 189790
rect 462320 181484 462372 181490
rect 462320 181426 462372 181432
rect 458180 159384 458232 159390
rect 458180 159326 458232 159332
rect 456064 8968 456116 8974
rect 456064 8910 456116 8916
rect 457260 4004 457312 4010
rect 457260 3946 457312 3952
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3946
rect 458192 3482 458220 159326
rect 460940 158024 460992 158030
rect 460940 157966 460992 157972
rect 459652 80708 459704 80714
rect 459652 80650 459704 80656
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 80650
rect 460848 4072 460900 4078
rect 460848 4014 460900 4020
rect 460860 480 460888 4014
rect 460952 3482 460980 157966
rect 462332 3482 462360 181426
rect 466460 140072 466512 140078
rect 466460 140014 466512 140020
rect 465080 28280 465132 28286
rect 465080 28222 465132 28228
rect 464436 3936 464488 3942
rect 464436 3878 464488 3884
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3878
rect 465092 3482 465120 28222
rect 466472 3482 466500 140014
rect 469876 111790 469904 237390
rect 471256 158710 471284 259422
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 479524 250504 479576 250510
rect 479524 250446 479576 250452
rect 472624 230512 472676 230518
rect 472624 230454 472676 230460
rect 471244 158704 471296 158710
rect 471244 158646 471296 158652
rect 469864 111784 469916 111790
rect 469864 111726 469916 111732
rect 469220 111104 469272 111110
rect 469220 111046 469272 111052
rect 467932 26920 467984 26926
rect 467932 26862 467984 26868
rect 467840 3868 467892 3874
rect 467840 3810 467892 3816
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 3210 467880 3810
rect 467944 3398 467972 26862
rect 469232 3482 469260 111046
rect 472636 88330 472664 230454
rect 478144 209840 478196 209846
rect 478144 209782 478196 209788
rect 476120 156664 476172 156670
rect 476120 156606 476172 156612
rect 473360 138712 473412 138718
rect 473360 138654 473412 138660
rect 472624 88324 472676 88330
rect 472624 88266 472676 88272
rect 471980 87644 472032 87650
rect 471980 87586 472032 87592
rect 471520 3800 471572 3806
rect 471520 3742 471572 3748
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 3182 467972 3210
rect 467944 480 467972 3182
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3742
rect 471992 3482 472020 87586
rect 473372 3482 473400 138654
rect 475108 3732 475160 3738
rect 475108 3674 475160 3680
rect 471992 3454 472756 3482
rect 473372 3454 473952 3482
rect 472728 480 472756 3454
rect 473924 480 473952 3454
rect 475120 480 475148 3674
rect 476132 3482 476160 156606
rect 477592 57248 477644 57254
rect 477592 57190 477644 57196
rect 477604 3482 477632 57190
rect 478156 41410 478184 209782
rect 479536 135250 479564 250446
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 483664 194608 483716 194614
rect 483664 194550 483716 194556
rect 480260 137284 480312 137290
rect 480260 137226 480312 137232
rect 479524 135244 479576 135250
rect 479524 135186 479576 135192
rect 478880 134564 478932 134570
rect 478880 134506 478932 134512
rect 478144 41404 478196 41410
rect 478144 41346 478196 41352
rect 478696 3664 478748 3670
rect 478696 3606 478748 3612
rect 476132 3454 476344 3482
rect 476316 480 476344 3454
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 3606
rect 478892 3482 478920 134506
rect 480272 3482 480300 137226
rect 483676 17950 483704 194550
rect 485780 189780 485832 189786
rect 485780 189722 485832 189728
rect 484400 155236 484452 155242
rect 484400 155178 484452 155184
rect 483664 17944 483716 17950
rect 483664 17886 483716 17892
rect 483480 4820 483532 4826
rect 483480 4762 483532 4768
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 478892 3454 479932 3482
rect 480272 3454 481128 3482
rect 479904 480 479932 3454
rect 481100 480 481128 3454
rect 482296 480 482324 3538
rect 483492 480 483520 4762
rect 484412 3482 484440 155178
rect 485792 3602 485820 189722
rect 489920 188352 489972 188358
rect 489920 188294 489972 188300
rect 487160 153876 487212 153882
rect 487160 153818 487212 153824
rect 485872 58676 485924 58682
rect 485872 58618 485924 58624
rect 485780 3596 485832 3602
rect 485780 3538 485832 3544
rect 485884 3482 485912 58618
rect 486976 3596 487028 3602
rect 486976 3538 487028 3544
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 3454 485912 3482
rect 485792 480 485820 3454
rect 486988 480 487016 3538
rect 487172 3482 487200 153818
rect 488540 60036 488592 60042
rect 488540 59978 488592 59984
rect 488552 3482 488580 59978
rect 489932 3482 489960 188294
rect 494060 186992 494112 186998
rect 494060 186934 494112 186940
rect 492680 61396 492732 61402
rect 492680 61338 492732 61344
rect 491300 32428 491352 32434
rect 491300 32370 491352 32376
rect 491312 3482 491340 32370
rect 492692 3482 492720 61338
rect 494072 3482 494100 186934
rect 500960 185632 501012 185638
rect 500960 185574 501012 185580
rect 498200 152516 498252 152522
rect 498200 152458 498252 152464
rect 495440 135924 495492 135930
rect 495440 135866 495492 135872
rect 494152 15904 494204 15910
rect 494152 15846 494204 15852
rect 494164 3602 494192 15846
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 489932 3454 490604 3482
rect 491312 3454 491800 3482
rect 492692 3454 492996 3482
rect 494072 3454 494192 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 490576 480 490604 3454
rect 491772 480 491800 3454
rect 492968 480 492996 3454
rect 494164 480 494192 3454
rect 495360 480 495388 3538
rect 495452 3482 495480 135866
rect 497740 6180 497792 6186
rect 497740 6122 497792 6128
rect 495452 3454 496584 3482
rect 496556 480 496584 3454
rect 497752 480 497780 6122
rect 498212 3482 498240 152458
rect 499580 62824 499632 62830
rect 499580 62766 499632 62772
rect 499592 3482 499620 62766
rect 500972 3482 501000 185574
rect 503720 184204 503772 184210
rect 503720 184146 503772 184152
rect 502340 108316 502392 108322
rect 502340 108258 502392 108264
rect 498212 3454 498976 3482
rect 499592 3454 500172 3482
rect 500972 3454 501276 3482
rect 498948 480 498976 3454
rect 500144 480 500172 3454
rect 501248 480 501276 3454
rect 502352 2786 502380 108258
rect 502432 10328 502484 10334
rect 502432 10270 502484 10276
rect 502340 2780 502392 2786
rect 502340 2722 502392 2728
rect 502444 480 502472 10270
rect 503732 3482 503760 184146
rect 507860 182844 507912 182850
rect 507860 182786 507912 182792
rect 505100 151088 505152 151094
rect 505100 151030 505152 151036
rect 505112 3482 505140 151030
rect 506480 82136 506532 82142
rect 506480 82078 506532 82084
rect 506492 3482 506520 82078
rect 507872 3482 507900 182786
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 512000 180124 512052 180130
rect 512000 180066 512052 180072
rect 510620 79348 510672 79354
rect 510620 79290 510672 79296
rect 509240 18624 509292 18630
rect 509240 18566 509292 18572
rect 509252 3482 509280 18566
rect 510632 3482 510660 79290
rect 503732 3454 504864 3482
rect 505112 3454 506060 3482
rect 506492 3454 507256 3482
rect 507872 3454 508452 3482
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 503628 2780 503680 2786
rect 503628 2722 503680 2728
rect 503640 480 503668 2722
rect 504836 480 504864 3454
rect 506032 480 506060 3454
rect 507228 480 507256 3454
rect 508424 480 508452 3454
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 480 512040 180066
rect 518900 178696 518952 178702
rect 518900 178638 518952 178644
rect 516140 149728 516192 149734
rect 516140 149670 516192 149676
rect 513380 133204 513432 133210
rect 513380 133146 513432 133152
rect 512092 35216 512144 35222
rect 512092 35158 512144 35164
rect 512104 3482 512132 35158
rect 513392 3482 513420 133146
rect 514760 11756 514812 11762
rect 514760 11698 514812 11704
rect 514772 3482 514800 11698
rect 516152 3482 516180 149670
rect 517520 65544 517572 65550
rect 517520 65486 517572 65492
rect 517532 3482 517560 65486
rect 518912 3482 518940 178638
rect 521660 177336 521712 177342
rect 521660 177278 521712 177284
rect 520280 68332 520332 68338
rect 520280 68274 520332 68280
rect 520292 3602 520320 68274
rect 520372 31068 520424 31074
rect 520372 31010 520424 31016
rect 520280 3596 520332 3602
rect 520280 3538 520332 3544
rect 512104 3454 513236 3482
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513208 480 513236 3454
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520384 1578 520412 31010
rect 521476 3596 521528 3602
rect 521476 3538 521528 3544
rect 520292 1550 520412 1578
rect 520292 480 520320 1550
rect 521488 480 521516 3538
rect 521672 3482 521700 177278
rect 525800 175976 525852 175982
rect 525800 175918 525852 175924
rect 524420 69692 524472 69698
rect 524420 69634 524472 69640
rect 523040 33788 523092 33794
rect 523040 33730 523092 33736
rect 523052 3482 523080 33730
rect 524432 3482 524460 69634
rect 525812 3482 525840 175918
rect 528560 174548 528612 174554
rect 528560 174490 528612 174496
rect 527180 21412 527232 21418
rect 527180 21354 527232 21360
rect 527192 3482 527220 21354
rect 528572 3602 528600 174490
rect 536840 173188 536892 173194
rect 536840 173130 536892 173136
rect 529940 148368 529992 148374
rect 529940 148310 529992 148316
rect 528652 66904 528704 66910
rect 528652 66846 528704 66852
rect 528560 3596 528612 3602
rect 528560 3538 528612 3544
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 525812 3454 526300 3482
rect 527192 3454 527496 3482
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 3454
rect 527468 480 527496 3454
rect 528664 480 528692 66846
rect 529848 3596 529900 3602
rect 529848 3538 529900 3544
rect 529860 480 529888 3538
rect 529952 3482 529980 148310
rect 534080 146940 534132 146946
rect 534080 146882 534132 146888
rect 531320 131776 531372 131782
rect 531320 131718 531372 131724
rect 531332 3482 531360 131718
rect 532700 13116 532752 13122
rect 532700 13058 532752 13064
rect 532712 3482 532740 13058
rect 534092 3482 534120 146882
rect 535460 77988 535512 77994
rect 535460 77930 535512 77936
rect 535472 3482 535500 77930
rect 536852 3482 536880 173130
rect 539600 171828 539652 171834
rect 539600 171770 539652 171776
rect 538220 72480 538272 72486
rect 538220 72422 538272 72428
rect 536932 22772 536984 22778
rect 536932 22714 536984 22720
rect 536944 3602 536972 22714
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 538128 3596 538180 3602
rect 538128 3538 538180 3544
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 3538
rect 538232 3482 538260 72422
rect 539612 3482 539640 171770
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 543740 169040 543792 169046
rect 543740 168982 543792 168988
rect 542360 75200 542412 75206
rect 542360 75142 542412 75148
rect 540980 37936 541032 37942
rect 540980 37878 541032 37884
rect 540992 3482 541020 37878
rect 542372 3482 542400 75142
rect 543752 3482 543780 168982
rect 546500 167680 546552 167686
rect 546500 167622 546552 167628
rect 545120 42084 545172 42090
rect 545120 42026 545172 42032
rect 545132 3482 545160 42026
rect 546512 3602 546540 167622
rect 554780 166320 554832 166326
rect 554780 166262 554832 166268
rect 547880 145580 547932 145586
rect 547880 145522 547932 145528
rect 546592 44872 546644 44878
rect 546592 44814 546644 44820
rect 546500 3596 546552 3602
rect 546500 3538 546552 3544
rect 546604 3482 546632 44814
rect 547696 3596 547748 3602
rect 547696 3538 547748 3544
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 3454 546632 3482
rect 546512 480 546540 3454
rect 547708 480 547736 3538
rect 547892 3482 547920 145522
rect 552020 144220 552072 144226
rect 552020 144162 552072 144168
rect 549260 49020 549312 49026
rect 549260 48962 549312 48968
rect 549272 3482 549300 48962
rect 550640 19984 550692 19990
rect 550640 19926 550692 19932
rect 550652 3482 550680 19926
rect 552032 3482 552060 144162
rect 553400 83496 553452 83502
rect 553400 83438 553452 83444
rect 553412 3482 553440 83438
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 166262
rect 557540 164892 557592 164898
rect 557540 164834 557592 164840
rect 556160 130416 556212 130422
rect 556160 130358 556212 130364
rect 554872 24132 554924 24138
rect 554872 24074 554924 24080
rect 554884 3482 554912 24074
rect 556172 3482 556200 130358
rect 557552 3482 557580 164834
rect 561680 163532 561732 163538
rect 561680 163474 561732 163480
rect 560300 71052 560352 71058
rect 560300 70994 560352 71000
rect 558920 43444 558972 43450
rect 558920 43386 558972 43392
rect 558932 3482 558960 43386
rect 560312 3482 560340 70994
rect 561692 3482 561720 163474
rect 564440 162172 564492 162178
rect 564440 162114 564492 162120
rect 563060 86284 563112 86290
rect 563060 86226 563112 86232
rect 554884 3454 556016 3482
rect 556172 3454 557212 3482
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 560312 3454 560800 3482
rect 561692 3454 561996 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3454
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3454
rect 561968 480 561996 3454
rect 563072 2786 563100 86226
rect 563152 14476 563204 14482
rect 563152 14418 563204 14424
rect 563060 2780 563112 2786
rect 563060 2722 563112 2728
rect 563164 480 563192 14418
rect 564452 3482 564480 162114
rect 571340 160744 571392 160750
rect 571340 160686 571392 160692
rect 565820 142860 565872 142866
rect 565820 142802 565872 142808
rect 565832 3482 565860 142802
rect 569960 141432 570012 141438
rect 569960 141374 570012 141380
rect 567200 46232 567252 46238
rect 567200 46174 567252 46180
rect 567212 3482 567240 46174
rect 568580 25560 568632 25566
rect 568580 25502 568632 25508
rect 568592 3482 568620 25502
rect 569972 3482 570000 141374
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 567212 3454 567884 3482
rect 568592 3454 569080 3482
rect 569972 3454 570276 3482
rect 564348 2780 564400 2786
rect 564348 2722 564400 2728
rect 564360 480 564388 2722
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3454
rect 569052 480 569080 3454
rect 570248 480 570276 3454
rect 571352 2786 571380 160686
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 573364 73840 573416 73846
rect 573364 73782 573416 73788
rect 571432 50380 571484 50386
rect 571432 50322 571484 50328
rect 571340 2780 571392 2786
rect 571340 2722 571392 2728
rect 571444 480 571472 50322
rect 572720 36576 572772 36582
rect 572720 36518 572772 36524
rect 572732 3346 572760 36518
rect 573376 3602 573404 73782
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 574744 47592 574796 47598
rect 574744 47534 574796 47540
rect 574756 4146 574784 47534
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 574836 39364 574888 39370
rect 574836 39306 574888 39312
rect 574744 4140 574796 4146
rect 574744 4082 574796 4088
rect 574848 3670 574876 39306
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 579804 8968 579856 8974
rect 579804 8910 579856 8916
rect 576216 7608 576268 7614
rect 576216 7550 576268 7556
rect 574836 3664 574888 3670
rect 574836 3606 574888 3612
rect 573364 3596 573416 3602
rect 573364 3538 573416 3544
rect 575020 3596 575072 3602
rect 575020 3538 575072 3544
rect 572732 3318 573864 3346
rect 572628 2780 572680 2786
rect 572628 2722 572680 2728
rect 572640 480 572668 2722
rect 573836 480 573864 3318
rect 575032 480 575060 3538
rect 576228 480 576256 7550
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 579816 480 579844 8910
rect 581000 3664 581052 3670
rect 581000 3606 581052 3612
rect 581012 480 581040 3606
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 582208 480 582236 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 4066 567316 4122 567352
rect 4066 567296 4068 567316
rect 4068 567296 4120 567316
rect 4120 567296 4122 567316
rect 3422 553016 3478 553072
rect 2870 509904 2926 509960
rect 3330 481072 3386 481128
rect 7930 540912 7986 540968
rect 8206 540912 8262 540968
rect 3698 538600 3754 538656
rect 8114 531256 8170 531312
rect 8298 531256 8354 531312
rect 3514 495488 3570 495544
rect 3146 452376 3202 452432
rect 3422 437960 3478 438016
rect 72974 608504 73030 608560
rect 73158 608504 73214 608560
rect 128358 508544 128414 508600
rect 128358 500928 128414 500984
rect 128358 493312 128414 493368
rect 128358 485732 128360 485752
rect 128360 485732 128412 485752
rect 128412 485732 128414 485752
rect 128358 485696 128414 485732
rect 128358 478080 128414 478136
rect 154210 540912 154266 540968
rect 154486 540912 154542 540968
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 284206 540912 284262 540968
rect 284390 540912 284446 540968
rect 284114 531256 284170 531312
rect 284298 531256 284354 531312
rect 347870 560224 347926 560280
rect 348054 560224 348110 560280
rect 364430 560224 364486 560280
rect 364614 560224 364670 560280
rect 347870 540912 347926 540968
rect 348054 540912 348110 540968
rect 364430 540912 364486 540968
rect 364614 540912 364670 540968
rect 453210 508816 453266 508872
rect 453394 501744 453450 501800
rect 453946 494536 454002 494592
rect 453762 487464 453818 487520
rect 453762 480392 453818 480448
rect 453946 473184 454002 473240
rect 129002 470464 129058 470520
rect 452750 466112 452806 466168
rect 128358 462848 128414 462904
rect 453394 459040 453450 459096
rect 128358 455232 128414 455288
rect 453946 451832 454002 451888
rect 3514 423680 3570 423736
rect 128358 447616 128414 447672
rect 453670 444760 453726 444816
rect 128358 440000 128414 440056
rect 128358 432248 128414 432304
rect 128358 424632 128414 424688
rect 128358 417016 128414 417072
rect 128358 409400 128414 409456
rect 452842 402056 452898 402112
rect 128358 401784 128414 401840
rect 3422 394984 3478 395040
rect 128358 394168 128414 394224
rect 453762 437688 453818 437744
rect 453946 430516 453948 430536
rect 453948 430516 454000 430536
rect 454000 430516 454002 430536
rect 453946 430480 454002 430516
rect 453946 423408 454002 423464
rect 453946 416372 453948 416392
rect 453948 416372 454000 416392
rect 454000 416372 454002 416392
rect 453946 416336 454002 416372
rect 453394 409128 453450 409184
rect 477590 560224 477646 560280
rect 477774 560224 477830 560280
rect 477590 540912 477646 540968
rect 477774 540912 477830 540968
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 494150 560224 494206 560280
rect 494334 560224 494390 560280
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 580170 697992 580226 698048
rect 580262 686296 580318 686352
rect 542358 683168 542414 683224
rect 542726 683168 542782 683224
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 579894 592456 579950 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 579894 545536 579950 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580354 639376 580410 639432
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580262 451696 580318 451752
rect 579894 439864 579950 439920
rect 580170 416472 580226 416528
rect 453762 394848 453818 394904
rect 453302 387776 453358 387832
rect 129002 386552 129058 386608
rect 453946 380704 454002 380760
rect 3238 380568 3294 380624
rect 129002 378936 129058 378992
rect 453394 373496 453450 373552
rect 129278 371320 129334 371376
rect 3146 366152 3202 366208
rect 129002 363704 129058 363760
rect 128358 348336 128414 348392
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 3330 308760 3386 308816
rect 128358 333104 128414 333160
rect 3514 294344 3570 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3146 265648 3202 265704
rect 3422 251232 3478 251288
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 3422 208120 3478 208176
rect 3146 193840 3202 193896
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 128358 325488 128414 325544
rect 129186 356088 129242 356144
rect 129094 340720 129150 340776
rect 129002 317872 129058 317928
rect 128358 310256 128414 310312
rect 3514 78920 3570 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 128358 302640 128414 302696
rect 128358 287408 128414 287464
rect 128358 264424 128414 264480
rect 128358 256808 128414 256864
rect 128358 241576 128414 241632
rect 580354 404776 580410 404832
rect 580170 392944 580226 393000
rect 580262 369552 580318 369608
rect 452658 366424 452714 366480
rect 453946 359352 454002 359408
rect 580262 357856 580318 357912
rect 453762 352144 453818 352200
rect 580170 346024 580226 346080
rect 453946 345072 454002 345128
rect 453486 338000 453542 338056
rect 453394 330792 453450 330848
rect 453302 323720 453358 323776
rect 452934 302388 452990 302424
rect 452934 302368 452936 302388
rect 452936 302368 452988 302388
rect 452988 302368 452990 302388
rect 580170 322632 580226 322688
rect 453578 316648 453634 316704
rect 453486 309440 453542 309496
rect 453394 295160 453450 295216
rect 129370 295024 129426 295080
rect 129094 279792 129150 279848
rect 129278 272040 129334 272096
rect 129186 249192 129242 249248
rect 128358 233960 128414 234016
rect 129094 226344 129150 226400
rect 128358 218728 128414 218784
rect 128358 211148 128360 211168
rect 128360 211148 128412 211168
rect 128412 211148 128414 211168
rect 128358 211112 128414 211148
rect 129002 203496 129058 203552
rect 128634 195880 128690 195936
rect 453302 288088 453358 288144
rect 453026 281016 453082 281072
rect 452842 252456 452898 252512
rect 453118 231104 453174 231160
rect 580170 310800 580226 310856
rect 453670 273808 453726 273864
rect 453578 266736 453634 266792
rect 453486 245384 453542 245440
rect 453394 224032 453450 224088
rect 452934 216960 452990 217016
rect 453302 202680 453358 202736
rect 3422 7112 3478 7168
rect 135350 183504 135406 183560
rect 135534 183504 135590 183560
rect 135350 154536 135406 154592
rect 135626 154536 135682 154592
rect 135350 135224 135406 135280
rect 135626 135224 135682 135280
rect 135350 115912 135406 115968
rect 135626 115912 135682 115968
rect 135350 96600 135406 96656
rect 135626 96600 135682 96656
rect 453946 259664 454002 259720
rect 579802 299104 579858 299160
rect 453946 238312 454002 238368
rect 453946 209788 453948 209808
rect 453948 209788 454000 209808
rect 454000 209788 454002 209808
rect 453946 209752 454002 209788
rect 453946 195608 454002 195664
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 542353 683226 542419 683229
rect 542721 683226 542787 683229
rect 542353 683224 542787 683226
rect 542353 683168 542358 683224
rect 542414 683168 542726 683224
rect 542782 683168 542787 683224
rect 542353 683166 542787 683168
rect 542353 683163 542419 683166
rect 542721 683163 542787 683166
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 72969 608562 73035 608565
rect 73153 608562 73219 608565
rect 72969 608560 73219 608562
rect 72969 608504 72974 608560
rect 73030 608504 73158 608560
rect 73214 608504 73219 608560
rect 72969 608502 73219 608504
rect 72969 608499 73035 608502
rect 73153 608499 73219 608502
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 579889 592514 579955 592517
rect 583520 592514 584960 592604
rect 579889 592512 584960 592514
rect 579889 592456 579894 592512
rect 579950 592456 584960 592512
rect 579889 592454 584960 592456
rect 579889 592451 579955 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 347865 560282 347931 560285
rect 348049 560282 348115 560285
rect 347865 560280 348115 560282
rect 347865 560224 347870 560280
rect 347926 560224 348054 560280
rect 348110 560224 348115 560280
rect 347865 560222 348115 560224
rect 347865 560219 347931 560222
rect 348049 560219 348115 560222
rect 364425 560282 364491 560285
rect 364609 560282 364675 560285
rect 364425 560280 364675 560282
rect 364425 560224 364430 560280
rect 364486 560224 364614 560280
rect 364670 560224 364675 560280
rect 364425 560222 364675 560224
rect 364425 560219 364491 560222
rect 364609 560219 364675 560222
rect 477585 560282 477651 560285
rect 477769 560282 477835 560285
rect 477585 560280 477835 560282
rect 477585 560224 477590 560280
rect 477646 560224 477774 560280
rect 477830 560224 477835 560280
rect 477585 560222 477835 560224
rect 477585 560219 477651 560222
rect 477769 560219 477835 560222
rect 494145 560282 494211 560285
rect 494329 560282 494395 560285
rect 494145 560280 494395 560282
rect 494145 560224 494150 560280
rect 494206 560224 494334 560280
rect 494390 560224 494395 560280
rect 494145 560222 494395 560224
rect 494145 560219 494211 560222
rect 494329 560219 494395 560222
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 579889 545594 579955 545597
rect 583520 545594 584960 545684
rect 579889 545592 584960 545594
rect 579889 545536 579894 545592
rect 579950 545536 584960 545592
rect 579889 545534 584960 545536
rect 579889 545531 579955 545534
rect 583520 545444 584960 545534
rect 7925 540970 7991 540973
rect 8201 540970 8267 540973
rect 7925 540968 8267 540970
rect 7925 540912 7930 540968
rect 7986 540912 8206 540968
rect 8262 540912 8267 540968
rect 7925 540910 8267 540912
rect 7925 540907 7991 540910
rect 8201 540907 8267 540910
rect 154205 540970 154271 540973
rect 154481 540970 154547 540973
rect 154205 540968 154547 540970
rect 154205 540912 154210 540968
rect 154266 540912 154486 540968
rect 154542 540912 154547 540968
rect 154205 540910 154547 540912
rect 154205 540907 154271 540910
rect 154481 540907 154547 540910
rect 284201 540970 284267 540973
rect 284385 540970 284451 540973
rect 284201 540968 284451 540970
rect 284201 540912 284206 540968
rect 284262 540912 284390 540968
rect 284446 540912 284451 540968
rect 284201 540910 284451 540912
rect 284201 540907 284267 540910
rect 284385 540907 284451 540910
rect 347865 540970 347931 540973
rect 348049 540970 348115 540973
rect 347865 540968 348115 540970
rect 347865 540912 347870 540968
rect 347926 540912 348054 540968
rect 348110 540912 348115 540968
rect 347865 540910 348115 540912
rect 347865 540907 347931 540910
rect 348049 540907 348115 540910
rect 364425 540970 364491 540973
rect 364609 540970 364675 540973
rect 364425 540968 364675 540970
rect 364425 540912 364430 540968
rect 364486 540912 364614 540968
rect 364670 540912 364675 540968
rect 364425 540910 364675 540912
rect 364425 540907 364491 540910
rect 364609 540907 364675 540910
rect 477585 540970 477651 540973
rect 477769 540970 477835 540973
rect 477585 540968 477835 540970
rect 477585 540912 477590 540968
rect 477646 540912 477774 540968
rect 477830 540912 477835 540968
rect 477585 540910 477835 540912
rect 477585 540907 477651 540910
rect 477769 540907 477835 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -960 538658 480 538748
rect 3693 538658 3759 538661
rect -960 538656 3759 538658
rect -960 538600 3698 538656
rect 3754 538600 3759 538656
rect -960 538598 3759 538600
rect -960 538508 480 538598
rect 3693 538595 3759 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 8109 531314 8175 531317
rect 8293 531314 8359 531317
rect 8109 531312 8359 531314
rect 8109 531256 8114 531312
rect 8170 531256 8298 531312
rect 8354 531256 8359 531312
rect 8109 531254 8359 531256
rect 8109 531251 8175 531254
rect 8293 531251 8359 531254
rect 284109 531314 284175 531317
rect 284293 531314 284359 531317
rect 284109 531312 284359 531314
rect 284109 531256 284114 531312
rect 284170 531256 284298 531312
rect 284354 531256 284359 531312
rect 284109 531254 284359 531256
rect 284109 531251 284175 531254
rect 284293 531251 284359 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 2865 509962 2931 509965
rect -960 509960 2931 509962
rect -960 509904 2870 509960
rect 2926 509904 2931 509960
rect -960 509902 2931 509904
rect -960 509812 480 509902
rect 2865 509899 2931 509902
rect 453205 508874 453271 508877
rect 450156 508872 453271 508874
rect 450156 508816 453210 508872
rect 453266 508816 453271 508872
rect 450156 508814 453271 508816
rect 453205 508811 453271 508814
rect 128353 508602 128419 508605
rect 128353 508600 132020 508602
rect 128353 508544 128358 508600
rect 128414 508544 132020 508600
rect 128353 508542 132020 508544
rect 128353 508539 128419 508542
rect 453389 501802 453455 501805
rect 450156 501800 453455 501802
rect 450156 501744 453394 501800
rect 453450 501744 453455 501800
rect 450156 501742 453455 501744
rect 453389 501739 453455 501742
rect 128353 500986 128419 500989
rect 128353 500984 132020 500986
rect 128353 500928 128358 500984
rect 128414 500928 132020 500984
rect 128353 500926 132020 500928
rect 128353 500923 128419 500926
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 453941 494594 454007 494597
rect 450156 494592 454007 494594
rect 450156 494536 453946 494592
rect 454002 494536 454007 494592
rect 450156 494534 454007 494536
rect 453941 494531 454007 494534
rect 128353 493370 128419 493373
rect 128353 493368 132020 493370
rect 128353 493312 128358 493368
rect 128414 493312 132020 493368
rect 128353 493310 132020 493312
rect 128353 493307 128419 493310
rect 453757 487522 453823 487525
rect 450156 487520 453823 487522
rect 450156 487464 453762 487520
rect 453818 487464 453823 487520
rect 450156 487462 453823 487464
rect 453757 487459 453823 487462
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 128353 485754 128419 485757
rect 128353 485752 132020 485754
rect 128353 485696 128358 485752
rect 128414 485696 132020 485752
rect 128353 485694 132020 485696
rect 128353 485691 128419 485694
rect -960 481130 480 481220
rect 3325 481130 3391 481133
rect -960 481128 3391 481130
rect -960 481072 3330 481128
rect 3386 481072 3391 481128
rect -960 481070 3391 481072
rect -960 480980 480 481070
rect 3325 481067 3391 481070
rect 453757 480450 453823 480453
rect 450156 480448 453823 480450
rect 450156 480392 453762 480448
rect 453818 480392 453823 480448
rect 450156 480390 453823 480392
rect 453757 480387 453823 480390
rect 128353 478138 128419 478141
rect 128353 478136 132020 478138
rect 128353 478080 128358 478136
rect 128414 478080 132020 478136
rect 128353 478078 132020 478080
rect 128353 478075 128419 478078
rect 583520 474996 584960 475236
rect 453941 473242 454007 473245
rect 450156 473240 454007 473242
rect 450156 473184 453946 473240
rect 454002 473184 454007 473240
rect 450156 473182 454007 473184
rect 453941 473179 454007 473182
rect 128997 470522 129063 470525
rect 128997 470520 132020 470522
rect 128997 470464 129002 470520
rect 129058 470464 132020 470520
rect 128997 470462 132020 470464
rect 128997 470459 129063 470462
rect -960 466700 480 466940
rect 452745 466170 452811 466173
rect 450156 466168 452811 466170
rect 450156 466112 452750 466168
rect 452806 466112 452811 466168
rect 450156 466110 452811 466112
rect 452745 466107 452811 466110
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 128353 462906 128419 462909
rect 128353 462904 132020 462906
rect 128353 462848 128358 462904
rect 128414 462848 132020 462904
rect 128353 462846 132020 462848
rect 128353 462843 128419 462846
rect 453389 459098 453455 459101
rect 450156 459096 453455 459098
rect 450156 459040 453394 459096
rect 453450 459040 453455 459096
rect 450156 459038 453455 459040
rect 453389 459035 453455 459038
rect 128353 455290 128419 455293
rect 128353 455288 132020 455290
rect 128353 455232 128358 455288
rect 128414 455232 132020 455288
rect 128353 455230 132020 455232
rect 128353 455227 128419 455230
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 453941 451890 454007 451893
rect 450156 451888 454007 451890
rect 450156 451832 453946 451888
rect 454002 451832 454007 451888
rect 450156 451830 454007 451832
rect 453941 451827 454007 451830
rect 580257 451754 580323 451757
rect 583520 451754 584960 451844
rect 580257 451752 584960 451754
rect 580257 451696 580262 451752
rect 580318 451696 584960 451752
rect 580257 451694 584960 451696
rect 580257 451691 580323 451694
rect 583520 451604 584960 451694
rect 128353 447674 128419 447677
rect 128353 447672 132020 447674
rect 128353 447616 128358 447672
rect 128414 447616 132020 447672
rect 128353 447614 132020 447616
rect 128353 447611 128419 447614
rect 453665 444818 453731 444821
rect 450156 444816 453731 444818
rect 450156 444760 453670 444816
rect 453726 444760 453731 444816
rect 450156 444758 453731 444760
rect 453665 444755 453731 444758
rect 128353 440058 128419 440061
rect 128353 440056 132020 440058
rect 128353 440000 128358 440056
rect 128414 440000 132020 440056
rect 128353 439998 132020 440000
rect 128353 439995 128419 439998
rect 579889 439922 579955 439925
rect 583520 439922 584960 440012
rect 579889 439920 584960 439922
rect 579889 439864 579894 439920
rect 579950 439864 584960 439920
rect 579889 439862 584960 439864
rect 579889 439859 579955 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3417 438018 3483 438021
rect -960 438016 3483 438018
rect -960 437960 3422 438016
rect 3478 437960 3483 438016
rect -960 437958 3483 437960
rect -960 437868 480 437958
rect 3417 437955 3483 437958
rect 453757 437746 453823 437749
rect 450156 437744 453823 437746
rect 450156 437688 453762 437744
rect 453818 437688 453823 437744
rect 450156 437686 453823 437688
rect 453757 437683 453823 437686
rect 128353 432306 128419 432309
rect 128353 432304 132020 432306
rect 128353 432248 128358 432304
rect 128414 432248 132020 432304
rect 128353 432246 132020 432248
rect 128353 432243 128419 432246
rect 453941 430538 454007 430541
rect 450156 430536 454007 430538
rect 450156 430480 453946 430536
rect 454002 430480 454007 430536
rect 450156 430478 454007 430480
rect 453941 430475 454007 430478
rect 583520 428076 584960 428316
rect 128353 424690 128419 424693
rect 128353 424688 132020 424690
rect 128353 424632 128358 424688
rect 128414 424632 132020 424688
rect 128353 424630 132020 424632
rect 128353 424627 128419 424630
rect -960 423738 480 423828
rect 3509 423738 3575 423741
rect -960 423736 3575 423738
rect -960 423680 3514 423736
rect 3570 423680 3575 423736
rect -960 423678 3575 423680
rect -960 423588 480 423678
rect 3509 423675 3575 423678
rect 453941 423466 454007 423469
rect 450156 423464 454007 423466
rect 450156 423408 453946 423464
rect 454002 423408 454007 423464
rect 450156 423406 454007 423408
rect 453941 423403 454007 423406
rect 128353 417074 128419 417077
rect 128353 417072 132020 417074
rect 128353 417016 128358 417072
rect 128414 417016 132020 417072
rect 128353 417014 132020 417016
rect 128353 417011 128419 417014
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 453941 416394 454007 416397
rect 450156 416392 454007 416394
rect 450156 416336 453946 416392
rect 454002 416336 454007 416392
rect 583520 416380 584960 416470
rect 450156 416334 454007 416336
rect 453941 416331 454007 416334
rect 128353 409458 128419 409461
rect 128353 409456 132020 409458
rect -960 409172 480 409412
rect 128353 409400 128358 409456
rect 128414 409400 132020 409456
rect 128353 409398 132020 409400
rect 128353 409395 128419 409398
rect 453389 409186 453455 409189
rect 450156 409184 453455 409186
rect 450156 409128 453394 409184
rect 453450 409128 453455 409184
rect 450156 409126 453455 409128
rect 453389 409123 453455 409126
rect 580349 404834 580415 404837
rect 583520 404834 584960 404924
rect 580349 404832 584960 404834
rect 580349 404776 580354 404832
rect 580410 404776 584960 404832
rect 580349 404774 584960 404776
rect 580349 404771 580415 404774
rect 583520 404684 584960 404774
rect 452837 402114 452903 402117
rect 450156 402112 452903 402114
rect 450156 402056 452842 402112
rect 452898 402056 452903 402112
rect 450156 402054 452903 402056
rect 452837 402051 452903 402054
rect 128353 401842 128419 401845
rect 128353 401840 132020 401842
rect 128353 401784 128358 401840
rect 128414 401784 132020 401840
rect 128353 401782 132020 401784
rect 128353 401779 128419 401782
rect -960 395042 480 395132
rect 3417 395042 3483 395045
rect -960 395040 3483 395042
rect -960 394984 3422 395040
rect 3478 394984 3483 395040
rect -960 394982 3483 394984
rect -960 394892 480 394982
rect 3417 394979 3483 394982
rect 453757 394906 453823 394909
rect 450156 394904 453823 394906
rect 450156 394848 453762 394904
rect 453818 394848 453823 394904
rect 450156 394846 453823 394848
rect 453757 394843 453823 394846
rect 128353 394226 128419 394229
rect 128353 394224 132020 394226
rect 128353 394168 128358 394224
rect 128414 394168 132020 394224
rect 128353 394166 132020 394168
rect 128353 394163 128419 394166
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 453297 387834 453363 387837
rect 450156 387832 453363 387834
rect 450156 387776 453302 387832
rect 453358 387776 453363 387832
rect 450156 387774 453363 387776
rect 453297 387771 453363 387774
rect 128997 386610 129063 386613
rect 128997 386608 132020 386610
rect 128997 386552 129002 386608
rect 129058 386552 132020 386608
rect 128997 386550 132020 386552
rect 128997 386547 129063 386550
rect 583520 381156 584960 381396
rect 453941 380762 454007 380765
rect 450156 380760 454007 380762
rect -960 380626 480 380716
rect 450156 380704 453946 380760
rect 454002 380704 454007 380760
rect 450156 380702 454007 380704
rect 453941 380699 454007 380702
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 128997 378994 129063 378997
rect 128997 378992 132020 378994
rect 128997 378936 129002 378992
rect 129058 378936 132020 378992
rect 128997 378934 132020 378936
rect 128997 378931 129063 378934
rect 453389 373554 453455 373557
rect 450156 373552 453455 373554
rect 450156 373496 453394 373552
rect 453450 373496 453455 373552
rect 450156 373494 453455 373496
rect 453389 373491 453455 373494
rect 129273 371378 129339 371381
rect 129273 371376 132020 371378
rect 129273 371320 129278 371376
rect 129334 371320 132020 371376
rect 129273 371318 132020 371320
rect 129273 371315 129339 371318
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 583520 369460 584960 369550
rect 452653 366482 452719 366485
rect 450156 366480 452719 366482
rect 450156 366424 452658 366480
rect 452714 366424 452719 366480
rect 450156 366422 452719 366424
rect 452653 366419 452719 366422
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 128997 363762 129063 363765
rect 128997 363760 132020 363762
rect 128997 363704 129002 363760
rect 129058 363704 132020 363760
rect 128997 363702 132020 363704
rect 128997 363699 129063 363702
rect 453941 359410 454007 359413
rect 450156 359408 454007 359410
rect 450156 359352 453946 359408
rect 454002 359352 454007 359408
rect 450156 359350 454007 359352
rect 453941 359347 454007 359350
rect 580257 357914 580323 357917
rect 583520 357914 584960 358004
rect 580257 357912 584960 357914
rect 580257 357856 580262 357912
rect 580318 357856 584960 357912
rect 580257 357854 584960 357856
rect 580257 357851 580323 357854
rect 583520 357764 584960 357854
rect 129181 356146 129247 356149
rect 129181 356144 132020 356146
rect 129181 356088 129186 356144
rect 129242 356088 132020 356144
rect 129181 356086 132020 356088
rect 129181 356083 129247 356086
rect 453757 352202 453823 352205
rect 450156 352200 453823 352202
rect 450156 352144 453762 352200
rect 453818 352144 453823 352200
rect 450156 352142 453823 352144
rect 453757 352139 453823 352142
rect -960 351780 480 352020
rect 128353 348394 128419 348397
rect 128353 348392 132020 348394
rect 128353 348336 128358 348392
rect 128414 348336 132020 348392
rect 128353 348334 132020 348336
rect 128353 348331 128419 348334
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 453941 345130 454007 345133
rect 450156 345128 454007 345130
rect 450156 345072 453946 345128
rect 454002 345072 454007 345128
rect 450156 345070 454007 345072
rect 453941 345067 454007 345070
rect 129089 340778 129155 340781
rect 129089 340776 132020 340778
rect 129089 340720 129094 340776
rect 129150 340720 132020 340776
rect 129089 340718 132020 340720
rect 129089 340715 129155 340718
rect 453481 338058 453547 338061
rect 450156 338056 453547 338058
rect 450156 338000 453486 338056
rect 453542 338000 453547 338056
rect 450156 337998 453547 338000
rect 453481 337995 453547 337998
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 583520 334236 584960 334476
rect 128353 333162 128419 333165
rect 128353 333160 132020 333162
rect 128353 333104 128358 333160
rect 128414 333104 132020 333160
rect 128353 333102 132020 333104
rect 128353 333099 128419 333102
rect 453389 330850 453455 330853
rect 450156 330848 453455 330850
rect 450156 330792 453394 330848
rect 453450 330792 453455 330848
rect 450156 330790 453455 330792
rect 453389 330787 453455 330790
rect 128353 325546 128419 325549
rect 128353 325544 132020 325546
rect 128353 325488 128358 325544
rect 128414 325488 132020 325544
rect 128353 325486 132020 325488
rect 128353 325483 128419 325486
rect 453297 323778 453363 323781
rect 450156 323776 453363 323778
rect 450156 323720 453302 323776
rect 453358 323720 453363 323776
rect 450156 323718 453363 323720
rect 453297 323715 453363 323718
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 128997 317930 129063 317933
rect 128997 317928 132020 317930
rect 128997 317872 129002 317928
rect 129058 317872 132020 317928
rect 128997 317870 132020 317872
rect 128997 317867 129063 317870
rect 453573 316706 453639 316709
rect 450156 316704 453639 316706
rect 450156 316648 453578 316704
rect 453634 316648 453639 316704
rect 450156 316646 453639 316648
rect 453573 316643 453639 316646
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 128353 310314 128419 310317
rect 128353 310312 132020 310314
rect 128353 310256 128358 310312
rect 128414 310256 132020 310312
rect 128353 310254 132020 310256
rect 128353 310251 128419 310254
rect 453481 309498 453547 309501
rect 450156 309496 453547 309498
rect 450156 309440 453486 309496
rect 453542 309440 453547 309496
rect 450156 309438 453547 309440
rect 453481 309435 453547 309438
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 128353 302698 128419 302701
rect 128353 302696 132020 302698
rect 128353 302640 128358 302696
rect 128414 302640 132020 302696
rect 128353 302638 132020 302640
rect 128353 302635 128419 302638
rect 452929 302426 452995 302429
rect 450156 302424 452995 302426
rect 450156 302368 452934 302424
rect 452990 302368 452995 302424
rect 450156 302366 452995 302368
rect 452929 302363 452995 302366
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 453389 295218 453455 295221
rect 450156 295216 453455 295218
rect 450156 295160 453394 295216
rect 453450 295160 453455 295216
rect 450156 295158 453455 295160
rect 453389 295155 453455 295158
rect 129365 295082 129431 295085
rect 129365 295080 132020 295082
rect 129365 295024 129370 295080
rect 129426 295024 132020 295080
rect 129365 295022 132020 295024
rect 129365 295019 129431 295022
rect -960 294402 480 294492
rect 3509 294402 3575 294405
rect -960 294400 3575 294402
rect -960 294344 3514 294400
rect 3570 294344 3575 294400
rect -960 294342 3575 294344
rect -960 294252 480 294342
rect 3509 294339 3575 294342
rect 453297 288146 453363 288149
rect 450156 288144 453363 288146
rect 450156 288088 453302 288144
rect 453358 288088 453363 288144
rect 450156 288086 453363 288088
rect 453297 288083 453363 288086
rect 128353 287466 128419 287469
rect 128353 287464 132020 287466
rect 128353 287408 128358 287464
rect 128414 287408 132020 287464
rect 128353 287406 132020 287408
rect 128353 287403 128419 287406
rect 583520 287316 584960 287556
rect 453021 281074 453087 281077
rect 450156 281072 453087 281074
rect 450156 281016 453026 281072
rect 453082 281016 453087 281072
rect 450156 281014 453087 281016
rect 453021 281011 453087 281014
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 129089 279850 129155 279853
rect 129089 279848 132020 279850
rect 129089 279792 129094 279848
rect 129150 279792 132020 279848
rect 129089 279790 132020 279792
rect 129089 279787 129155 279790
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 453665 273866 453731 273869
rect 450156 273864 453731 273866
rect 450156 273808 453670 273864
rect 453726 273808 453731 273864
rect 450156 273806 453731 273808
rect 453665 273803 453731 273806
rect 129273 272098 129339 272101
rect 129273 272096 132020 272098
rect 129273 272040 129278 272096
rect 129334 272040 132020 272096
rect 129273 272038 132020 272040
rect 129273 272035 129339 272038
rect 453573 266794 453639 266797
rect 450156 266792 453639 266794
rect 450156 266736 453578 266792
rect 453634 266736 453639 266792
rect 450156 266734 453639 266736
rect 453573 266731 453639 266734
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 128353 264482 128419 264485
rect 128353 264480 132020 264482
rect 128353 264424 128358 264480
rect 128414 264424 132020 264480
rect 128353 264422 132020 264424
rect 128353 264419 128419 264422
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 453941 259722 454007 259725
rect 450156 259720 454007 259722
rect 450156 259664 453946 259720
rect 454002 259664 454007 259720
rect 450156 259662 454007 259664
rect 453941 259659 454007 259662
rect 128353 256866 128419 256869
rect 128353 256864 132020 256866
rect 128353 256808 128358 256864
rect 128414 256808 132020 256864
rect 128353 256806 132020 256808
rect 128353 256803 128419 256806
rect 452837 252514 452903 252517
rect 450156 252512 452903 252514
rect 450156 252456 452842 252512
rect 452898 252456 452903 252512
rect 450156 252454 452903 252456
rect 452837 252451 452903 252454
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 129181 249250 129247 249253
rect 129181 249248 132020 249250
rect 129181 249192 129186 249248
rect 129242 249192 132020 249248
rect 129181 249190 132020 249192
rect 129181 249187 129247 249190
rect 453481 245442 453547 245445
rect 450156 245440 453547 245442
rect 450156 245384 453486 245440
rect 453542 245384 453547 245440
rect 450156 245382 453547 245384
rect 453481 245379 453547 245382
rect 128353 241634 128419 241637
rect 128353 241632 132020 241634
rect 128353 241576 128358 241632
rect 128414 241576 132020 241632
rect 128353 241574 132020 241576
rect 128353 241571 128419 241574
rect 583520 240396 584960 240636
rect 453941 238370 454007 238373
rect 450156 238368 454007 238370
rect 450156 238312 453946 238368
rect 454002 238312 454007 238368
rect 450156 238310 454007 238312
rect 453941 238307 454007 238310
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 128353 234018 128419 234021
rect 128353 234016 132020 234018
rect 128353 233960 128358 234016
rect 128414 233960 132020 234016
rect 128353 233958 132020 233960
rect 128353 233955 128419 233958
rect 453113 231162 453179 231165
rect 450156 231160 453179 231162
rect 450156 231104 453118 231160
rect 453174 231104 453179 231160
rect 450156 231102 453179 231104
rect 453113 231099 453179 231102
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 129089 226402 129155 226405
rect 129089 226400 132020 226402
rect 129089 226344 129094 226400
rect 129150 226344 132020 226400
rect 129089 226342 132020 226344
rect 129089 226339 129155 226342
rect 453389 224090 453455 224093
rect 450156 224088 453455 224090
rect 450156 224032 453394 224088
rect 453450 224032 453455 224088
rect 450156 224030 453455 224032
rect 453389 224027 453455 224030
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 128353 218786 128419 218789
rect 128353 218784 132020 218786
rect 128353 218728 128358 218784
rect 128414 218728 132020 218784
rect 128353 218726 132020 218728
rect 128353 218723 128419 218726
rect 452929 217018 452995 217021
rect 450156 217016 452995 217018
rect 450156 216960 452934 217016
rect 452990 216960 452995 217016
rect 450156 216958 452995 216960
rect 452929 216955 452995 216958
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 128353 211170 128419 211173
rect 128353 211168 132020 211170
rect 128353 211112 128358 211168
rect 128414 211112 132020 211168
rect 128353 211110 132020 211112
rect 128353 211107 128419 211110
rect 453941 209810 454007 209813
rect 450156 209808 454007 209810
rect 450156 209752 453946 209808
rect 454002 209752 454007 209808
rect 450156 209750 454007 209752
rect 453941 209747 454007 209750
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 128997 203554 129063 203557
rect 128997 203552 132020 203554
rect 128997 203496 129002 203552
rect 129058 203496 132020 203552
rect 128997 203494 132020 203496
rect 128997 203491 129063 203494
rect 453297 202738 453363 202741
rect 450156 202736 453363 202738
rect 450156 202680 453302 202736
rect 453358 202680 453363 202736
rect 450156 202678 453363 202680
rect 453297 202675 453363 202678
rect 128629 195938 128695 195941
rect 128629 195936 132020 195938
rect 128629 195880 128634 195936
rect 128690 195880 132020 195936
rect 128629 195878 132020 195880
rect 128629 195875 128695 195878
rect 453941 195666 454007 195669
rect 450156 195664 454007 195666
rect 450156 195608 453946 195664
rect 454002 195608 454007 195664
rect 450156 195606 454007 195608
rect 453941 195603 454007 195606
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 135345 183562 135411 183565
rect 135529 183562 135595 183565
rect 135345 183560 135595 183562
rect 135345 183504 135350 183560
rect 135406 183504 135534 183560
rect 135590 183504 135595 183560
rect 135345 183502 135595 183504
rect 135345 183499 135411 183502
rect 135529 183499 135595 183502
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 135345 154594 135411 154597
rect 135621 154594 135687 154597
rect 135345 154592 135687 154594
rect 135345 154536 135350 154592
rect 135406 154536 135626 154592
rect 135682 154536 135687 154592
rect 135345 154534 135687 154536
rect 135345 154531 135411 154534
rect 135621 154531 135687 154534
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 135345 135282 135411 135285
rect 135621 135282 135687 135285
rect 135345 135280 135687 135282
rect 135345 135224 135350 135280
rect 135406 135224 135626 135280
rect 135682 135224 135687 135280
rect 135345 135222 135687 135224
rect 135345 135219 135411 135222
rect 135621 135219 135687 135222
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 135345 115970 135411 115973
rect 135621 115970 135687 115973
rect 135345 115968 135687 115970
rect 135345 115912 135350 115968
rect 135406 115912 135626 115968
rect 135682 115912 135687 115968
rect 135345 115910 135687 115912
rect 135345 115907 135411 115910
rect 135621 115907 135687 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect 135345 96658 135411 96661
rect 135621 96658 135687 96661
rect 135345 96656 135687 96658
rect 135345 96600 135350 96656
rect 135406 96600 135626 96656
rect 135682 96600 135687 96656
rect 135345 96598 135687 96600
rect 135345 96595 135411 96598
rect 135621 96595 135687 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 514437 145404 541898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 514437 163404 523898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 514437 181404 541898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 514437 199404 523898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 514437 217404 541898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 514437 235404 523898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 514437 253404 541898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 514437 271404 523898
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 514437 289404 541898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 514437 307404 523898
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 514437 325404 541898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 514437 343404 523898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 514437 361404 541898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 514437 379404 523898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 514437 397404 541898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 514437 415404 523898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 514437 433404 541898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 514437 451404 523898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 136208 506454 136528 506476
rect 136208 506218 136250 506454
rect 136486 506218 136528 506454
rect 136208 506134 136528 506218
rect 136208 505898 136250 506134
rect 136486 505898 136528 506134
rect 136208 505876 136528 505898
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 151568 488454 151888 488476
rect 151568 488218 151610 488454
rect 151846 488218 151888 488454
rect 151568 488134 151888 488218
rect 151568 487898 151610 488134
rect 151846 487898 151888 488134
rect 151568 487876 151888 487898
rect 136208 470454 136528 470476
rect 136208 470218 136250 470454
rect 136486 470218 136528 470454
rect 136208 470134 136528 470218
rect 136208 469898 136250 470134
rect 136486 469898 136528 470134
rect 136208 469876 136528 469898
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 151568 452454 151888 452476
rect 151568 452218 151610 452454
rect 151846 452218 151888 452454
rect 151568 452134 151888 452218
rect 151568 451898 151610 452134
rect 151846 451898 151888 452134
rect 151568 451876 151888 451898
rect 136208 434454 136528 434476
rect 136208 434218 136250 434454
rect 136486 434218 136528 434454
rect 136208 434134 136528 434218
rect 136208 433898 136250 434134
rect 136486 433898 136528 434134
rect 136208 433876 136528 433898
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 151568 416454 151888 416476
rect 151568 416218 151610 416454
rect 151846 416218 151888 416454
rect 151568 416134 151888 416218
rect 151568 415898 151610 416134
rect 151846 415898 151888 416134
rect 151568 415876 151888 415898
rect 136208 398454 136528 398476
rect 136208 398218 136250 398454
rect 136486 398218 136528 398454
rect 136208 398134 136528 398218
rect 136208 397898 136250 398134
rect 136486 397898 136528 398134
rect 136208 397876 136528 397898
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 151568 380454 151888 380476
rect 151568 380218 151610 380454
rect 151846 380218 151888 380454
rect 151568 380134 151888 380218
rect 151568 379898 151610 380134
rect 151846 379898 151888 380134
rect 151568 379876 151888 379898
rect 136208 362454 136528 362476
rect 136208 362218 136250 362454
rect 136486 362218 136528 362454
rect 136208 362134 136528 362218
rect 136208 361898 136250 362134
rect 136486 361898 136528 362134
rect 136208 361876 136528 361898
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 151568 344454 151888 344476
rect 151568 344218 151610 344454
rect 151846 344218 151888 344454
rect 151568 344134 151888 344218
rect 151568 343898 151610 344134
rect 151846 343898 151888 344134
rect 151568 343876 151888 343898
rect 136208 326454 136528 326476
rect 136208 326218 136250 326454
rect 136486 326218 136528 326454
rect 136208 326134 136528 326218
rect 136208 325898 136250 326134
rect 136486 325898 136528 326134
rect 136208 325876 136528 325898
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 151568 308454 151888 308476
rect 151568 308218 151610 308454
rect 151846 308218 151888 308454
rect 151568 308134 151888 308218
rect 151568 307898 151610 308134
rect 151846 307898 151888 308134
rect 151568 307876 151888 307898
rect 136208 290454 136528 290476
rect 136208 290218 136250 290454
rect 136486 290218 136528 290454
rect 136208 290134 136528 290218
rect 136208 289898 136250 290134
rect 136486 289898 136528 290134
rect 136208 289876 136528 289898
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 151568 272454 151888 272476
rect 151568 272218 151610 272454
rect 151846 272218 151888 272454
rect 151568 272134 151888 272218
rect 151568 271898 151610 272134
rect 151846 271898 151888 272134
rect 151568 271876 151888 271898
rect 136208 254454 136528 254476
rect 136208 254218 136250 254454
rect 136486 254218 136528 254454
rect 136208 254134 136528 254218
rect 136208 253898 136250 254134
rect 136486 253898 136528 254134
rect 136208 253876 136528 253898
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 151568 236454 151888 236476
rect 151568 236218 151610 236454
rect 151846 236218 151888 236454
rect 151568 236134 151888 236218
rect 151568 235898 151610 236134
rect 151846 235898 151888 236134
rect 151568 235876 151888 235898
rect 136208 218454 136528 218476
rect 136208 218218 136250 218454
rect 136486 218218 136528 218454
rect 136208 218134 136528 218218
rect 136208 217898 136250 218134
rect 136486 217898 136528 218134
rect 136208 217876 136528 217898
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 151568 200454 151888 200476
rect 151568 200218 151610 200454
rect 151846 200218 151888 200454
rect 151568 200134 151888 200218
rect 151568 199898 151610 200134
rect 151846 199898 151888 200134
rect 151568 199876 151888 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 182454 145404 190000
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 164454 163404 190000
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 182454 181404 190000
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 164454 199404 190000
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 182454 217404 190000
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 164454 235404 190000
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 182454 253404 190000
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 164454 271404 190000
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 182454 289404 190000
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 164454 307404 190000
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 182454 325404 190000
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 164454 343404 190000
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 182454 361404 190000
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 164454 379404 190000
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 182454 397404 190000
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 164454 415404 190000
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 182454 433404 190000
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 164454 451404 190000
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 136250 506218 136486 506454
rect 136250 505898 136486 506134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 151610 488218 151846 488454
rect 151610 487898 151846 488134
rect 136250 470218 136486 470454
rect 136250 469898 136486 470134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 151610 452218 151846 452454
rect 151610 451898 151846 452134
rect 136250 434218 136486 434454
rect 136250 433898 136486 434134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 151610 416218 151846 416454
rect 151610 415898 151846 416134
rect 136250 398218 136486 398454
rect 136250 397898 136486 398134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 151610 380218 151846 380454
rect 151610 379898 151846 380134
rect 136250 362218 136486 362454
rect 136250 361898 136486 362134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 151610 344218 151846 344454
rect 151610 343898 151846 344134
rect 136250 326218 136486 326454
rect 136250 325898 136486 326134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 151610 308218 151846 308454
rect 151610 307898 151846 308134
rect 136250 290218 136486 290454
rect 136250 289898 136486 290134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 151610 272218 151846 272454
rect 151610 271898 151846 272134
rect 136250 254218 136486 254454
rect 136250 253898 136486 254134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 151610 236218 151846 236454
rect 151610 235898 151846 236134
rect 136250 218218 136486 218454
rect 136250 217898 136486 218134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 151610 200218 151846 200454
rect 151610 199898 151846 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 136208 506476 136528 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 136250 506454
rect 136486 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 136250 506134
rect 136486 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 136208 505874 136528 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 151568 488476 151888 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 151610 488454
rect 151846 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 151610 488134
rect 151846 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 151568 487874 151888 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 136208 470476 136528 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 136250 470454
rect 136486 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 136250 470134
rect 136486 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 136208 469874 136528 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 151568 452476 151888 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 151610 452454
rect 151846 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 151610 452134
rect 151846 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 151568 451874 151888 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 136208 434476 136528 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 136250 434454
rect 136486 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 136250 434134
rect 136486 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 136208 433874 136528 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 151568 416476 151888 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 151610 416454
rect 151846 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 151610 416134
rect 151846 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 151568 415874 151888 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 136208 398476 136528 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 136250 398454
rect 136486 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 136250 398134
rect 136486 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 136208 397874 136528 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 151568 380476 151888 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 151610 380454
rect 151846 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 151610 380134
rect 151846 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 151568 379874 151888 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 136208 362476 136528 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 136250 362454
rect 136486 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 136250 362134
rect 136486 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 136208 361874 136528 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 151568 344476 151888 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 151610 344454
rect 151846 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 151610 344134
rect 151846 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 151568 343874 151888 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 136208 326476 136528 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 136250 326454
rect 136486 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 136250 326134
rect 136486 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 136208 325874 136528 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 151568 308476 151888 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 151610 308454
rect 151846 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 151610 308134
rect 151846 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 151568 307874 151888 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 136208 290476 136528 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 136250 290454
rect 136486 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 136250 290134
rect 136486 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 136208 289874 136528 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 151568 272476 151888 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 151610 272454
rect 151846 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 151610 272134
rect 151846 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 151568 271874 151888 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 136208 254476 136528 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 136250 254454
rect 136486 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 136250 254134
rect 136486 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 136208 253874 136528 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 151568 236476 151888 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 151610 236454
rect 151846 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 151610 236134
rect 151846 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 151568 235874 151888 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 136208 218476 136528 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 136250 218454
rect 136486 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 136250 218134
rect 136486 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 136208 217874 136528 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 151568 200476 151888 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 151610 200454
rect 151846 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 151610 200134
rect 151846 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 151568 199874 151888 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use Ibtida_top_dffram_cv  mprj
timestamp 1611548290
transform 1 0 132000 0 1 192000
box 0 0 318293 320437
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
