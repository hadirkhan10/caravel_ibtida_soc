magic
tech sky130A
magscale 1 2
timestamp 1607406405
<< locali >>
rect 72525 684607 72559 694093
rect 72801 676107 72835 684437
rect 170137 666587 170171 683077
rect 72985 647275 73019 656829
rect 72801 627963 72835 637517
rect 72985 608719 73019 618137
rect 122849 605999 122883 606645
rect 140697 606067 140731 606645
rect 97859 605965 97917 605999
rect 103379 605965 103437 605999
rect 142169 605999 142203 606101
rect 142353 605999 142387 606101
rect 142169 605965 142387 605999
rect 75837 602327 75871 605965
rect 103195 605829 103345 605863
rect 143549 603687 143583 606101
rect 150449 605795 150483 606033
rect 155233 605795 155267 606033
rect 91109 600423 91143 601273
rect 97917 600967 97951 601273
rect 105829 600355 105863 601273
rect 113189 600559 113223 601273
rect 123125 600899 123159 601273
rect 131037 600355 131071 601273
rect 183017 600423 183051 601273
rect 187341 600491 187375 601273
rect 215033 600559 215067 601273
rect 217609 600491 217643 601273
rect 271429 600695 271463 601273
rect 274465 600695 274499 601273
rect 95191 599981 95375 600015
rect 95341 599879 95375 599981
rect 113189 599879 113223 600049
rect 122757 599947 122791 600049
rect 143365 599947 143399 599981
rect 143549 599947 143583 600049
rect 124263 599913 124321 599947
rect 143365 599913 143457 599947
rect 146033 599947 146067 600049
rect 157935 599913 157993 599947
rect 160109 599879 160143 600117
rect 169769 600015 169803 600185
rect 179429 600015 179463 600117
rect 188997 599947 189031 600117
rect 202889 599947 202923 600049
rect 195839 599913 195897 599947
rect 212457 599947 212491 600049
rect 222209 599947 222243 600049
rect 215159 599913 215401 599947
rect 231777 599947 231811 600049
rect 241529 599947 241563 600049
rect 234479 599913 234721 599947
rect 251097 599947 251131 600049
rect 260849 599947 260883 600049
rect 253799 599913 254041 599947
rect 270417 599947 270451 600049
rect 270509 599947 270543 600117
rect 280077 600015 280111 600117
rect 283757 600015 283791 601273
rect 347973 600627 348007 601273
rect 365729 600627 365763 601273
rect 406577 600967 406611 603109
rect 407221 601647 407255 603653
rect 425161 600287 425195 601273
rect 437305 600831 437339 601273
rect 38669 599675 38703 599777
rect 22051 599641 22109 599675
rect 6193 599267 6227 599573
rect 9689 599471 9723 599573
rect 19257 599471 19291 599641
rect 31769 599539 31803 599641
rect 48237 599607 48271 599777
rect 51089 599539 51123 599641
rect 501521 599607 501555 603585
rect 504373 596207 504407 601749
rect 504373 531335 504407 534157
rect 504465 524331 504499 531233
rect 501613 510663 501647 520217
rect 504373 512023 504407 514777
rect 79241 496791 79275 501721
rect 82921 501619 82955 507841
rect 501613 498219 501647 507773
rect 512837 481695 512871 491249
rect 82921 469251 82955 474929
rect 512837 462383 512871 471937
rect 82829 441983 82863 444329
rect 82921 441711 82955 448545
rect 504373 434775 504407 444329
rect 512837 443003 512871 452489
rect 504373 415463 504407 425017
rect 512837 423691 512871 433245
rect 512837 404379 512871 413933
rect 82829 374799 82863 386257
rect 512837 385135 512871 394621
rect 512837 365755 512871 375241
rect 512837 346443 512871 355997
rect 82921 336855 82955 342465
rect 512837 327131 512871 336685
rect 82829 294287 82863 294729
rect 82921 294627 82955 299489
rect 82921 259471 82955 273785
rect 82829 217447 82863 219521
rect 82737 209831 82771 210681
rect 82829 207519 82863 209933
rect 82921 207723 82955 218977
rect 82737 172295 82771 173485
rect 82737 157403 82771 158661
rect 82829 158423 82863 173349
rect 82921 158015 82955 195245
rect 82645 144891 82679 148257
rect 82737 143599 82771 144993
rect 82829 143735 82863 145197
rect 82921 144823 82955 157845
rect 512837 153255 512871 162809
rect 82829 137207 82863 140233
rect 512837 133943 512871 143497
rect 82829 111027 82863 124185
rect 82921 118711 82955 124049
rect 51031 103105 51123 103139
rect 19349 102867 19383 102969
rect 38669 102799 38703 103105
rect 51089 103071 51123 103105
rect 56609 102799 56643 103037
rect 66177 102799 66211 102901
rect 9689 102595 9723 102697
rect 19257 102595 19291 102765
rect 80161 102459 80195 102493
rect 80011 102425 80195 102459
rect 82921 102323 82955 115209
rect 512837 114563 512871 124117
rect 416605 102833 416823 102867
rect 416605 102799 416639 102833
rect 416789 102799 416823 102833
rect 91293 102459 91327 102765
rect 86969 102391 87003 102425
rect 103529 102391 103563 102493
rect 104173 102459 104207 102765
rect 113833 102459 113867 102765
rect 120733 102459 120767 102765
rect 127357 102459 127391 102765
rect 142721 102459 142755 102765
rect 144929 102527 144963 102765
rect 153209 102391 153243 102493
rect 86969 102357 87061 102391
rect 115949 102187 115983 102357
rect 162777 102391 162811 102765
rect 162869 102527 162903 102765
rect 172529 102391 172563 102493
rect 182097 102391 182131 102765
rect 183569 102663 183603 102697
rect 193229 102663 193263 102765
rect 215251 102697 215309 102731
rect 183569 102629 183661 102663
rect 138029 102323 138063 102357
rect 137971 102289 138063 102323
rect 125609 102187 125643 102289
rect 183569 101847 183603 102561
rect 222209 102527 222243 102629
rect 226993 102527 227027 102697
rect 85037 100147 85071 100521
rect 280537 99331 280571 102697
rect 386337 102663 386371 102765
rect 394617 102663 394651 102765
rect 416697 102663 416731 102765
rect 356529 96679 356563 100249
rect 176703 96577 176853 96611
rect 212215 96577 212457 96611
rect 356471 96577 356621 96611
rect 176611 96509 176945 96543
rect 356379 96509 356713 96543
rect 212399 96441 212457 96475
rect 83289 89403 83323 95897
rect 86969 94707 87003 94809
rect 96537 94571 96571 94809
rect 115949 93279 115983 94605
rect 176761 89675 176795 96441
rect 512561 96339 512595 96509
rect 512653 95251 512687 104805
rect 512779 96577 512929 96611
rect 411177 87023 411211 93653
rect 79793 75939 79827 85493
rect 151553 77367 151587 81073
rect 198473 77299 198507 86921
rect 280445 77299 280479 86921
rect 212399 77197 212457 77231
rect 151461 67643 151495 77129
rect 176761 67643 176795 77129
rect 198473 67643 198507 77129
rect 356713 70295 356747 77129
rect 411177 67643 411211 77129
rect 512837 75939 512871 85493
rect 79885 50915 79919 57885
rect 83381 57851 83415 66181
rect 89913 48331 89947 57885
rect 140697 46971 140731 56525
rect 144745 48331 144779 57885
rect 176761 48331 176795 57885
rect 198473 48331 198507 57885
rect 212457 48331 212491 57885
rect 280353 48331 280387 57885
rect 333897 48331 333931 57885
rect 356621 48331 356655 57885
rect 411177 48331 411211 57885
rect 512837 56627 512871 66181
rect 140789 35955 140823 45509
rect 151553 38675 151587 48229
rect 210985 46971 211019 48297
rect 90005 29087 90039 31773
rect 144745 29019 144779 38573
rect 176761 31739 176795 38573
rect 198473 31671 198507 38573
rect 280353 31739 280387 38573
rect 512837 37315 512871 46869
rect 89821 21947 89855 27557
rect 140789 9707 140823 22661
rect 210985 19295 211019 27557
rect 144745 9707 144779 19261
rect 176853 9707 176887 19261
rect 212457 9707 212491 19261
rect 333897 9707 333931 19261
rect 338129 9707 338163 19261
rect 389189 9707 389223 19261
rect 391765 9707 391799 19261
rect 411177 9775 411211 19261
rect 488181 9707 488215 12461
rect 512469 9707 512503 27557
rect 73077 3451 73111 3689
rect 93869 3247 93903 4029
rect 103437 3247 103471 4029
rect 113189 3315 113223 4029
rect 122757 3315 122791 4029
rect 132509 3315 132543 4029
rect 146953 3315 146987 4029
rect 157349 3383 157383 4029
rect 253949 3383 253983 3621
rect 203901 595 203935 2805
rect 393053 595 393087 2805
rect 410901 595 410935 9605
rect 445677 6715 445711 9537
rect 496461 3383 496495 3893
rect 502441 595 502475 9605
rect 503729 3315 503763 4029
rect 508513 3927 508547 4029
<< viali >>
rect 72525 694093 72559 694127
rect 72525 684573 72559 684607
rect 72801 684437 72835 684471
rect 72801 676073 72835 676107
rect 170137 683077 170171 683111
rect 170137 666553 170171 666587
rect 72985 656829 73019 656863
rect 72985 647241 73019 647275
rect 72801 637517 72835 637551
rect 72801 627929 72835 627963
rect 72985 618137 73019 618171
rect 72985 608685 73019 608719
rect 122849 606645 122883 606679
rect 140697 606645 140731 606679
rect 140697 606033 140731 606067
rect 142169 606101 142203 606135
rect 75837 605965 75871 605999
rect 97825 605965 97859 605999
rect 97917 605965 97951 605999
rect 103345 605965 103379 605999
rect 103437 605965 103471 605999
rect 122849 605965 122883 605999
rect 142353 606101 142387 606135
rect 143549 606101 143583 606135
rect 103161 605829 103195 605863
rect 103345 605829 103379 605863
rect 150449 606033 150483 606067
rect 150449 605761 150483 605795
rect 155233 606033 155267 606067
rect 155233 605761 155267 605795
rect 143549 603653 143583 603687
rect 407221 603653 407255 603687
rect 75837 602293 75871 602327
rect 406577 603109 406611 603143
rect 91109 601273 91143 601307
rect 97917 601273 97951 601307
rect 97917 600933 97951 600967
rect 105829 601273 105863 601307
rect 91109 600389 91143 600423
rect 113189 601273 113223 601307
rect 123125 601273 123159 601307
rect 123125 600865 123159 600899
rect 131037 601273 131071 601307
rect 113189 600525 113223 600559
rect 105829 600321 105863 600355
rect 183017 601273 183051 601307
rect 187341 601273 187375 601307
rect 215033 601273 215067 601307
rect 215033 600525 215067 600559
rect 217609 601273 217643 601307
rect 187341 600457 187375 600491
rect 271429 601273 271463 601307
rect 271429 600661 271463 600695
rect 274465 601273 274499 601307
rect 274465 600661 274499 600695
rect 283757 601273 283791 601307
rect 217609 600457 217643 600491
rect 183017 600389 183051 600423
rect 131037 600321 131071 600355
rect 169769 600185 169803 600219
rect 160109 600117 160143 600151
rect 113189 600049 113223 600083
rect 95157 599981 95191 600015
rect 95341 599845 95375 599879
rect 122757 600049 122791 600083
rect 143549 600049 143583 600083
rect 143365 599981 143399 600015
rect 122757 599913 122791 599947
rect 124229 599913 124263 599947
rect 124321 599913 124355 599947
rect 143457 599913 143491 599947
rect 143549 599913 143583 599947
rect 146033 600049 146067 600083
rect 146033 599913 146067 599947
rect 157901 599913 157935 599947
rect 157993 599913 158027 599947
rect 113189 599845 113223 599879
rect 169769 599981 169803 600015
rect 179429 600117 179463 600151
rect 179429 599981 179463 600015
rect 188997 600117 189031 600151
rect 270509 600117 270543 600151
rect 202889 600049 202923 600083
rect 188997 599913 189031 599947
rect 195805 599913 195839 599947
rect 195897 599913 195931 599947
rect 202889 599913 202923 599947
rect 212457 600049 212491 600083
rect 222209 600049 222243 600083
rect 212457 599913 212491 599947
rect 215125 599913 215159 599947
rect 215401 599913 215435 599947
rect 222209 599913 222243 599947
rect 231777 600049 231811 600083
rect 241529 600049 241563 600083
rect 231777 599913 231811 599947
rect 234445 599913 234479 599947
rect 234721 599913 234755 599947
rect 241529 599913 241563 599947
rect 251097 600049 251131 600083
rect 260849 600049 260883 600083
rect 251097 599913 251131 599947
rect 253765 599913 253799 599947
rect 254041 599913 254075 599947
rect 260849 599913 260883 599947
rect 270417 600049 270451 600083
rect 270417 599913 270451 599947
rect 280077 600117 280111 600151
rect 280077 599981 280111 600015
rect 347973 601273 348007 601307
rect 347973 600593 348007 600627
rect 365729 601273 365763 601307
rect 407221 601613 407255 601647
rect 501521 603585 501555 603619
rect 406577 600933 406611 600967
rect 425161 601273 425195 601307
rect 365729 600593 365763 600627
rect 437305 601273 437339 601307
rect 437305 600797 437339 600831
rect 425161 600253 425195 600287
rect 283757 599981 283791 600015
rect 270509 599913 270543 599947
rect 160109 599845 160143 599879
rect 38669 599777 38703 599811
rect 19257 599641 19291 599675
rect 22017 599641 22051 599675
rect 22109 599641 22143 599675
rect 31769 599641 31803 599675
rect 38669 599641 38703 599675
rect 48237 599777 48271 599811
rect 6193 599573 6227 599607
rect 9689 599573 9723 599607
rect 9689 599437 9723 599471
rect 48237 599573 48271 599607
rect 51089 599641 51123 599675
rect 31769 599505 31803 599539
rect 501521 599573 501555 599607
rect 504373 601749 504407 601783
rect 51089 599505 51123 599539
rect 19257 599437 19291 599471
rect 6193 599233 6227 599267
rect 504373 596173 504407 596207
rect 504373 534157 504407 534191
rect 504373 531301 504407 531335
rect 504465 531233 504499 531267
rect 504465 524297 504499 524331
rect 501613 520217 501647 520251
rect 504373 514777 504407 514811
rect 504373 511989 504407 512023
rect 501613 510629 501647 510663
rect 82921 507841 82955 507875
rect 79241 501721 79275 501755
rect 82921 501585 82955 501619
rect 501613 507773 501647 507807
rect 501613 498185 501647 498219
rect 79241 496757 79275 496791
rect 512837 491249 512871 491283
rect 512837 481661 512871 481695
rect 82921 474929 82955 474963
rect 82921 469217 82955 469251
rect 512837 471937 512871 471971
rect 512837 462349 512871 462383
rect 512837 452489 512871 452523
rect 82921 448545 82955 448579
rect 82829 444329 82863 444363
rect 82829 441949 82863 441983
rect 82921 441677 82955 441711
rect 504373 444329 504407 444363
rect 512837 442969 512871 443003
rect 504373 434741 504407 434775
rect 512837 433245 512871 433279
rect 504373 425017 504407 425051
rect 512837 423657 512871 423691
rect 504373 415429 504407 415463
rect 512837 413933 512871 413967
rect 512837 404345 512871 404379
rect 512837 394621 512871 394655
rect 82829 386257 82863 386291
rect 512837 385101 512871 385135
rect 82829 374765 82863 374799
rect 512837 375241 512871 375275
rect 512837 365721 512871 365755
rect 512837 355997 512871 356031
rect 512837 346409 512871 346443
rect 82921 342465 82955 342499
rect 82921 336821 82955 336855
rect 512837 336685 512871 336719
rect 512837 327097 512871 327131
rect 82921 299489 82955 299523
rect 82829 294729 82863 294763
rect 82921 294593 82955 294627
rect 82829 294253 82863 294287
rect 82921 273785 82955 273819
rect 82921 259437 82955 259471
rect 82829 219521 82863 219555
rect 82829 217413 82863 217447
rect 82921 218977 82955 219011
rect 82737 210681 82771 210715
rect 82737 209797 82771 209831
rect 82829 209933 82863 209967
rect 82921 207689 82955 207723
rect 82829 207485 82863 207519
rect 82921 195245 82955 195279
rect 82737 173485 82771 173519
rect 82737 172261 82771 172295
rect 82829 173349 82863 173383
rect 82737 158661 82771 158695
rect 82829 158389 82863 158423
rect 82921 157981 82955 158015
rect 512837 162809 512871 162843
rect 82737 157369 82771 157403
rect 82921 157845 82955 157879
rect 82645 148257 82679 148291
rect 82829 145197 82863 145231
rect 82645 144857 82679 144891
rect 82737 144993 82771 145027
rect 512837 153221 512871 153255
rect 82921 144789 82955 144823
rect 82829 143701 82863 143735
rect 82737 143565 82771 143599
rect 512837 143497 512871 143531
rect 82829 140233 82863 140267
rect 82829 137173 82863 137207
rect 512837 133909 512871 133943
rect 82829 124185 82863 124219
rect 512837 124117 512871 124151
rect 82921 124049 82955 124083
rect 82921 118677 82955 118711
rect 82829 110993 82863 111027
rect 82921 115209 82955 115243
rect 38669 103105 38703 103139
rect 50997 103105 51031 103139
rect 19349 102969 19383 103003
rect 19349 102833 19383 102867
rect 51089 103037 51123 103071
rect 56609 103037 56643 103071
rect 19257 102765 19291 102799
rect 38669 102765 38703 102799
rect 56609 102765 56643 102799
rect 66177 102901 66211 102935
rect 66177 102765 66211 102799
rect 9689 102697 9723 102731
rect 9689 102561 9723 102595
rect 19257 102561 19291 102595
rect 80161 102493 80195 102527
rect 79977 102425 80011 102459
rect 512837 114529 512871 114563
rect 512653 104805 512687 104839
rect 91293 102765 91327 102799
rect 104173 102765 104207 102799
rect 86969 102425 87003 102459
rect 91293 102425 91327 102459
rect 103529 102493 103563 102527
rect 104173 102425 104207 102459
rect 113833 102765 113867 102799
rect 113833 102425 113867 102459
rect 120733 102765 120767 102799
rect 120733 102425 120767 102459
rect 127357 102765 127391 102799
rect 127357 102425 127391 102459
rect 142721 102765 142755 102799
rect 144929 102765 144963 102799
rect 162777 102765 162811 102799
rect 144929 102493 144963 102527
rect 153209 102493 153243 102527
rect 142721 102425 142755 102459
rect 87061 102357 87095 102391
rect 103529 102357 103563 102391
rect 115949 102357 115983 102391
rect 82921 102289 82955 102323
rect 138029 102357 138063 102391
rect 153209 102357 153243 102391
rect 162869 102765 162903 102799
rect 182097 102765 182131 102799
rect 162869 102493 162903 102527
rect 172529 102493 172563 102527
rect 162777 102357 162811 102391
rect 172529 102357 172563 102391
rect 193229 102765 193263 102799
rect 183569 102697 183603 102731
rect 386337 102765 386371 102799
rect 215217 102697 215251 102731
rect 215309 102697 215343 102731
rect 226993 102697 227027 102731
rect 183661 102629 183695 102663
rect 193229 102629 193263 102663
rect 222209 102629 222243 102663
rect 182097 102357 182131 102391
rect 183569 102561 183603 102595
rect 115949 102153 115983 102187
rect 125609 102289 125643 102323
rect 137937 102289 137971 102323
rect 125609 102153 125643 102187
rect 222209 102493 222243 102527
rect 226993 102493 227027 102527
rect 280537 102697 280571 102731
rect 183569 101813 183603 101847
rect 85037 100521 85071 100555
rect 85037 100113 85071 100147
rect 386337 102629 386371 102663
rect 394617 102765 394651 102799
rect 416605 102765 416639 102799
rect 416697 102765 416731 102799
rect 416789 102765 416823 102799
rect 394617 102629 394651 102663
rect 416697 102629 416731 102663
rect 280537 99297 280571 99331
rect 356529 100249 356563 100283
rect 356529 96645 356563 96679
rect 176669 96577 176703 96611
rect 176853 96577 176887 96611
rect 212181 96577 212215 96611
rect 212457 96577 212491 96611
rect 356437 96577 356471 96611
rect 356621 96577 356655 96611
rect 176577 96509 176611 96543
rect 176945 96509 176979 96543
rect 356345 96509 356379 96543
rect 356713 96509 356747 96543
rect 512561 96509 512595 96543
rect 176761 96441 176795 96475
rect 212365 96441 212399 96475
rect 212457 96441 212491 96475
rect 83289 95897 83323 95931
rect 86969 94809 87003 94843
rect 86969 94673 87003 94707
rect 96537 94809 96571 94843
rect 96537 94537 96571 94571
rect 115949 94605 115983 94639
rect 115949 93245 115983 93279
rect 512561 96305 512595 96339
rect 512745 96577 512779 96611
rect 512929 96577 512963 96611
rect 512653 95217 512687 95251
rect 176761 89641 176795 89675
rect 411177 93653 411211 93687
rect 83289 89369 83323 89403
rect 411177 86989 411211 87023
rect 198473 86921 198507 86955
rect 79793 85493 79827 85527
rect 151553 81073 151587 81107
rect 151553 77333 151587 77367
rect 198473 77265 198507 77299
rect 280445 86921 280479 86955
rect 280445 77265 280479 77299
rect 512837 85493 512871 85527
rect 212365 77197 212399 77231
rect 212457 77197 212491 77231
rect 79793 75905 79827 75939
rect 151461 77129 151495 77163
rect 151461 67609 151495 67643
rect 176761 77129 176795 77163
rect 176761 67609 176795 67643
rect 198473 77129 198507 77163
rect 356713 77129 356747 77163
rect 356713 70261 356747 70295
rect 411177 77129 411211 77163
rect 198473 67609 198507 67643
rect 512837 75905 512871 75939
rect 411177 67609 411211 67643
rect 83381 66181 83415 66215
rect 79885 57885 79919 57919
rect 512837 66181 512871 66215
rect 83381 57817 83415 57851
rect 89913 57885 89947 57919
rect 79885 50881 79919 50915
rect 144745 57885 144779 57919
rect 89913 48297 89947 48331
rect 140697 56525 140731 56559
rect 144745 48297 144779 48331
rect 176761 57885 176795 57919
rect 176761 48297 176795 48331
rect 198473 57885 198507 57919
rect 212457 57885 212491 57919
rect 198473 48297 198507 48331
rect 210985 48297 211019 48331
rect 212457 48297 212491 48331
rect 280353 57885 280387 57919
rect 280353 48297 280387 48331
rect 333897 57885 333931 57919
rect 333897 48297 333931 48331
rect 356621 57885 356655 57919
rect 356621 48297 356655 48331
rect 411177 57885 411211 57919
rect 512837 56593 512871 56627
rect 411177 48297 411211 48331
rect 140697 46937 140731 46971
rect 151553 48229 151587 48263
rect 140789 45509 140823 45543
rect 210985 46937 211019 46971
rect 151553 38641 151587 38675
rect 512837 46869 512871 46903
rect 140789 35921 140823 35955
rect 144745 38573 144779 38607
rect 90005 31773 90039 31807
rect 90005 29053 90039 29087
rect 176761 38573 176795 38607
rect 176761 31705 176795 31739
rect 198473 38573 198507 38607
rect 280353 38573 280387 38607
rect 512837 37281 512871 37315
rect 280353 31705 280387 31739
rect 198473 31637 198507 31671
rect 144745 28985 144779 29019
rect 89821 27557 89855 27591
rect 210985 27557 211019 27591
rect 89821 21913 89855 21947
rect 140789 22661 140823 22695
rect 512469 27557 512503 27591
rect 140789 9673 140823 9707
rect 144745 19261 144779 19295
rect 144745 9673 144779 9707
rect 176853 19261 176887 19295
rect 210985 19261 211019 19295
rect 212457 19261 212491 19295
rect 176853 9673 176887 9707
rect 212457 9673 212491 9707
rect 333897 19261 333931 19295
rect 333897 9673 333931 9707
rect 338129 19261 338163 19295
rect 338129 9673 338163 9707
rect 389189 19261 389223 19295
rect 389189 9673 389223 9707
rect 391765 19261 391799 19295
rect 411177 19261 411211 19295
rect 411177 9741 411211 9775
rect 488181 12461 488215 12495
rect 391765 9673 391799 9707
rect 488181 9673 488215 9707
rect 512469 9673 512503 9707
rect 410901 9605 410935 9639
rect 93869 4029 93903 4063
rect 73077 3689 73111 3723
rect 73077 3417 73111 3451
rect 93869 3213 93903 3247
rect 103437 4029 103471 4063
rect 113189 4029 113223 4063
rect 113189 3281 113223 3315
rect 122757 4029 122791 4063
rect 122757 3281 122791 3315
rect 132509 4029 132543 4063
rect 132509 3281 132543 3315
rect 146953 4029 146987 4063
rect 157349 4029 157383 4063
rect 157349 3349 157383 3383
rect 253949 3621 253983 3655
rect 253949 3349 253983 3383
rect 146953 3281 146987 3315
rect 103437 3213 103471 3247
rect 203901 2805 203935 2839
rect 203901 561 203935 595
rect 393053 2805 393087 2839
rect 393053 561 393087 595
rect 502441 9605 502475 9639
rect 445677 9537 445711 9571
rect 445677 6681 445711 6715
rect 496461 3893 496495 3927
rect 496461 3349 496495 3383
rect 410901 561 410935 595
rect 503729 4029 503763 4063
rect 508513 4029 508547 4063
rect 508513 3893 508547 3927
rect 503729 3281 503763 3315
rect 502441 561 502475 595
<< metal1 >>
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 138658 700720 138664 700732
rect 137888 700692 138664 700720
rect 137888 700680 137894 700692
rect 138658 700680 138664 700692
rect 138716 700680 138722 700732
rect 70302 700612 70308 700664
rect 70360 700652 70366 700664
rect 154114 700652 154120 700664
rect 70360 700624 154120 700652
rect 70360 700612 70366 700624
rect 154114 700612 154120 700624
rect 154172 700612 154178 700664
rect 81342 700544 81348 700596
rect 81400 700584 81406 700596
rect 218974 700584 218980 700596
rect 81400 700556 218980 700584
rect 81400 700544 81406 700556
rect 218974 700544 218980 700556
rect 219032 700544 219038 700596
rect 75822 700476 75828 700528
rect 75880 700516 75886 700528
rect 235166 700516 235172 700528
rect 75880 700488 235172 700516
rect 75880 700476 75886 700488
rect 235166 700476 235172 700488
rect 235224 700476 235230 700528
rect 283834 700476 283840 700528
rect 283892 700516 283898 700528
rect 298738 700516 298744 700528
rect 283892 700488 298744 700516
rect 283892 700476 283898 700488
rect 298738 700476 298744 700488
rect 298796 700476 298802 700528
rect 332502 700476 332508 700528
rect 332560 700516 332566 700528
rect 520458 700516 520464 700528
rect 332560 700488 520464 700516
rect 332560 700476 332566 700488
rect 520458 700476 520464 700488
rect 520516 700476 520522 700528
rect 77202 700408 77208 700460
rect 77260 700448 77266 700460
rect 348786 700448 348792 700460
rect 77260 700420 348792 700448
rect 77260 700408 77266 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 364978 700408 364984 700460
rect 365036 700448 365042 700460
rect 509970 700448 509976 700460
rect 365036 700420 509976 700448
rect 365036 700408 365042 700420
rect 509970 700408 509976 700420
rect 510028 700408 510034 700460
rect 67450 700340 67456 700392
rect 67508 700380 67514 700392
rect 413646 700380 413652 700392
rect 67508 700352 413652 700380
rect 67508 700340 67514 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 68738 700272 68744 700324
rect 68796 700312 68802 700324
rect 462314 700312 462320 700324
rect 68796 700284 462320 700312
rect 68796 700272 68802 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 529198 700272 529204 700324
rect 529256 700312 529262 700324
rect 543458 700312 543464 700324
rect 529256 700284 543464 700312
rect 529256 700272 529262 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 543550 700272 543556 700324
rect 543608 700312 543614 700324
rect 559650 700312 559656 700324
rect 543608 700284 559656 700312
rect 543608 700272 543614 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 8110 700204 8116 700256
rect 8168 700244 8174 700256
rect 14458 700244 14464 700256
rect 8168 700216 14464 700244
rect 8168 700204 8174 700216
rect 14458 700204 14464 700216
rect 14516 700204 14522 700256
rect 397454 699932 397460 699984
rect 397512 699972 397518 699984
rect 398742 699972 398748 699984
rect 397512 699944 398748 699972
rect 397512 699932 397518 699944
rect 398742 699932 398748 699944
rect 398800 699932 398806 699984
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 40494 699660 40500 699712
rect 40552 699700 40558 699712
rect 43438 699700 43444 699712
rect 40552 699672 43444 699700
rect 40552 699660 40558 699672
rect 43438 699660 43444 699672
rect 43496 699660 43502 699712
rect 88334 699660 88340 699712
rect 88392 699700 88398 699712
rect 89162 699700 89168 699712
rect 88392 699672 89168 699700
rect 88392 699660 88398 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 104894 699660 104900 699712
rect 104952 699700 104958 699712
rect 105446 699700 105452 699712
rect 104952 699672 105452 699700
rect 104952 699660 104958 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 542998 699660 543004 699712
rect 543056 699700 543062 699712
rect 543550 699700 543556 699712
rect 543056 699672 543556 699700
rect 543056 699660 543062 699672
rect 543550 699660 543556 699672
rect 543608 699660 543614 699712
rect 259362 698912 259368 698964
rect 259420 698952 259426 698964
rect 300118 698952 300124 698964
rect 259420 698924 300124 698952
rect 259420 698912 259426 698924
rect 300118 698912 300124 698924
rect 300176 698912 300182 698964
rect 202782 697552 202788 697604
rect 202840 697592 202846 697604
rect 502334 697592 502340 697604
rect 202840 697564 502340 697592
rect 202840 697552 202846 697564
rect 502334 697552 502340 697564
rect 502392 697552 502398 697604
rect 169938 695444 169944 695496
rect 169996 695484 170002 695496
rect 170306 695484 170312 695496
rect 169996 695456 170312 695484
rect 169996 695444 170002 695456
rect 170306 695444 170312 695456
rect 170364 695444 170370 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 429194 692792 429200 692844
rect 429252 692832 429258 692844
rect 429930 692832 429936 692844
rect 429252 692804 429936 692832
rect 429252 692792 429258 692804
rect 429930 692792 429936 692804
rect 429988 692792 429994 692844
rect 477494 692792 477500 692844
rect 477552 692832 477558 692844
rect 478598 692832 478604 692844
rect 477552 692804 478604 692832
rect 477552 692792 477558 692804
rect 478598 692792 478604 692804
rect 478656 692792 478662 692844
rect 169938 687896 169944 687948
rect 169996 687936 170002 687948
rect 170122 687936 170128 687948
rect 169996 687908 170128 687936
rect 169996 687896 170002 687908
rect 170122 687896 170128 687908
rect 170180 687896 170186 687948
rect 522298 685856 522304 685908
rect 522356 685896 522362 685908
rect 580166 685896 580172 685908
rect 522356 685868 580172 685896
rect 522356 685856 522362 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 169754 683068 169760 683120
rect 169812 683108 169818 683120
rect 170125 683111 170183 683117
rect 170125 683108 170137 683111
rect 169812 683080 170137 683108
rect 169812 683068 169818 683080
rect 170125 683077 170137 683080
rect 170171 683077 170183 683111
rect 170125 683071 170183 683077
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 173894 673956 173900 674008
rect 173952 673996 173958 674008
rect 178310 673996 178316 674008
rect 173952 673968 178316 673996
rect 173952 673956 173958 673968
rect 178310 673956 178316 673968
rect 178368 673956 178374 674008
rect 154574 673752 154580 673804
rect 154632 673792 154638 673804
rect 162210 673792 162216 673804
rect 154632 673764 162216 673792
rect 154632 673752 154638 673764
rect 162210 673752 162216 673764
rect 162268 673752 162274 673804
rect 477494 673480 477500 673532
rect 477552 673520 477558 673532
rect 477678 673520 477684 673532
rect 477552 673492 477684 673520
rect 477552 673480 477558 673492
rect 477678 673480 477684 673492
rect 477736 673480 477742 673532
rect 429194 673412 429200 673464
rect 429252 673452 429258 673464
rect 429470 673452 429476 673464
rect 429252 673424 429476 673452
rect 429252 673412 429258 673424
rect 429470 673412 429476 673424
rect 429528 673412 429534 673464
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 502426 667944 502432 667956
rect 3476 667916 502432 667944
rect 3476 667904 3482 667916
rect 502426 667904 502432 667916
rect 502484 667904 502490 667956
rect 170125 666587 170183 666593
rect 170125 666553 170137 666587
rect 170171 666584 170183 666587
rect 170214 666584 170220 666596
rect 170171 666556 170220 666584
rect 170171 666553 170183 666556
rect 170125 666547 170183 666553
rect 170214 666544 170220 666556
rect 170272 666544 170278 666596
rect 72878 659608 72884 659660
rect 72936 659648 72942 659660
rect 73062 659648 73068 659660
rect 72936 659620 73068 659648
rect 72936 659608 72942 659620
rect 73062 659608 73068 659620
rect 73120 659608 73126 659660
rect 72973 656863 73031 656869
rect 72973 656829 72985 656863
rect 73019 656860 73031 656863
rect 73062 656860 73068 656872
rect 73019 656832 73068 656860
rect 73019 656829 73031 656832
rect 72973 656823 73031 656829
rect 73062 656820 73068 656832
rect 73120 656820 73126 656872
rect 477494 654100 477500 654152
rect 477552 654140 477558 654152
rect 477678 654140 477684 654152
rect 477552 654112 477684 654140
rect 477552 654100 477558 654112
rect 477678 654100 477684 654112
rect 477736 654100 477742 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 17218 652780 17224 652792
rect 3108 652752 17224 652780
rect 3108 652740 3114 652752
rect 17218 652740 17224 652752
rect 17276 652740 17282 652792
rect 177942 650020 177948 650072
rect 178000 650060 178006 650072
rect 580166 650060 580172 650072
rect 178000 650032 580172 650060
rect 178000 650020 178006 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 72970 647272 72976 647284
rect 72931 647244 72976 647272
rect 72970 647232 72976 647244
rect 73028 647232 73034 647284
rect 169938 647232 169944 647284
rect 169996 647272 170002 647284
rect 170030 647272 170036 647284
rect 169996 647244 170036 647272
rect 169996 647232 170002 647244
rect 170030 647232 170036 647244
rect 170088 647232 170094 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 72970 640404 72976 640416
rect 72804 640376 72976 640404
rect 72804 640280 72832 640376
rect 72970 640364 72976 640376
rect 73028 640364 73034 640416
rect 169938 640364 169944 640416
rect 169996 640404 170002 640416
rect 170030 640404 170036 640416
rect 169996 640376 170036 640404
rect 169996 640364 170002 640376
rect 170030 640364 170036 640376
rect 170088 640364 170094 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 72786 640228 72792 640280
rect 72844 640228 72850 640280
rect 515398 638936 515404 638988
rect 515456 638976 515462 638988
rect 580166 638976 580172 638988
rect 515456 638948 580172 638976
rect 515456 638936 515462 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 72786 637548 72792 637560
rect 72747 637520 72792 637548
rect 72786 637508 72792 637520
rect 72844 637508 72850 637560
rect 477494 634788 477500 634840
rect 477552 634828 477558 634840
rect 477678 634828 477684 634840
rect 477552 634800 477684 634828
rect 477552 634788 477558 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 169846 630640 169852 630692
rect 169904 630680 169910 630692
rect 170030 630680 170036 630692
rect 169904 630652 170036 630680
rect 169904 630640 169910 630652
rect 170030 630640 170036 630652
rect 170088 630640 170094 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 398742 628532 398748 628584
rect 398800 628572 398806 628584
rect 501598 628572 501604 628584
rect 398800 628544 501604 628572
rect 398800 628532 398806 628544
rect 501598 628532 501604 628544
rect 501656 628532 501662 628584
rect 72789 627963 72847 627969
rect 72789 627929 72801 627963
rect 72835 627960 72847 627963
rect 73062 627960 73068 627972
rect 72835 627932 73068 627960
rect 72835 627929 72847 627932
rect 72789 627923 72847 627929
rect 73062 627920 73068 627932
rect 73120 627920 73126 627972
rect 81710 626560 81716 626612
rect 81768 626600 81774 626612
rect 580166 626600 580172 626612
rect 81768 626572 580172 626600
rect 81768 626560 81774 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 55858 623812 55864 623824
rect 3476 623784 55864 623812
rect 3476 623772 3482 623784
rect 55858 623772 55864 623784
rect 55916 623772 55922 623824
rect 72970 618264 72976 618316
rect 73028 618304 73034 618316
rect 73062 618304 73068 618316
rect 73028 618276 73068 618304
rect 73028 618264 73034 618276
rect 73062 618264 73068 618276
rect 73120 618264 73126 618316
rect 72970 618168 72976 618180
rect 72931 618140 72976 618168
rect 72970 618128 72976 618140
rect 73028 618128 73034 618180
rect 79870 617516 79876 617568
rect 79928 617556 79934 617568
rect 477678 617556 477684 617568
rect 79928 617528 477684 617556
rect 79928 617516 79934 617528
rect 477678 617516 477684 617528
rect 477736 617516 477742 617568
rect 43438 616088 43444 616140
rect 43496 616128 43502 616140
rect 398834 616128 398840 616140
rect 43496 616100 398840 616128
rect 43496 616088 43502 616100
rect 398834 616088 398840 616100
rect 398892 616088 398898 616140
rect 138658 614728 138664 614780
rect 138716 614768 138722 614780
rect 382274 614768 382280 614780
rect 138716 614740 382280 614768
rect 138716 614728 138722 614740
rect 382274 614728 382280 614740
rect 382332 614728 382338 614780
rect 169754 611328 169760 611380
rect 169812 611368 169818 611380
rect 170030 611368 170036 611380
rect 169812 611340 170036 611368
rect 169812 611328 169818 611340
rect 170030 611328 170036 611340
rect 170088 611328 170094 611380
rect 429194 611328 429200 611380
rect 429252 611368 429258 611380
rect 429470 611368 429476 611380
rect 429252 611340 429476 611368
rect 429252 611328 429258 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 128354 610580 128360 610632
rect 128412 610620 128418 610632
rect 542998 610620 543004 610632
rect 128412 610592 543004 610620
rect 128412 610580 128418 610592
rect 542998 610580 543004 610592
rect 543056 610580 543062 610632
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 48958 610008 48964 610020
rect 3476 609980 48964 610008
rect 3476 609968 3482 609980
rect 48958 609968 48964 609980
rect 49016 609968 49022 610020
rect 72973 608719 73031 608725
rect 72973 608685 72985 608719
rect 73019 608716 73031 608719
rect 73062 608716 73068 608728
rect 73019 608688 73068 608716
rect 73019 608685 73031 608688
rect 72973 608679 73031 608685
rect 73062 608676 73068 608688
rect 73120 608676 73126 608728
rect 380434 608676 380440 608728
rect 380492 608716 380498 608728
rect 521838 608716 521844 608728
rect 380492 608688 521844 608716
rect 380492 608676 380498 608688
rect 521838 608676 521844 608688
rect 521896 608676 521902 608728
rect 57882 608608 57888 608660
rect 57940 608648 57946 608660
rect 313642 608648 313648 608660
rect 57940 608620 313648 608648
rect 57940 608608 57946 608620
rect 313642 608608 313648 608620
rect 313700 608608 313706 608660
rect 375466 608608 375472 608660
rect 375524 608648 375530 608660
rect 520366 608648 520372 608660
rect 375524 608620 520372 608648
rect 375524 608608 375530 608620
rect 520366 608608 520372 608620
rect 520424 608608 520430 608660
rect 501782 608540 501788 608592
rect 501840 608580 501846 608592
rect 501966 608580 501972 608592
rect 501840 608552 501972 608580
rect 501840 608540 501846 608552
rect 501966 608540 501972 608552
rect 502024 608540 502030 608592
rect 81618 607860 81624 607912
rect 81676 607900 81682 607912
rect 169754 607900 169760 607912
rect 81676 607872 169760 607900
rect 81676 607860 81682 607872
rect 169754 607860 169760 607872
rect 169812 607860 169818 607912
rect 298738 607860 298744 607912
rect 298796 607900 298802 607912
rect 338298 607900 338304 607912
rect 298796 607872 338304 607900
rect 298796 607860 298802 607872
rect 338298 607860 338304 607872
rect 338356 607860 338362 607912
rect 67542 607316 67548 607368
rect 67600 607356 67606 607368
rect 155586 607356 155592 607368
rect 67600 607328 155592 607356
rect 67600 607316 67606 607328
rect 155586 607316 155592 607328
rect 155644 607316 155650 607368
rect 372890 607316 372896 607368
rect 372948 607356 372954 607368
rect 521654 607356 521660 607368
rect 372948 607328 521660 607356
rect 372948 607316 372954 607328
rect 521654 607316 521660 607328
rect 521712 607316 521718 607368
rect 64782 607248 64788 607300
rect 64840 607288 64846 607300
rect 180242 607288 180248 607300
rect 64840 607260 180248 607288
rect 64840 607248 64846 607260
rect 180242 607248 180248 607260
rect 180300 607248 180306 607300
rect 353202 607248 353208 607300
rect 353260 607288 353266 607300
rect 504818 607288 504824 607300
rect 353260 607260 504824 607288
rect 353260 607248 353266 607260
rect 504818 607248 504824 607260
rect 504876 607248 504882 607300
rect 81250 607180 81256 607232
rect 81308 607220 81314 607232
rect 204898 607220 204904 607232
rect 81308 607192 204904 607220
rect 81308 607180 81314 607192
rect 204898 607180 204904 607192
rect 204956 607180 204962 607232
rect 340874 607180 340880 607232
rect 340932 607220 340938 607232
rect 505738 607220 505744 607232
rect 340932 607192 505744 607220
rect 340932 607180 340938 607192
rect 505738 607180 505744 607192
rect 505796 607180 505802 607232
rect 122837 606679 122895 606685
rect 122837 606645 122849 606679
rect 122883 606676 122895 606679
rect 140685 606679 140743 606685
rect 140685 606676 140697 606679
rect 122883 606648 140697 606676
rect 122883 606645 122895 606648
rect 122837 606639 122895 606645
rect 140685 606645 140697 606648
rect 140731 606645 140743 606679
rect 140685 606639 140743 606645
rect 69750 606568 69756 606620
rect 69808 606608 69814 606620
rect 461946 606608 461952 606620
rect 69808 606580 461952 606608
rect 69808 606568 69814 606580
rect 461946 606568 461952 606580
rect 462004 606568 462010 606620
rect 66162 606500 66168 606552
rect 66220 606540 66226 606552
rect 190178 606540 190184 606552
rect 66220 606512 190184 606540
rect 66220 606500 66226 606512
rect 190178 606500 190184 606512
rect 190236 606500 190242 606552
rect 61838 606432 61844 606484
rect 61896 606472 61902 606484
rect 224770 606472 224776 606484
rect 61896 606444 224776 606472
rect 61896 606432 61902 606444
rect 224770 606432 224776 606444
rect 224828 606432 224834 606484
rect 328546 606432 328552 606484
rect 328604 606472 328610 606484
rect 429194 606472 429200 606484
rect 328604 606444 429200 606472
rect 328604 606432 328610 606444
rect 429194 606432 429200 606444
rect 429252 606432 429258 606484
rect 61746 606364 61752 606416
rect 61804 606404 61810 606416
rect 244458 606404 244464 606416
rect 61804 606376 244464 606404
rect 61804 606364 61810 606376
rect 244458 606364 244464 606376
rect 244516 606364 244522 606416
rect 81158 606296 81164 606348
rect 81216 606336 81222 606348
rect 318610 606336 318616 606348
rect 81216 606308 318616 606336
rect 81216 606296 81222 606308
rect 318610 606296 318616 606308
rect 318668 606296 318674 606348
rect 471698 606296 471704 606348
rect 471756 606336 471762 606348
rect 514938 606336 514944 606348
rect 471756 606308 514944 606336
rect 471756 606296 471762 606308
rect 514938 606296 514944 606308
rect 514996 606296 515002 606348
rect 74258 606228 74264 606280
rect 74316 606268 74322 606280
rect 323578 606268 323584 606280
rect 74316 606240 323584 606268
rect 74316 606228 74322 606240
rect 323578 606228 323584 606240
rect 323636 606228 323642 606280
rect 390186 606228 390192 606280
rect 390244 606268 390250 606280
rect 520550 606268 520556 606280
rect 390244 606240 520556 606268
rect 390244 606228 390250 606240
rect 520550 606228 520556 606240
rect 520608 606228 520614 606280
rect 71590 606160 71596 606212
rect 71648 606200 71654 606212
rect 199930 606200 199936 606212
rect 71648 606172 199936 606200
rect 71648 606160 71654 606172
rect 199930 606160 199936 606172
rect 199988 606160 199994 606212
rect 209866 606160 209872 606212
rect 209924 606200 209930 606212
rect 554038 606200 554044 606212
rect 209924 606172 554044 606200
rect 209924 606160 209930 606172
rect 554038 606160 554044 606172
rect 554096 606160 554102 606212
rect 82078 606092 82084 606144
rect 82136 606132 82142 606144
rect 142157 606135 142215 606141
rect 142157 606132 142169 606135
rect 82136 606104 142169 606132
rect 82136 606092 82142 606104
rect 142157 606101 142169 606104
rect 142203 606101 142215 606135
rect 142157 606095 142215 606101
rect 142341 606135 142399 606141
rect 142341 606101 142353 606135
rect 142387 606132 142399 606135
rect 143537 606135 143595 606141
rect 143537 606132 143549 606135
rect 142387 606104 143549 606132
rect 142387 606101 142399 606104
rect 142341 606095 142399 606101
rect 143537 606101 143549 606104
rect 143583 606101 143595 606135
rect 143537 606095 143595 606101
rect 165338 606092 165344 606144
rect 165396 606132 165402 606144
rect 508498 606132 508504 606144
rect 165396 606104 508504 606132
rect 165396 606092 165402 606104
rect 508498 606092 508504 606104
rect 508556 606092 508562 606144
rect 140685 606067 140743 606073
rect 140685 606033 140697 606067
rect 140731 606064 140743 606067
rect 150437 606067 150495 606073
rect 150437 606064 150449 606067
rect 140731 606036 150449 606064
rect 140731 606033 140743 606036
rect 140685 606027 140743 606033
rect 150437 606033 150449 606036
rect 150483 606033 150495 606067
rect 150437 606027 150495 606033
rect 155221 606067 155279 606073
rect 155221 606033 155233 606067
rect 155267 606064 155279 606067
rect 167914 606064 167920 606076
rect 155267 606036 167920 606064
rect 155267 606033 155279 606036
rect 155221 606027 155279 606033
rect 167914 606024 167920 606036
rect 167972 606024 167978 606076
rect 456978 606024 456984 606076
rect 457036 606064 457042 606076
rect 517790 606064 517796 606076
rect 457036 606036 517796 606064
rect 457036 606024 457042 606036
rect 517790 606024 517796 606036
rect 517848 606024 517854 606076
rect 75825 605999 75883 606005
rect 75825 605965 75837 605999
rect 75871 605996 75883 605999
rect 97813 605999 97871 606005
rect 97813 605996 97825 605999
rect 75871 605968 97825 605996
rect 75871 605965 75883 605968
rect 75825 605959 75883 605965
rect 97813 605965 97825 605968
rect 97859 605965 97871 605999
rect 97813 605959 97871 605965
rect 97905 605999 97963 606005
rect 97905 605965 97917 605999
rect 97951 605996 97963 605999
rect 103333 605999 103391 606005
rect 103333 605996 103345 605999
rect 97951 605968 103345 605996
rect 97951 605965 97963 605968
rect 97905 605959 97963 605965
rect 103333 605965 103345 605968
rect 103379 605965 103391 605999
rect 103333 605959 103391 605965
rect 103425 605999 103483 606005
rect 103425 605965 103437 605999
rect 103471 605996 103483 605999
rect 122837 605999 122895 606005
rect 122837 605996 122849 605999
rect 103471 605968 122849 605996
rect 103471 605965 103483 605968
rect 103425 605959 103483 605965
rect 122837 605965 122849 605968
rect 122883 605965 122895 605999
rect 122837 605959 122895 605965
rect 168282 605956 168288 606008
rect 168340 605996 168346 606008
rect 573358 605996 573364 606008
rect 168340 605968 573364 605996
rect 168340 605956 168346 605968
rect 573358 605956 573364 605968
rect 573416 605956 573422 606008
rect 86402 605888 86408 605940
rect 86460 605928 86466 605940
rect 523034 605928 523040 605940
rect 86460 605900 523040 605928
rect 86460 605888 86466 605900
rect 523034 605888 523040 605900
rect 523092 605888 523098 605940
rect 39390 605820 39396 605872
rect 39448 605860 39454 605872
rect 103149 605863 103207 605869
rect 103149 605860 103161 605863
rect 39448 605832 103161 605860
rect 39448 605820 39454 605832
rect 103149 605829 103161 605832
rect 103195 605829 103207 605863
rect 103149 605823 103207 605829
rect 103333 605863 103391 605869
rect 103333 605829 103345 605863
rect 103379 605860 103391 605863
rect 503898 605860 503904 605872
rect 103379 605832 503904 605860
rect 103379 605829 103391 605832
rect 103333 605823 103391 605829
rect 503898 605820 503904 605832
rect 503956 605820 503962 605872
rect 150437 605795 150495 605801
rect 150437 605761 150449 605795
rect 150483 605792 150495 605795
rect 155221 605795 155279 605801
rect 155221 605792 155233 605795
rect 150483 605764 155233 605792
rect 150483 605761 150495 605764
rect 150437 605755 150495 605761
rect 155221 605761 155233 605764
rect 155267 605761 155279 605795
rect 155221 605755 155279 605761
rect 72418 605276 72424 605328
rect 72476 605316 72482 605328
rect 246850 605316 246856 605328
rect 72476 605288 246856 605316
rect 72476 605276 72482 605288
rect 246850 605276 246856 605288
rect 246908 605276 246914 605328
rect 72970 605208 72976 605260
rect 73028 605248 73034 605260
rect 192570 605248 192576 605260
rect 73028 605220 192576 605248
rect 73028 605208 73034 605220
rect 192570 605208 192576 605220
rect 192628 605208 192634 605260
rect 82262 605140 82268 605192
rect 82320 605180 82326 605192
rect 360562 605180 360568 605192
rect 82320 605152 360568 605180
rect 82320 605140 82326 605152
rect 360562 605140 360568 605152
rect 360620 605140 360626 605192
rect 83274 605072 83280 605124
rect 83332 605112 83338 605124
rect 145650 605112 145656 605124
rect 83332 605084 145656 605112
rect 83332 605072 83338 605084
rect 145650 605072 145656 605084
rect 145708 605072 145714 605124
rect 79318 605004 79324 605056
rect 79376 605044 79382 605056
rect 160370 605044 160376 605056
rect 79376 605016 160376 605044
rect 79376 605004 79382 605016
rect 160370 605004 160376 605016
rect 160428 605004 160434 605056
rect 444650 605004 444656 605056
rect 444708 605044 444714 605056
rect 521746 605044 521752 605056
rect 444708 605016 521752 605044
rect 444708 605004 444714 605016
rect 521746 605004 521752 605016
rect 521804 605004 521810 605056
rect 67266 604936 67272 604988
rect 67324 604976 67330 604988
rect 222194 604976 222200 604988
rect 67324 604948 222200 604976
rect 67324 604936 67330 604948
rect 222194 604936 222200 604948
rect 222252 604936 222258 604988
rect 419810 604936 419816 604988
rect 419868 604976 419874 604988
rect 513558 604976 513564 604988
rect 419868 604948 513564 604976
rect 419868 604936 419874 604948
rect 513558 604936 513564 604948
rect 513616 604936 513622 604988
rect 57238 604868 57244 604920
rect 57296 604908 57302 604920
rect 276658 604908 276664 604920
rect 57296 604880 276664 604908
rect 57296 604868 57302 604880
rect 276658 604868 276664 604880
rect 276716 604868 276722 604920
rect 412450 604868 412456 604920
rect 412508 604908 412514 604920
rect 513374 604908 513380 604920
rect 412508 604880 513380 604908
rect 412508 604868 412514 604880
rect 513374 604868 513380 604880
rect 513432 604868 513438 604920
rect 21358 604800 21364 604852
rect 21416 604840 21422 604852
rect 256786 604840 256792 604852
rect 21416 604812 256792 604840
rect 21416 604800 21422 604812
rect 256786 604800 256792 604812
rect 256844 604800 256850 604852
rect 387794 604800 387800 604852
rect 387852 604840 387858 604852
rect 516410 604840 516416 604852
rect 387852 604812 516416 604840
rect 387852 604800 387858 604812
rect 516410 604800 516416 604812
rect 516468 604800 516474 604852
rect 79962 604732 79968 604784
rect 80020 604772 80026 604784
rect 325970 604772 325976 604784
rect 80020 604744 325976 604772
rect 80020 604732 80026 604744
rect 325970 604732 325976 604744
rect 326028 604732 326034 604784
rect 333330 604732 333336 604784
rect 333388 604772 333394 604784
rect 502978 604772 502984 604784
rect 333388 604744 502984 604772
rect 333388 604732 333394 604744
rect 502978 604732 502984 604744
rect 503036 604732 503042 604784
rect 68922 604664 68928 604716
rect 68980 604704 68986 604716
rect 101122 604704 101128 604716
rect 68980 604676 101128 604704
rect 68980 604664 68986 604676
rect 101122 604664 101128 604676
rect 101180 604664 101186 604716
rect 358170 604664 358176 604716
rect 358228 604704 358234 604716
rect 503806 604704 503812 604716
rect 358228 604676 503812 604704
rect 358228 604664 358234 604676
rect 503806 604664 503812 604676
rect 503864 604664 503870 604716
rect 242066 604596 242072 604648
rect 242124 604636 242130 604648
rect 554774 604636 554780 604648
rect 242124 604608 554780 604636
rect 242124 604596 242130 604608
rect 554774 604596 554780 604608
rect 554832 604596 554838 604648
rect 68278 604528 68284 604580
rect 68336 604568 68342 604580
rect 153010 604568 153016 604580
rect 68336 604540 153016 604568
rect 68336 604528 68342 604540
rect 153010 604528 153016 604540
rect 153068 604528 153074 604580
rect 172882 604528 172888 604580
rect 172940 604568 172946 604580
rect 514110 604568 514116 604580
rect 172940 604540 514116 604568
rect 172940 604528 172946 604540
rect 514110 604528 514116 604540
rect 514168 604528 514174 604580
rect 140682 604460 140688 604512
rect 140740 604500 140746 604512
rect 503714 604500 503720 604512
rect 140740 604472 503720 604500
rect 140740 604460 140746 604472
rect 503714 604460 503720 604472
rect 503772 604460 503778 604512
rect 289814 604052 289820 604104
rect 289872 604092 289878 604104
rect 299382 604092 299388 604104
rect 289872 604064 299388 604092
rect 289872 604052 289878 604064
rect 299382 604052 299388 604064
rect 299440 604052 299446 604104
rect 328454 604052 328460 604104
rect 328512 604092 328518 604104
rect 338022 604092 338028 604104
rect 328512 604064 338028 604092
rect 328512 604052 328518 604064
rect 338022 604052 338028 604064
rect 338080 604052 338086 604104
rect 347774 604052 347780 604104
rect 347832 604092 347838 604104
rect 357342 604092 357348 604104
rect 347832 604064 357348 604092
rect 347832 604052 347838 604064
rect 357342 604052 357348 604064
rect 357400 604052 357406 604104
rect 345842 603916 345848 603968
rect 345900 603956 345906 603968
rect 492674 603956 492680 603968
rect 345900 603928 492680 603956
rect 345900 603916 345906 603928
rect 492674 603916 492680 603928
rect 492732 603916 492738 603968
rect 64598 603848 64604 603900
rect 64656 603888 64662 603900
rect 98730 603888 98736 603900
rect 64656 603860 98736 603888
rect 64656 603848 64662 603860
rect 98730 603848 98736 603860
rect 98788 603848 98794 603900
rect 363138 603848 363144 603900
rect 363196 603888 363202 603900
rect 481726 603888 481732 603900
rect 363196 603860 481732 603888
rect 363196 603848 363202 603860
rect 481726 603848 481732 603860
rect 481784 603848 481790 603900
rect 483014 603848 483020 603900
rect 483072 603888 483078 603900
rect 492766 603888 492772 603900
rect 483072 603860 492772 603888
rect 483072 603848 483078 603860
rect 492766 603848 492772 603860
rect 492824 603848 492830 603900
rect 81434 603780 81440 603832
rect 81492 603820 81498 603832
rect 410058 603820 410064 603832
rect 81492 603792 410064 603820
rect 81492 603780 81498 603792
rect 410058 603780 410064 603792
rect 410116 603780 410122 603832
rect 452010 603780 452016 603832
rect 452068 603820 452074 603832
rect 502058 603820 502064 603832
rect 452068 603792 502064 603820
rect 452068 603780 452074 603792
rect 502058 603780 502064 603792
rect 502116 603780 502122 603832
rect 71038 603712 71044 603764
rect 71096 603752 71102 603764
rect 96154 603752 96160 603764
rect 71096 603724 96160 603752
rect 71096 603712 71102 603724
rect 96154 603712 96160 603724
rect 96212 603712 96218 603764
rect 190086 603712 190092 603764
rect 190144 603752 190150 603764
rect 417418 603752 417424 603764
rect 190144 603724 417424 603752
rect 190144 603712 190150 603724
rect 417418 603712 417424 603724
rect 417476 603712 417482 603764
rect 444466 603712 444472 603764
rect 444524 603752 444530 603764
rect 449158 603752 449164 603764
rect 444524 603724 449164 603752
rect 444524 603712 444530 603724
rect 449158 603712 449164 603724
rect 449216 603712 449222 603764
rect 454402 603712 454408 603764
rect 454460 603752 454466 603764
rect 513466 603752 513472 603764
rect 454460 603724 513472 603752
rect 454460 603712 454466 603724
rect 513466 603712 513472 603724
rect 513524 603712 513530 603764
rect 516870 603712 516876 603764
rect 516928 603752 516934 603764
rect 525702 603752 525708 603764
rect 516928 603724 525708 603752
rect 516928 603712 516934 603724
rect 525702 603712 525708 603724
rect 525760 603712 525766 603764
rect 79410 603644 79416 603696
rect 79468 603684 79474 603696
rect 108482 603684 108488 603696
rect 79468 603656 108488 603684
rect 79468 603644 79474 603656
rect 108482 603644 108488 603656
rect 108540 603644 108546 603696
rect 143537 603687 143595 603693
rect 143537 603653 143549 603687
rect 143583 603684 143595 603687
rect 148042 603684 148048 603696
rect 143583 603656 148048 603684
rect 143583 603653 143595 603656
rect 143537 603647 143595 603653
rect 148042 603644 148048 603656
rect 148100 603644 148106 603696
rect 309226 603644 309232 603696
rect 309284 603684 309290 603696
rect 318702 603684 318708 603696
rect 309284 603656 318708 603684
rect 309284 603644 309290 603656
rect 318702 603644 318708 603656
rect 318760 603644 318766 603696
rect 407209 603687 407267 603693
rect 407209 603653 407221 603687
rect 407255 603684 407267 603687
rect 469306 603684 469312 603696
rect 407255 603656 469312 603684
rect 407255 603653 407267 603656
rect 407209 603647 407267 603653
rect 469306 603644 469312 603656
rect 469364 603644 469370 603696
rect 479242 603644 479248 603696
rect 479300 603684 479306 603696
rect 502242 603684 502248 603696
rect 479300 603656 502248 603684
rect 479300 603644 479306 603656
rect 502242 603644 502248 603656
rect 502300 603644 502306 603696
rect 533982 603644 533988 603696
rect 534040 603684 534046 603696
rect 540882 603684 540888 603696
rect 534040 603656 540888 603684
rect 534040 603644 534046 603656
rect 540882 603644 540888 603656
rect 540940 603644 540946 603696
rect 71682 603576 71688 603628
rect 71740 603616 71746 603628
rect 125778 603616 125784 603628
rect 71740 603588 125784 603616
rect 71740 603576 71746 603588
rect 125778 603576 125784 603588
rect 125836 603576 125842 603628
rect 422386 603576 422392 603628
rect 422444 603616 422450 603628
rect 501509 603619 501567 603625
rect 501509 603616 501521 603619
rect 422444 603588 501521 603616
rect 422444 603576 422450 603588
rect 501509 603585 501521 603588
rect 501555 603585 501567 603619
rect 501509 603579 501567 603585
rect 56502 603508 56508 603560
rect 56560 603548 56566 603560
rect 111058 603548 111064 603560
rect 56560 603520 111064 603548
rect 56560 603508 56566 603520
rect 111058 603508 111064 603520
rect 111116 603508 111122 603560
rect 321002 603508 321008 603560
rect 321060 603548 321066 603560
rect 381446 603548 381452 603560
rect 321060 603520 381452 603548
rect 321060 603508 321066 603520
rect 381446 603508 381452 603520
rect 381504 603508 381510 603560
rect 432322 603508 432328 603560
rect 432380 603548 432386 603560
rect 515490 603548 515496 603560
rect 432380 603520 515496 603548
rect 432380 603508 432386 603520
rect 515490 603508 515496 603520
rect 515548 603508 515554 603560
rect 97902 603440 97908 603492
rect 97960 603480 97966 603492
rect 197538 603480 197544 603492
rect 97960 603452 197544 603480
rect 97960 603440 97966 603452
rect 197538 603440 197544 603452
rect 197596 603440 197602 603492
rect 351822 603440 351828 603492
rect 351880 603480 351886 603492
rect 466914 603480 466920 603492
rect 351880 603452 466920 603480
rect 351880 603440 351886 603452
rect 466914 603440 466920 603452
rect 466972 603440 466978 603492
rect 484210 603440 484216 603492
rect 484268 603480 484274 603492
rect 517606 603480 517612 603492
rect 484268 603452 517612 603480
rect 484268 603440 484274 603452
rect 517606 603440 517612 603452
rect 517664 603440 517670 603492
rect 67174 603372 67180 603424
rect 67232 603412 67238 603424
rect 202506 603412 202512 603424
rect 67232 603384 202512 603412
rect 67232 603372 67238 603384
rect 202506 603372 202512 603384
rect 202564 603372 202570 603424
rect 481634 603372 481640 603424
rect 481692 603412 481698 603424
rect 531958 603412 531964 603424
rect 481692 603384 531964 603412
rect 481692 603372 481698 603384
rect 531958 603372 531964 603384
rect 532016 603372 532022 603424
rect 64138 603304 64144 603356
rect 64196 603344 64202 603356
rect 150618 603344 150624 603356
rect 64196 603316 150624 603344
rect 64196 603304 64202 603316
rect 150618 603304 150624 603316
rect 150676 603304 150682 603356
rect 175274 603304 175280 603356
rect 175332 603344 175338 603356
rect 318794 603344 318800 603356
rect 175332 603316 318800 603344
rect 175332 603304 175338 603316
rect 318794 603304 318800 603316
rect 318852 603304 318858 603356
rect 493962 603304 493968 603356
rect 494020 603344 494026 603356
rect 516318 603344 516324 603356
rect 494020 603316 516324 603344
rect 494020 603304 494026 603316
rect 516318 603304 516324 603316
rect 516376 603304 516382 603356
rect 83182 603236 83188 603288
rect 83240 603276 83246 603288
rect 261754 603276 261760 603288
rect 83240 603248 261760 603276
rect 83240 603236 83246 603248
rect 261754 603236 261760 603248
rect 261812 603236 261818 603288
rect 343266 603236 343272 603288
rect 343324 603276 343330 603288
rect 512086 603276 512092 603288
rect 343324 603248 512092 603276
rect 343324 603236 343330 603248
rect 512086 603236 512092 603248
rect 512144 603236 512150 603288
rect 28258 603168 28264 603220
rect 28316 603208 28322 603220
rect 303706 603208 303712 603220
rect 28316 603180 303712 603208
rect 28316 603168 28322 603180
rect 303706 603168 303712 603180
rect 303764 603168 303770 603220
rect 311250 603168 311256 603220
rect 311308 603208 311314 603220
rect 552658 603208 552664 603220
rect 311308 603180 552664 603208
rect 311308 603168 311314 603180
rect 552658 603168 552664 603180
rect 552716 603168 552722 603220
rect 60550 603100 60556 603152
rect 60608 603140 60614 603152
rect 88794 603140 88800 603152
rect 60608 603112 88800 603140
rect 60608 603100 60614 603112
rect 88794 603100 88800 603112
rect 88852 603100 88858 603152
rect 301314 603100 301320 603152
rect 301372 603140 301378 603152
rect 346394 603140 346400 603152
rect 301372 603112 346400 603140
rect 301372 603100 301378 603112
rect 346394 603100 346400 603112
rect 346452 603100 346458 603152
rect 395154 603100 395160 603152
rect 395212 603140 395218 603152
rect 406565 603143 406623 603149
rect 406565 603140 406577 603143
rect 395212 603112 406577 603140
rect 395212 603100 395218 603112
rect 406565 603109 406577 603112
rect 406611 603109 406623 603143
rect 406565 603103 406623 603109
rect 407482 603100 407488 603152
rect 407540 603140 407546 603152
rect 507210 603140 507216 603152
rect 407540 603112 507216 603140
rect 407540 603100 407546 603112
rect 507210 603100 507216 603112
rect 507268 603100 507274 603152
rect 88334 603032 88340 603084
rect 88392 603072 88398 603084
rect 351822 603072 351828 603084
rect 88392 603044 351828 603072
rect 88392 603032 88398 603044
rect 351822 603032 351828 603044
rect 351880 603032 351886 603084
rect 492674 602760 492680 602812
rect 492732 602800 492738 602812
rect 498194 602800 498200 602812
rect 492732 602772 498200 602800
rect 492732 602760 492738 602772
rect 498194 602760 498200 602772
rect 498252 602760 498258 602812
rect 31662 602624 31668 602676
rect 31720 602664 31726 602676
rect 239490 602664 239496 602676
rect 31720 602636 239496 602664
rect 31720 602624 31726 602636
rect 239490 602624 239496 602636
rect 239548 602624 239554 602676
rect 70210 602556 70216 602608
rect 70268 602596 70274 602608
rect 232130 602596 232136 602608
rect 70268 602568 232136 602596
rect 70268 602556 70274 602568
rect 232130 602556 232136 602568
rect 232188 602556 232194 602608
rect 8938 602488 8944 602540
rect 8996 602528 9002 602540
rect 133322 602528 133328 602540
rect 8996 602500 133328 602528
rect 8996 602488 9002 602500
rect 133322 602488 133328 602500
rect 133380 602488 133386 602540
rect 59262 602420 59268 602472
rect 59320 602460 59326 602472
rect 59320 602432 68784 602460
rect 59320 602420 59326 602432
rect 68756 602324 68784 602432
rect 68830 602420 68836 602472
rect 68888 602460 68894 602472
rect 88242 602460 88248 602472
rect 68888 602432 88248 602460
rect 68888 602420 68894 602432
rect 88242 602420 88248 602432
rect 88300 602420 88306 602472
rect 481726 602420 481732 602472
rect 481784 602460 481790 602472
rect 517698 602460 517704 602472
rect 481784 602432 517704 602460
rect 481784 602420 481790 602432
rect 517698 602420 517704 602432
rect 517756 602420 517762 602472
rect 71498 602352 71504 602404
rect 71556 602392 71562 602404
rect 104802 602392 104808 602404
rect 71556 602364 104808 602392
rect 71556 602352 71562 602364
rect 104802 602352 104808 602364
rect 104860 602352 104866 602404
rect 381446 602352 381452 602404
rect 381504 602392 381510 602404
rect 580258 602392 580264 602404
rect 381504 602364 580264 602392
rect 381504 602352 381510 602364
rect 580258 602352 580264 602364
rect 580316 602352 580322 602404
rect 75825 602327 75883 602333
rect 75825 602324 75837 602327
rect 68756 602296 75837 602324
rect 75825 602293 75837 602296
rect 75871 602293 75883 602327
rect 75825 602287 75883 602293
rect 104894 602284 104900 602336
rect 104952 602324 104958 602336
rect 464338 602324 464344 602336
rect 104952 602296 464344 602324
rect 104952 602284 104958 602296
rect 464338 602284 464344 602296
rect 464396 602284 464402 602336
rect 82170 602216 82176 602268
rect 82228 602256 82234 602268
rect 143074 602256 143080 602268
rect 82228 602228 143080 602256
rect 82228 602216 82234 602228
rect 143074 602216 143080 602228
rect 143132 602216 143138 602268
rect 474274 602216 474280 602268
rect 474332 602256 474338 602268
rect 507854 602256 507860 602268
rect 474332 602228 507860 602256
rect 474332 602216 474338 602228
rect 507854 602216 507860 602228
rect 507912 602216 507918 602268
rect 74442 602148 74448 602200
rect 74500 602188 74506 602200
rect 135714 602188 135720 602200
rect 74500 602160 135720 602188
rect 74500 602148 74506 602160
rect 135714 602148 135720 602160
rect 135772 602148 135778 602200
rect 377858 602148 377864 602200
rect 377916 602188 377922 602200
rect 524414 602188 524420 602200
rect 377916 602160 524420 602188
rect 377916 602148 377922 602160
rect 524414 602148 524420 602160
rect 524472 602148 524478 602200
rect 9030 602080 9036 602132
rect 9088 602120 9094 602132
rect 120994 602120 121000 602132
rect 9088 602092 121000 602120
rect 9088 602080 9094 602092
rect 120994 602080 121000 602092
rect 121052 602080 121058 602132
rect 370498 602080 370504 602132
rect 370556 602120 370562 602132
rect 569954 602120 569960 602132
rect 370556 602092 569960 602120
rect 370556 602080 370562 602092
rect 569954 602080 569960 602092
rect 570012 602080 570018 602132
rect 83458 602012 83464 602064
rect 83516 602052 83522 602064
rect 226886 602052 226892 602064
rect 83516 602024 226892 602052
rect 83516 602012 83522 602024
rect 226886 602012 226892 602024
rect 226944 602012 226950 602064
rect 269482 602012 269488 602064
rect 269540 602052 269546 602064
rect 481818 602052 481824 602064
rect 269540 602024 481824 602052
rect 269540 602012 269546 602024
rect 481818 602012 481824 602024
rect 481876 602012 481882 602064
rect 27522 601944 27528 601996
rect 27580 601984 27586 601996
rect 263870 601984 263876 601996
rect 27580 601956 263876 601984
rect 27580 601944 27586 601956
rect 263870 601944 263876 601956
rect 263928 601944 263934 601996
rect 309042 601944 309048 601996
rect 309100 601984 309106 601996
rect 542998 601984 543004 601996
rect 309100 601956 543004 601984
rect 309100 601944 309106 601956
rect 542998 601944 543004 601956
rect 543056 601944 543062 601996
rect 237282 601876 237288 601928
rect 237340 601916 237346 601928
rect 514754 601916 514760 601928
rect 237340 601888 514760 601916
rect 237340 601876 237346 601888
rect 514754 601876 514760 601888
rect 514812 601876 514818 601928
rect 229922 601808 229928 601860
rect 229980 601848 229986 601860
rect 510614 601848 510620 601860
rect 229980 601820 510620 601848
rect 229980 601808 229986 601820
rect 510614 601808 510620 601820
rect 510672 601808 510678 601860
rect 72510 601740 72516 601792
rect 72568 601780 72574 601792
rect 115934 601780 115940 601792
rect 72568 601752 115940 601780
rect 72568 601740 72574 601752
rect 115934 601740 115940 601752
rect 115992 601740 115998 601792
rect 459554 601740 459560 601792
rect 459612 601780 459618 601792
rect 504361 601783 504419 601789
rect 504361 601780 504373 601783
rect 459612 601752 504373 601780
rect 459612 601740 459618 601752
rect 504361 601749 504373 601752
rect 504407 601749 504419 601783
rect 504361 601743 504419 601749
rect 118602 601672 118608 601724
rect 118660 601712 118666 601724
rect 507118 601712 507124 601724
rect 118660 601684 507124 601712
rect 118660 601672 118666 601684
rect 507118 601672 507124 601684
rect 507176 601672 507182 601724
rect 92382 601604 92388 601656
rect 92440 601644 92446 601656
rect 407209 601647 407267 601653
rect 407209 601644 407221 601647
rect 92440 601616 407221 601644
rect 92440 601604 92446 601616
rect 407209 601613 407221 601616
rect 407255 601613 407267 601647
rect 407209 601607 407267 601613
rect 504818 601332 504824 601384
rect 504876 601372 504882 601384
rect 507302 601372 507308 601384
rect 504876 601344 507308 601372
rect 504876 601332 504882 601344
rect 507302 601332 507308 601344
rect 507360 601332 507366 601384
rect 91094 601304 91100 601316
rect 91055 601276 91100 601304
rect 91094 601264 91100 601276
rect 91152 601264 91158 601316
rect 97902 601304 97908 601316
rect 97863 601276 97908 601304
rect 97902 601264 97908 601276
rect 97960 601264 97966 601316
rect 105814 601304 105820 601316
rect 105775 601276 105820 601304
rect 105814 601264 105820 601276
rect 105872 601264 105878 601316
rect 113174 601304 113180 601316
rect 113135 601276 113180 601304
rect 113174 601264 113180 601276
rect 113232 601264 113238 601316
rect 123110 601304 123116 601316
rect 123071 601276 123116 601304
rect 123110 601264 123116 601276
rect 123168 601264 123174 601316
rect 131022 601304 131028 601316
rect 130983 601276 131028 601304
rect 131022 601264 131028 601276
rect 131080 601264 131086 601316
rect 183002 601304 183008 601316
rect 182963 601276 183008 601304
rect 183002 601264 183008 601276
rect 183060 601264 183066 601316
rect 187326 601304 187332 601316
rect 187287 601276 187332 601304
rect 187326 601264 187332 601276
rect 187384 601264 187390 601316
rect 215018 601304 215024 601316
rect 214979 601276 215024 601304
rect 215018 601264 215024 601276
rect 215076 601264 215082 601316
rect 217594 601304 217600 601316
rect 217555 601276 217600 601304
rect 217594 601264 217600 601276
rect 217652 601264 217658 601316
rect 234246 601264 234252 601316
rect 234304 601264 234310 601316
rect 254210 601264 254216 601316
rect 254268 601264 254274 601316
rect 271414 601304 271420 601316
rect 271375 601276 271420 601304
rect 271414 601264 271420 601276
rect 271472 601264 271478 601316
rect 274450 601304 274456 601316
rect 274411 601276 274456 601304
rect 274450 601264 274456 601276
rect 274508 601264 274514 601316
rect 283742 601304 283748 601316
rect 283703 601276 283748 601304
rect 283742 601264 283748 601276
rect 283800 601264 283806 601316
rect 291194 601264 291200 601316
rect 291252 601264 291258 601316
rect 347958 601304 347964 601316
rect 347919 601276 347964 601304
rect 347958 601264 347964 601276
rect 348016 601264 348022 601316
rect 355870 601264 355876 601316
rect 355928 601264 355934 601316
rect 365714 601304 365720 601316
rect 365675 601276 365720 601304
rect 365714 601264 365720 601276
rect 365772 601264 365778 601316
rect 425146 601304 425152 601316
rect 425107 601276 425152 601304
rect 425146 601264 425152 601276
rect 425204 601264 425210 601316
rect 437290 601304 437296 601316
rect 437251 601276 437296 601304
rect 437290 601264 437296 601276
rect 437348 601264 437354 601316
rect 498194 601264 498200 601316
rect 498252 601304 498258 601316
rect 503990 601304 503996 601316
rect 498252 601276 503996 601304
rect 498252 601264 498258 601276
rect 503990 601264 503996 601276
rect 504048 601264 504054 601316
rect 83458 601060 83464 601112
rect 83516 601100 83522 601112
rect 83642 601100 83648 601112
rect 83516 601072 83648 601100
rect 83516 601060 83522 601072
rect 83642 601060 83648 601072
rect 83700 601060 83706 601112
rect 75546 600992 75552 601044
rect 75604 601032 75610 601044
rect 234264 601032 234292 601264
rect 75604 601004 234292 601032
rect 75604 600992 75610 601004
rect 81066 600924 81072 600976
rect 81124 600964 81130 600976
rect 97905 600967 97963 600973
rect 97905 600964 97917 600967
rect 81124 600936 97917 600964
rect 81124 600924 81130 600936
rect 97905 600933 97917 600936
rect 97951 600933 97963 600967
rect 97905 600927 97963 600933
rect 74350 600856 74356 600908
rect 74408 600896 74414 600908
rect 123113 600899 123171 600905
rect 123113 600896 123125 600899
rect 74408 600868 123125 600896
rect 74408 600856 74414 600868
rect 123113 600865 123125 600868
rect 123159 600865 123171 600899
rect 123113 600859 123171 600865
rect 71130 600788 71136 600840
rect 71188 600828 71194 600840
rect 254228 600828 254256 601264
rect 71188 600800 254256 600828
rect 71188 600788 71194 600800
rect 72878 600720 72884 600772
rect 72936 600760 72942 600772
rect 291212 600760 291240 601264
rect 72936 600732 291240 600760
rect 355888 600760 355916 601264
rect 406565 600967 406623 600973
rect 406565 600933 406577 600967
rect 406611 600964 406623 600967
rect 543734 600964 543740 600976
rect 406611 600936 543740 600964
rect 406611 600933 406623 600936
rect 406565 600927 406623 600933
rect 543734 600924 543740 600936
rect 543792 600924 543798 600976
rect 437293 600831 437351 600837
rect 437293 600797 437305 600831
rect 437339 600828 437351 600831
rect 509326 600828 509332 600840
rect 437339 600800 509332 600828
rect 437339 600797 437351 600800
rect 437293 600791 437351 600797
rect 509326 600788 509332 600800
rect 509384 600788 509390 600840
rect 511350 600760 511356 600772
rect 355888 600732 511356 600760
rect 72936 600720 72942 600732
rect 511350 600720 511356 600732
rect 511408 600720 511414 600772
rect 76558 600652 76564 600704
rect 76616 600692 76622 600704
rect 271417 600695 271475 600701
rect 271417 600692 271429 600695
rect 76616 600664 271429 600692
rect 76616 600652 76622 600664
rect 271417 600661 271429 600664
rect 271463 600661 271475 600695
rect 271417 600655 271475 600661
rect 274453 600695 274511 600701
rect 274453 600661 274465 600695
rect 274499 600692 274511 600695
rect 516226 600692 516232 600704
rect 274499 600664 516232 600692
rect 274499 600661 274511 600664
rect 274453 600655 274511 600661
rect 516226 600652 516232 600664
rect 516284 600652 516290 600704
rect 69658 600584 69664 600636
rect 69716 600624 69722 600636
rect 347961 600627 348019 600633
rect 347961 600624 347973 600627
rect 69716 600596 347973 600624
rect 69716 600584 69722 600596
rect 347961 600593 347973 600596
rect 348007 600593 348019 600627
rect 347961 600587 348019 600593
rect 365717 600627 365775 600633
rect 365717 600593 365729 600627
rect 365763 600624 365775 600627
rect 556154 600624 556160 600636
rect 365763 600596 556160 600624
rect 365763 600593 365775 600596
rect 365717 600587 365775 600593
rect 556154 600584 556160 600596
rect 556212 600584 556218 600636
rect 62022 600516 62028 600568
rect 62080 600556 62086 600568
rect 113177 600559 113235 600565
rect 113177 600556 113189 600559
rect 62080 600528 113189 600556
rect 62080 600516 62086 600528
rect 113177 600525 113189 600528
rect 113223 600525 113235 600559
rect 113177 600519 113235 600525
rect 215021 600559 215079 600565
rect 215021 600525 215033 600559
rect 215067 600556 215079 600559
rect 518158 600556 518164 600568
rect 215067 600528 518164 600556
rect 215067 600525 215079 600528
rect 215021 600519 215079 600525
rect 518158 600516 518164 600528
rect 518216 600516 518222 600568
rect 83642 600448 83648 600500
rect 83700 600488 83706 600500
rect 187329 600491 187387 600497
rect 187329 600488 187341 600491
rect 83700 600460 187341 600488
rect 83700 600448 83706 600460
rect 187329 600457 187341 600460
rect 187375 600457 187387 600491
rect 187329 600451 187387 600457
rect 217597 600491 217655 600497
rect 217597 600457 217609 600491
rect 217643 600488 217655 600491
rect 532694 600488 532700 600500
rect 217643 600460 532700 600488
rect 217643 600457 217655 600460
rect 217597 600451 217655 600457
rect 532694 600448 532700 600460
rect 532752 600448 532758 600500
rect 61930 600380 61936 600432
rect 61988 600420 61994 600432
rect 91097 600423 91155 600429
rect 91097 600420 91109 600423
rect 61988 600392 91109 600420
rect 61988 600380 61994 600392
rect 91097 600389 91109 600392
rect 91143 600389 91155 600423
rect 91097 600383 91155 600389
rect 183005 600423 183063 600429
rect 183005 600389 183017 600423
rect 183051 600420 183063 600423
rect 518894 600420 518900 600432
rect 183051 600392 518900 600420
rect 183051 600389 183063 600392
rect 183005 600383 183063 600389
rect 518894 600380 518900 600392
rect 518952 600380 518958 600432
rect 15838 600312 15844 600364
rect 15896 600352 15902 600364
rect 105817 600355 105875 600361
rect 105817 600352 105829 600355
rect 15896 600324 105829 600352
rect 15896 600312 15902 600324
rect 105817 600321 105829 600324
rect 105863 600321 105875 600355
rect 105817 600315 105875 600321
rect 131025 600355 131083 600361
rect 131025 600321 131037 600355
rect 131071 600352 131083 600355
rect 509878 600352 509884 600364
rect 131071 600324 509884 600352
rect 131071 600321 131083 600324
rect 131025 600315 131083 600321
rect 509878 600312 509884 600324
rect 509936 600312 509942 600364
rect 425149 600287 425207 600293
rect 425149 600253 425161 600287
rect 425195 600284 425207 600287
rect 501506 600284 501512 600296
rect 425195 600256 501512 600284
rect 425195 600253 425207 600256
rect 425149 600247 425207 600253
rect 501506 600244 501512 600256
rect 501564 600244 501570 600296
rect 169757 600219 169815 600225
rect 169757 600216 169769 600219
rect 169680 600188 169769 600216
rect 160097 600151 160155 600157
rect 160097 600117 160109 600151
rect 160143 600148 160155 600151
rect 169680 600148 169708 600188
rect 169757 600185 169769 600188
rect 169803 600185 169815 600219
rect 169757 600179 169815 600185
rect 160143 600120 169708 600148
rect 179417 600151 179475 600157
rect 160143 600117 160155 600120
rect 160097 600111 160155 600117
rect 179417 600117 179429 600151
rect 179463 600148 179475 600151
rect 188985 600151 189043 600157
rect 188985 600148 188997 600151
rect 179463 600120 188997 600148
rect 179463 600117 179475 600120
rect 179417 600111 179475 600117
rect 188985 600117 188997 600120
rect 189031 600117 189043 600151
rect 188985 600111 189043 600117
rect 270497 600151 270555 600157
rect 270497 600117 270509 600151
rect 270543 600148 270555 600151
rect 280065 600151 280123 600157
rect 280065 600148 280077 600151
rect 270543 600120 280077 600148
rect 270543 600117 270555 600120
rect 270497 600111 270555 600117
rect 280065 600117 280077 600120
rect 280111 600117 280123 600151
rect 280065 600111 280123 600117
rect 113177 600083 113235 600089
rect 113177 600049 113189 600083
rect 113223 600080 113235 600083
rect 122745 600083 122803 600089
rect 122745 600080 122757 600083
rect 113223 600052 122757 600080
rect 113223 600049 113235 600052
rect 113177 600043 113235 600049
rect 122745 600049 122757 600052
rect 122791 600049 122803 600083
rect 122745 600043 122803 600049
rect 143537 600083 143595 600089
rect 143537 600049 143549 600083
rect 143583 600080 143595 600083
rect 146021 600083 146079 600089
rect 146021 600080 146033 600083
rect 143583 600052 146033 600080
rect 143583 600049 143595 600052
rect 143537 600043 143595 600049
rect 146021 600049 146033 600052
rect 146067 600049 146079 600083
rect 146021 600043 146079 600049
rect 202877 600083 202935 600089
rect 202877 600049 202889 600083
rect 202923 600080 202935 600083
rect 212445 600083 212503 600089
rect 212445 600080 212457 600083
rect 202923 600052 212457 600080
rect 202923 600049 202935 600052
rect 202877 600043 202935 600049
rect 212445 600049 212457 600052
rect 212491 600049 212503 600083
rect 212445 600043 212503 600049
rect 222197 600083 222255 600089
rect 222197 600049 222209 600083
rect 222243 600080 222255 600083
rect 231765 600083 231823 600089
rect 231765 600080 231777 600083
rect 222243 600052 231777 600080
rect 222243 600049 222255 600052
rect 222197 600043 222255 600049
rect 231765 600049 231777 600052
rect 231811 600049 231823 600083
rect 231765 600043 231823 600049
rect 241517 600083 241575 600089
rect 241517 600049 241529 600083
rect 241563 600080 241575 600083
rect 251085 600083 251143 600089
rect 251085 600080 251097 600083
rect 241563 600052 251097 600080
rect 241563 600049 241575 600052
rect 241517 600043 241575 600049
rect 251085 600049 251097 600052
rect 251131 600049 251143 600083
rect 251085 600043 251143 600049
rect 260837 600083 260895 600089
rect 260837 600049 260849 600083
rect 260883 600080 260895 600083
rect 270405 600083 270463 600089
rect 270405 600080 270417 600083
rect 260883 600052 270417 600080
rect 260883 600049 260895 600052
rect 260837 600043 260895 600049
rect 270405 600049 270417 600052
rect 270451 600049 270463 600083
rect 270405 600043 270463 600049
rect 83458 600012 83464 600024
rect 75196 599984 83464 600012
rect 38657 599811 38715 599817
rect 38657 599777 38669 599811
rect 38703 599808 38715 599811
rect 48225 599811 48283 599817
rect 48225 599808 48237 599811
rect 38703 599780 48237 599808
rect 38703 599777 38715 599780
rect 38657 599771 38715 599777
rect 48225 599777 48237 599780
rect 48271 599777 48283 599811
rect 48225 599771 48283 599777
rect 60568 599712 62804 599740
rect 19245 599675 19303 599681
rect 19245 599641 19257 599675
rect 19291 599672 19303 599675
rect 22005 599675 22063 599681
rect 22005 599672 22017 599675
rect 19291 599644 22017 599672
rect 19291 599641 19303 599644
rect 19245 599635 19303 599641
rect 22005 599641 22017 599644
rect 22051 599641 22063 599675
rect 22005 599635 22063 599641
rect 22097 599675 22155 599681
rect 22097 599641 22109 599675
rect 22143 599672 22155 599675
rect 31757 599675 31815 599681
rect 22143 599644 23336 599672
rect 22143 599641 22155 599644
rect 22097 599635 22155 599641
rect 6181 599607 6239 599613
rect 6181 599573 6193 599607
rect 6227 599604 6239 599607
rect 9677 599607 9735 599613
rect 9677 599604 9689 599607
rect 6227 599576 9689 599604
rect 6227 599573 6239 599576
rect 6181 599567 6239 599573
rect 9677 599573 9689 599576
rect 9723 599573 9735 599607
rect 23308 599604 23336 599644
rect 31757 599641 31769 599675
rect 31803 599672 31815 599675
rect 38657 599675 38715 599681
rect 38657 599672 38669 599675
rect 31803 599644 38669 599672
rect 31803 599641 31815 599644
rect 31757 599635 31815 599641
rect 38657 599641 38669 599644
rect 38703 599641 38715 599675
rect 38657 599635 38715 599641
rect 51077 599675 51135 599681
rect 51077 599641 51089 599675
rect 51123 599672 51135 599675
rect 60568 599672 60596 599712
rect 51123 599644 60596 599672
rect 51123 599641 51135 599644
rect 51077 599635 51135 599641
rect 48225 599607 48283 599613
rect 23308 599576 31708 599604
rect 9677 599567 9735 599573
rect 31680 599536 31708 599576
rect 48225 599573 48237 599607
rect 48271 599604 48283 599607
rect 62776 599604 62804 599712
rect 75196 599604 75224 599984
rect 83458 599972 83464 599984
rect 83516 599972 83522 600024
rect 95145 600015 95203 600021
rect 95145 600012 95157 600015
rect 91756 599984 95157 600012
rect 91756 599876 91784 599984
rect 95145 599981 95157 599984
rect 95191 599981 95203 600015
rect 143353 600015 143411 600021
rect 143353 600012 143365 600015
rect 95145 599975 95203 599981
rect 138676 599984 143365 600012
rect 122745 599947 122803 599953
rect 122745 599913 122757 599947
rect 122791 599944 122803 599947
rect 124217 599947 124275 599953
rect 124217 599944 124229 599947
rect 122791 599916 124229 599944
rect 122791 599913 122803 599916
rect 122745 599907 122803 599913
rect 124217 599913 124229 599916
rect 124263 599913 124275 599947
rect 124217 599907 124275 599913
rect 124309 599947 124367 599953
rect 124309 599913 124321 599947
rect 124355 599944 124367 599947
rect 138676 599944 138704 599984
rect 143353 599981 143365 599984
rect 143399 599981 143411 600015
rect 143353 599975 143411 599981
rect 169757 600015 169815 600021
rect 169757 599981 169769 600015
rect 169803 600012 169815 600015
rect 179417 600015 179475 600021
rect 179417 600012 179429 600015
rect 169803 599984 179429 600012
rect 169803 599981 169815 599984
rect 169757 599975 169815 599981
rect 179417 599981 179429 599984
rect 179463 599981 179475 600015
rect 179417 599975 179475 599981
rect 280065 600015 280123 600021
rect 280065 599981 280077 600015
rect 280111 600012 280123 600015
rect 283745 600015 283803 600021
rect 283745 600012 283757 600015
rect 280111 599984 283757 600012
rect 280111 599981 280123 599984
rect 280065 599975 280123 599981
rect 283745 599981 283757 599984
rect 283791 599981 283803 600015
rect 283745 599975 283803 599981
rect 124355 599916 138704 599944
rect 143445 599947 143503 599953
rect 124355 599913 124367 599916
rect 124309 599907 124367 599913
rect 143445 599913 143457 599947
rect 143491 599944 143503 599947
rect 143537 599947 143595 599953
rect 143537 599944 143549 599947
rect 143491 599916 143549 599944
rect 143491 599913 143503 599916
rect 143445 599907 143503 599913
rect 143537 599913 143549 599916
rect 143583 599913 143595 599947
rect 143537 599907 143595 599913
rect 146021 599947 146079 599953
rect 146021 599913 146033 599947
rect 146067 599944 146079 599947
rect 157889 599947 157947 599953
rect 157889 599944 157901 599947
rect 146067 599916 157901 599944
rect 146067 599913 146079 599916
rect 146021 599907 146079 599913
rect 157889 599913 157901 599916
rect 157935 599913 157947 599947
rect 157889 599907 157947 599913
rect 157981 599947 158039 599953
rect 157981 599913 157993 599947
rect 158027 599913 158039 599947
rect 157981 599907 158039 599913
rect 188985 599947 189043 599953
rect 188985 599913 188997 599947
rect 189031 599913 189043 599947
rect 195793 599947 195851 599953
rect 195793 599944 195805 599947
rect 188985 599907 189043 599913
rect 195716 599916 195805 599944
rect 83016 599848 91784 599876
rect 95329 599879 95387 599885
rect 75638 599768 75644 599820
rect 75696 599808 75702 599820
rect 83016 599808 83044 599848
rect 95329 599845 95341 599879
rect 95375 599876 95387 599879
rect 113177 599879 113235 599885
rect 113177 599876 113189 599879
rect 95375 599848 113189 599876
rect 95375 599845 95387 599848
rect 95329 599839 95387 599845
rect 113177 599845 113189 599848
rect 113223 599845 113235 599879
rect 157996 599876 158024 599907
rect 160097 599879 160155 599885
rect 160097 599876 160109 599879
rect 157996 599848 160109 599876
rect 113177 599839 113235 599845
rect 160097 599845 160109 599848
rect 160143 599845 160155 599879
rect 189000 599876 189028 599907
rect 195716 599876 195744 599916
rect 195793 599913 195805 599916
rect 195839 599913 195851 599947
rect 195793 599907 195851 599913
rect 195885 599947 195943 599953
rect 195885 599913 195897 599947
rect 195931 599913 195943 599947
rect 202877 599947 202935 599953
rect 202877 599944 202889 599947
rect 195885 599907 195943 599913
rect 198016 599916 202889 599944
rect 189000 599848 195744 599876
rect 195900 599876 195928 599907
rect 198016 599876 198044 599916
rect 202877 599913 202889 599916
rect 202923 599913 202935 599947
rect 202877 599907 202935 599913
rect 212445 599947 212503 599953
rect 212445 599913 212457 599947
rect 212491 599913 212503 599947
rect 212445 599907 212503 599913
rect 215113 599947 215171 599953
rect 215113 599913 215125 599947
rect 215159 599913 215171 599947
rect 215113 599907 215171 599913
rect 215389 599947 215447 599953
rect 215389 599913 215401 599947
rect 215435 599944 215447 599947
rect 222197 599947 222255 599953
rect 222197 599944 222209 599947
rect 215435 599916 222209 599944
rect 215435 599913 215447 599916
rect 215389 599907 215447 599913
rect 222197 599913 222209 599916
rect 222243 599913 222255 599947
rect 222197 599907 222255 599913
rect 231765 599947 231823 599953
rect 231765 599913 231777 599947
rect 231811 599913 231823 599947
rect 231765 599907 231823 599913
rect 234433 599947 234491 599953
rect 234433 599913 234445 599947
rect 234479 599913 234491 599947
rect 234433 599907 234491 599913
rect 234709 599947 234767 599953
rect 234709 599913 234721 599947
rect 234755 599944 234767 599947
rect 241517 599947 241575 599953
rect 241517 599944 241529 599947
rect 234755 599916 241529 599944
rect 234755 599913 234767 599916
rect 234709 599907 234767 599913
rect 241517 599913 241529 599916
rect 241563 599913 241575 599947
rect 241517 599907 241575 599913
rect 251085 599947 251143 599953
rect 251085 599913 251097 599947
rect 251131 599913 251143 599947
rect 251085 599907 251143 599913
rect 253753 599947 253811 599953
rect 253753 599913 253765 599947
rect 253799 599913 253811 599947
rect 253753 599907 253811 599913
rect 254029 599947 254087 599953
rect 254029 599913 254041 599947
rect 254075 599944 254087 599947
rect 260837 599947 260895 599953
rect 260837 599944 260849 599947
rect 254075 599916 260849 599944
rect 254075 599913 254087 599916
rect 254029 599907 254087 599913
rect 260837 599913 260849 599916
rect 260883 599913 260895 599947
rect 260837 599907 260895 599913
rect 270405 599947 270463 599953
rect 270405 599913 270417 599947
rect 270451 599913 270463 599947
rect 270405 599907 270463 599913
rect 270497 599947 270555 599953
rect 270497 599913 270509 599947
rect 270543 599913 270555 599947
rect 270497 599907 270555 599913
rect 195900 599848 198044 599876
rect 212460 599876 212488 599907
rect 215128 599876 215156 599907
rect 212460 599848 215156 599876
rect 231780 599876 231808 599907
rect 234448 599876 234476 599907
rect 231780 599848 234476 599876
rect 251100 599876 251128 599907
rect 253768 599876 253796 599907
rect 251100 599848 253796 599876
rect 270420 599876 270448 599907
rect 270512 599876 270540 599907
rect 270420 599848 270540 599876
rect 160097 599839 160155 599845
rect 75696 599780 83044 599808
rect 75696 599768 75702 599780
rect 501690 599632 501696 599684
rect 501748 599672 501754 599684
rect 514018 599672 514024 599684
rect 501748 599644 514024 599672
rect 501748 599632 501754 599644
rect 514018 599632 514024 599644
rect 514076 599632 514082 599684
rect 48271 599576 51028 599604
rect 62776 599576 75224 599604
rect 501509 599607 501567 599613
rect 48271 599573 48283 599576
rect 48225 599567 48283 599573
rect 31757 599539 31815 599545
rect 31757 599536 31769 599539
rect 31680 599508 31769 599536
rect 31757 599505 31769 599508
rect 31803 599505 31815 599539
rect 51000 599536 51028 599576
rect 501509 599573 501521 599607
rect 501555 599604 501567 599607
rect 580350 599604 580356 599616
rect 501555 599576 580356 599604
rect 501555 599573 501567 599576
rect 501509 599567 501567 599573
rect 580350 599564 580356 599576
rect 580408 599564 580414 599616
rect 51077 599539 51135 599545
rect 51077 599536 51089 599539
rect 51000 599508 51089 599536
rect 31757 599499 31815 599505
rect 51077 599505 51089 599508
rect 51123 599505 51135 599539
rect 51077 599499 51135 599505
rect 9677 599471 9735 599477
rect 9677 599437 9689 599471
rect 9723 599468 9735 599471
rect 19245 599471 19303 599477
rect 19245 599468 19257 599471
rect 9723 599440 19257 599468
rect 9723 599437 9735 599440
rect 9677 599431 9735 599437
rect 19245 599437 19257 599440
rect 19291 599437 19303 599471
rect 19245 599431 19303 599437
rect 2682 599224 2688 599276
rect 2740 599264 2746 599276
rect 6181 599267 6239 599273
rect 6181 599264 6193 599267
rect 2740 599236 6193 599264
rect 2740 599224 2746 599236
rect 6181 599233 6193 599236
rect 6227 599233 6239 599267
rect 6181 599227 6239 599233
rect 64690 598952 64696 599004
rect 64748 598992 64754 599004
rect 78674 598992 78680 599004
rect 64748 598964 78680 598992
rect 64748 598952 64754 598964
rect 78674 598952 78680 598964
rect 78732 598952 78738 599004
rect 503990 598272 503996 598324
rect 504048 598312 504054 598324
rect 523126 598312 523132 598324
rect 504048 598284 523132 598312
rect 504048 598272 504054 598284
rect 523126 598272 523132 598284
rect 523184 598272 523190 598324
rect 502058 598204 502064 598256
rect 502116 598244 502122 598256
rect 534074 598244 534080 598256
rect 502116 598216 534080 598244
rect 502116 598204 502122 598216
rect 534074 598204 534080 598216
rect 534132 598204 534138 598256
rect 30282 596776 30288 596828
rect 30340 596816 30346 596828
rect 81434 596816 81440 596828
rect 30340 596788 81440 596816
rect 30340 596776 30346 596788
rect 81434 596776 81440 596788
rect 81492 596776 81498 596828
rect 502242 596776 502248 596828
rect 502300 596816 502306 596828
rect 512822 596816 512828 596828
rect 502300 596788 512828 596816
rect 502300 596776 502306 596788
rect 512822 596776 512828 596788
rect 512880 596776 512886 596828
rect 504358 596204 504364 596216
rect 504319 596176 504364 596204
rect 504358 596164 504364 596176
rect 504416 596164 504422 596216
rect 2866 594804 2872 594856
rect 2924 594844 2930 594856
rect 32398 594844 32404 594856
rect 2924 594816 32404 594844
rect 2924 594804 2930 594816
rect 32398 594804 32404 594816
rect 32456 594804 32462 594856
rect 20070 594056 20076 594108
rect 20128 594096 20134 594108
rect 78674 594096 78680 594108
rect 20128 594068 78680 594096
rect 20128 594056 20134 594068
rect 78674 594056 78680 594068
rect 78732 594056 78738 594108
rect 42702 592628 42708 592680
rect 42760 592668 42766 592680
rect 82906 592668 82912 592680
rect 42760 592640 82912 592668
rect 42760 592628 42766 592640
rect 82906 592628 82912 592640
rect 82964 592628 82970 592680
rect 60458 592016 60464 592068
rect 60516 592056 60522 592068
rect 78674 592056 78680 592068
rect 60516 592028 78680 592056
rect 60516 592016 60522 592028
rect 78674 592016 78680 592028
rect 78732 592016 78738 592068
rect 511258 592016 511264 592068
rect 511316 592056 511322 592068
rect 579890 592056 579896 592068
rect 511316 592028 579896 592056
rect 511316 592016 511322 592028
rect 579890 592016 579896 592028
rect 579948 592016 579954 592068
rect 507302 587120 507308 587172
rect 507360 587160 507366 587172
rect 523218 587160 523224 587172
rect 507360 587132 523224 587160
rect 507360 587120 507366 587132
rect 523218 587120 523224 587132
rect 523276 587120 523282 587172
rect 503898 586508 503904 586560
rect 503956 586548 503962 586560
rect 540238 586548 540244 586560
rect 503956 586520 540244 586548
rect 503956 586508 503962 586520
rect 540238 586508 540244 586520
rect 540296 586508 540302 586560
rect 72786 586440 72792 586492
rect 72844 586480 72850 586492
rect 73062 586480 73068 586492
rect 72844 586452 73068 586480
rect 72844 586440 72850 586452
rect 73062 586440 73068 586452
rect 73120 586440 73126 586492
rect 503898 582360 503904 582412
rect 503956 582400 503962 582412
rect 574094 582400 574100 582412
rect 503956 582372 574100 582400
rect 503956 582360 503962 582372
rect 574094 582360 574100 582372
rect 574152 582360 574158 582412
rect 560938 579640 560944 579692
rect 560996 579680 561002 579692
rect 580166 579680 580172 579692
rect 560996 579652 580172 579680
rect 560996 579640 561002 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 504358 578212 504364 578264
rect 504416 578252 504422 578264
rect 504450 578252 504456 578264
rect 504416 578224 504456 578252
rect 504416 578212 504422 578224
rect 504450 578212 504456 578224
rect 504508 578212 504514 578264
rect 75730 577124 75736 577176
rect 75788 577164 75794 577176
rect 78950 577164 78956 577176
rect 75788 577136 78956 577164
rect 75788 577124 75794 577136
rect 78950 577124 78956 577136
rect 79008 577124 79014 577176
rect 72786 576852 72792 576904
rect 72844 576892 72850 576904
rect 73062 576892 73068 576904
rect 72844 576864 73068 576892
rect 72844 576852 72850 576864
rect 73062 576852 73068 576864
rect 73120 576852 73126 576904
rect 501690 574064 501696 574116
rect 501748 574104 501754 574116
rect 501966 574104 501972 574116
rect 501748 574076 501972 574104
rect 501748 574064 501754 574076
rect 501966 574064 501972 574076
rect 502024 574064 502030 574116
rect 504358 572812 504364 572824
rect 504284 572784 504364 572812
rect 76926 572704 76932 572756
rect 76984 572744 76990 572756
rect 78766 572744 78772 572756
rect 76984 572716 78772 572744
rect 76984 572704 76990 572716
rect 78766 572704 78772 572716
rect 78824 572704 78830 572756
rect 504284 572688 504312 572784
rect 504358 572772 504364 572784
rect 504416 572772 504422 572824
rect 504266 572636 504272 572688
rect 504324 572636 504330 572688
rect 503898 571344 503904 571396
rect 503956 571384 503962 571396
rect 538858 571384 538864 571396
rect 503956 571356 538864 571384
rect 503956 571344 503962 571356
rect 538858 571344 538864 571356
rect 538916 571344 538922 571396
rect 50338 569916 50344 569968
rect 50396 569956 50402 569968
rect 78674 569956 78680 569968
rect 50396 569928 78680 569956
rect 50396 569916 50402 569928
rect 78674 569916 78680 569928
rect 78732 569916 78738 569968
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 25498 567236 25504 567248
rect 3476 567208 25504 567236
rect 3476 567196 3482 567208
rect 25498 567196 25504 567208
rect 25556 567196 25562 567248
rect 503898 567196 503904 567248
rect 503956 567236 503962 567248
rect 517974 567236 517980 567248
rect 503956 567208 517980 567236
rect 503956 567196 503962 567208
rect 517974 567196 517980 567208
rect 518032 567196 518038 567248
rect 46842 565836 46848 565888
rect 46900 565876 46906 565888
rect 78674 565876 78680 565888
rect 46900 565848 78680 565876
rect 46900 565836 46906 565848
rect 78674 565836 78680 565848
rect 78732 565836 78738 565888
rect 503898 564408 503904 564460
rect 503956 564448 503962 564460
rect 514846 564448 514852 564460
rect 503956 564420 514852 564448
rect 503956 564408 503962 564420
rect 514846 564408 514852 564420
rect 514904 564408 514910 564460
rect 504358 562912 504364 562964
rect 504416 562952 504422 562964
rect 504542 562952 504548 562964
rect 504416 562924 504548 562952
rect 504416 562912 504422 562924
rect 504542 562912 504548 562924
rect 504600 562912 504606 562964
rect 67358 561688 67364 561740
rect 67416 561728 67422 561740
rect 78674 561728 78680 561740
rect 67416 561700 78680 561728
rect 67416 561688 67422 561700
rect 78674 561688 78680 561700
rect 78732 561688 78738 561740
rect 503898 560260 503904 560312
rect 503956 560300 503962 560312
rect 520642 560300 520648 560312
rect 503956 560272 520648 560300
rect 503956 560260 503962 560272
rect 520642 560260 520648 560272
rect 520700 560260 520706 560312
rect 77018 558900 77024 558952
rect 77076 558940 77082 558952
rect 79594 558940 79600 558952
rect 77076 558912 79600 558940
rect 77076 558900 77082 558912
rect 79594 558900 79600 558912
rect 79652 558900 79658 558952
rect 512822 558900 512828 558952
rect 512880 558940 512886 558952
rect 513006 558940 513012 558952
rect 512880 558912 513012 558940
rect 512880 558900 512886 558912
rect 513006 558900 513012 558912
rect 513064 558900 513070 558952
rect 569310 556180 569316 556232
rect 569368 556220 569374 556232
rect 580166 556220 580172 556232
rect 569368 556192 580172 556220
rect 569368 556180 569374 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 501506 556112 501512 556164
rect 501564 556112 501570 556164
rect 501524 556028 501552 556112
rect 501506 555976 501512 556028
rect 501564 555976 501570 556028
rect 501690 554860 501696 554872
rect 501616 554832 501696 554860
rect 501616 554804 501644 554832
rect 501690 554820 501696 554832
rect 501748 554820 501754 554872
rect 63402 554752 63408 554804
rect 63460 554792 63466 554804
rect 78674 554792 78680 554804
rect 63460 554764 78680 554792
rect 63460 554752 63466 554764
rect 78674 554752 78680 554764
rect 78732 554752 78738 554804
rect 501598 554752 501604 554804
rect 501656 554752 501662 554804
rect 503898 554684 503904 554736
rect 503956 554724 503962 554736
rect 529198 554724 529204 554736
rect 503956 554696 529204 554724
rect 503956 554684 503962 554696
rect 529198 554684 529204 554696
rect 529256 554684 529262 554736
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 39298 552072 39304 552084
rect 3200 552044 39304 552072
rect 3200 552032 3206 552044
rect 39298 552032 39304 552044
rect 39356 552032 39362 552084
rect 503898 549244 503904 549296
rect 503956 549284 503962 549296
rect 518986 549284 518992 549296
rect 503956 549256 518992 549284
rect 503956 549244 503962 549256
rect 518986 549244 518992 549256
rect 519044 549244 519050 549296
rect 72786 547816 72792 547868
rect 72844 547856 72850 547868
rect 73062 547856 73068 547868
rect 72844 547828 73068 547856
rect 72844 547816 72850 547828
rect 73062 547816 73068 547828
rect 73120 547816 73126 547868
rect 504450 547136 504456 547188
rect 504508 547176 504514 547188
rect 536834 547176 536840 547188
rect 504508 547148 536840 547176
rect 504508 547136 504514 547148
rect 536834 547136 536840 547148
rect 536892 547136 536898 547188
rect 503898 545164 503904 545216
rect 503956 545204 503962 545216
rect 515030 545204 515036 545216
rect 503956 545176 515036 545204
rect 503956 545164 503962 545176
rect 515030 545164 515036 545176
rect 515088 545164 515094 545216
rect 512638 545096 512644 545148
rect 512696 545136 512702 545148
rect 579890 545136 579896 545148
rect 512696 545108 579896 545136
rect 512696 545096 512702 545108
rect 579890 545096 579896 545108
rect 579948 545096 579954 545148
rect 503898 541628 503904 541680
rect 503956 541668 503962 541680
rect 565078 541668 565084 541680
rect 503956 541640 565084 541668
rect 503956 541628 503962 541640
rect 565078 541628 565084 541640
rect 565136 541628 565142 541680
rect 3418 538228 3424 538280
rect 3476 538268 3482 538280
rect 43438 538268 43444 538280
rect 3476 538240 43444 538268
rect 3476 538228 3482 538240
rect 43438 538228 43444 538240
rect 43496 538228 43502 538280
rect 72786 538228 72792 538280
rect 72844 538268 72850 538280
rect 73062 538268 73068 538280
rect 72844 538240 73068 538268
rect 72844 538228 72850 538240
rect 73062 538228 73068 538240
rect 73120 538228 73126 538280
rect 503898 538228 503904 538280
rect 503956 538268 503962 538280
rect 521930 538268 521936 538280
rect 503956 538240 521936 538268
rect 503956 538228 503962 538240
rect 521930 538228 521936 538240
rect 521988 538228 521994 538280
rect 501598 536800 501604 536852
rect 501656 536800 501662 536852
rect 501616 536704 501644 536800
rect 501690 536704 501696 536716
rect 501616 536676 501696 536704
rect 501690 536664 501696 536676
rect 501748 536664 501754 536716
rect 504361 534191 504419 534197
rect 504361 534157 504373 534191
rect 504407 534188 504419 534191
rect 504450 534188 504456 534200
rect 504407 534160 504456 534188
rect 504407 534157 504419 534160
rect 504361 534151 504419 534157
rect 504450 534148 504456 534160
rect 504508 534148 504514 534200
rect 507210 534012 507216 534064
rect 507268 534052 507274 534064
rect 580166 534052 580172 534064
rect 507268 534024 580172 534052
rect 507268 534012 507274 534024
rect 580166 534012 580172 534024
rect 580224 534012 580230 534064
rect 504358 531332 504364 531344
rect 504319 531304 504364 531332
rect 504358 531292 504364 531304
rect 504416 531292 504422 531344
rect 512822 531292 512828 531344
rect 512880 531332 512886 531344
rect 513006 531332 513012 531344
rect 512880 531304 513012 531332
rect 512880 531292 512886 531304
rect 513006 531292 513012 531304
rect 513064 531292 513070 531344
rect 504450 531264 504456 531276
rect 504411 531236 504456 531264
rect 504450 531224 504456 531236
rect 504508 531224 504514 531276
rect 512822 529864 512828 529916
rect 512880 529904 512886 529916
rect 513006 529904 513012 529916
rect 512880 529876 513012 529904
rect 512880 529864 512886 529876
rect 513006 529864 513012 529876
rect 513064 529864 513070 529916
rect 76834 525784 76840 525836
rect 76892 525824 76898 525836
rect 78674 525824 78680 525836
rect 76892 525796 78680 525824
rect 76892 525784 76898 525796
rect 78674 525784 78680 525796
rect 78732 525784 78738 525836
rect 503898 524424 503904 524476
rect 503956 524464 503962 524476
rect 506474 524464 506480 524476
rect 503956 524436 506480 524464
rect 503956 524424 503962 524436
rect 506474 524424 506480 524436
rect 506532 524424 506538 524476
rect 504450 524328 504456 524340
rect 504411 524300 504456 524328
rect 504450 524288 504456 524300
rect 504508 524288 504514 524340
rect 503898 520276 503904 520328
rect 503956 520316 503962 520328
rect 520734 520316 520740 520328
rect 503956 520288 520740 520316
rect 503956 520276 503962 520288
rect 520734 520276 520740 520288
rect 520792 520276 520798 520328
rect 501601 520251 501659 520257
rect 501601 520217 501613 520251
rect 501647 520248 501659 520251
rect 501690 520248 501696 520260
rect 501647 520220 501696 520248
rect 501647 520217 501659 520220
rect 501601 520211 501659 520217
rect 501690 520208 501696 520220
rect 501748 520208 501754 520260
rect 75454 518916 75460 518968
rect 75512 518956 75518 518968
rect 78858 518956 78864 518968
rect 75512 518928 78864 518956
rect 75512 518916 75518 518928
rect 78858 518916 78864 518928
rect 78916 518916 78922 518968
rect 504358 514808 504364 514820
rect 504319 514780 504364 514808
rect 504358 514768 504364 514780
rect 504416 514768 504422 514820
rect 504358 512020 504364 512032
rect 504319 511992 504364 512020
rect 504358 511980 504364 511992
rect 504416 511980 504422 512032
rect 512822 511980 512828 512032
rect 512880 512020 512886 512032
rect 513006 512020 513012 512032
rect 512880 511992 513012 512020
rect 512880 511980 512886 511992
rect 513006 511980 513012 511992
rect 513064 511980 513070 512032
rect 63310 510620 63316 510672
rect 63368 510660 63374 510672
rect 78674 510660 78680 510672
rect 63368 510632 78680 510660
rect 63368 510620 63374 510632
rect 78674 510620 78680 510632
rect 78732 510620 78738 510672
rect 501598 510660 501604 510672
rect 501559 510632 501604 510660
rect 501598 510620 501604 510632
rect 501656 510620 501662 510672
rect 512822 510552 512828 510604
rect 512880 510592 512886 510604
rect 513006 510592 513012 510604
rect 512880 510564 513012 510592
rect 512880 510552 512886 510564
rect 513006 510552 513012 510564
rect 513064 510552 513070 510604
rect 565078 510552 565084 510604
rect 565136 510592 565142 510604
rect 580166 510592 580172 510604
rect 565136 510564 580172 510592
rect 565136 510552 565142 510564
rect 580166 510552 580172 510564
rect 580224 510552 580230 510604
rect 3142 509260 3148 509312
rect 3200 509300 3206 509312
rect 9122 509300 9128 509312
rect 3200 509272 9128 509300
rect 3200 509260 3206 509272
rect 9122 509260 9128 509272
rect 9180 509260 9186 509312
rect 64506 507832 64512 507884
rect 64564 507872 64570 507884
rect 78674 507872 78680 507884
rect 64564 507844 78680 507872
rect 64564 507832 64570 507844
rect 78674 507832 78680 507844
rect 78732 507832 78738 507884
rect 82906 507872 82912 507884
rect 82867 507844 82912 507872
rect 82906 507832 82912 507844
rect 82964 507832 82970 507884
rect 501598 507804 501604 507816
rect 501559 507776 501604 507804
rect 501598 507764 501604 507776
rect 501656 507764 501662 507816
rect 504358 505112 504364 505164
rect 504416 505112 504422 505164
rect 504376 505016 504404 505112
rect 504450 505016 504456 505028
rect 504376 504988 504456 505016
rect 504450 504976 504456 504988
rect 504508 504976 504514 505028
rect 66070 503684 66076 503736
rect 66128 503724 66134 503736
rect 78674 503724 78680 503736
rect 66128 503696 78680 503724
rect 66128 503684 66134 503696
rect 78674 503684 78680 503696
rect 78732 503684 78738 503736
rect 79229 501755 79287 501761
rect 79229 501721 79241 501755
rect 79275 501752 79287 501755
rect 82906 501752 82912 501764
rect 79275 501724 82912 501752
rect 79275 501721 79287 501724
rect 79229 501715 79287 501721
rect 82906 501712 82912 501724
rect 82964 501712 82970 501764
rect 82906 501616 82912 501628
rect 82867 501588 82912 501616
rect 82906 501576 82912 501588
rect 82964 501576 82970 501628
rect 77110 500012 77116 500064
rect 77168 500052 77174 500064
rect 79042 500052 79048 500064
rect 77168 500024 79048 500052
rect 77168 500012 77174 500024
rect 79042 500012 79048 500024
rect 79100 500012 79106 500064
rect 508498 499468 508504 499520
rect 508556 499508 508562 499520
rect 580166 499508 580172 499520
rect 508556 499480 580172 499508
rect 508556 499468 508562 499480
rect 580166 499468 580172 499480
rect 580224 499468 580230 499520
rect 501601 498219 501659 498225
rect 501601 498185 501613 498219
rect 501647 498216 501659 498219
rect 501690 498216 501696 498228
rect 501647 498188 501696 498216
rect 501647 498185 501659 498188
rect 501601 498179 501659 498185
rect 501690 498176 501696 498188
rect 501748 498176 501754 498228
rect 503898 498176 503904 498228
rect 503956 498216 503962 498228
rect 507946 498216 507952 498228
rect 503956 498188 507952 498216
rect 503956 498176 503962 498188
rect 507946 498176 507952 498188
rect 508004 498176 508010 498228
rect 504174 497496 504180 497548
rect 504232 497536 504238 497548
rect 504358 497536 504364 497548
rect 504232 497508 504364 497536
rect 504232 497496 504238 497508
rect 504358 497496 504364 497508
rect 504416 497496 504422 497548
rect 61654 496816 61660 496868
rect 61712 496856 61718 496868
rect 78674 496856 78680 496868
rect 61712 496828 78680 496856
rect 61712 496816 61718 496828
rect 78674 496816 78680 496828
rect 78732 496816 78738 496868
rect 3418 496748 3424 496800
rect 3476 496788 3482 496800
rect 79229 496791 79287 496797
rect 79229 496788 79241 496791
rect 3476 496760 79241 496788
rect 3476 496748 3482 496760
rect 79229 496757 79241 496760
rect 79275 496757 79287 496791
rect 79229 496751 79287 496757
rect 503898 494028 503904 494080
rect 503956 494068 503962 494080
rect 513650 494068 513656 494080
rect 503956 494040 513656 494068
rect 503956 494028 503962 494040
rect 513650 494028 513656 494040
rect 513708 494028 513714 494080
rect 512822 491280 512828 491292
rect 512783 491252 512828 491280
rect 512822 491240 512828 491252
rect 512880 491240 512886 491292
rect 72786 489812 72792 489864
rect 72844 489852 72850 489864
rect 73062 489852 73068 489864
rect 72844 489824 73068 489852
rect 72844 489812 72850 489824
rect 73062 489812 73068 489824
rect 73120 489812 73126 489864
rect 503898 487160 503904 487212
rect 503956 487200 503962 487212
rect 571978 487200 571984 487212
rect 503956 487172 571984 487200
rect 503956 487160 503962 487172
rect 571978 487160 571984 487172
rect 572036 487160 572042 487212
rect 65978 485800 65984 485852
rect 66036 485840 66042 485852
rect 78674 485840 78680 485852
rect 66036 485812 78680 485840
rect 66036 485800 66042 485812
rect 78674 485800 78680 485812
rect 78732 485800 78738 485852
rect 504358 485800 504364 485852
rect 504416 485800 504422 485852
rect 567838 485800 567844 485852
rect 567896 485840 567902 485852
rect 580166 485840 580172 485852
rect 567896 485812 580172 485840
rect 567896 485800 567902 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 504376 485704 504404 485800
rect 504450 485704 504456 485716
rect 504376 485676 504456 485704
rect 504450 485664 504456 485676
rect 504508 485664 504514 485716
rect 503898 483012 503904 483064
rect 503956 483052 503962 483064
rect 522022 483052 522028 483064
rect 503956 483024 522028 483052
rect 503956 483012 503962 483024
rect 522022 483012 522028 483024
rect 522080 483012 522086 483064
rect 504450 482944 504456 482996
rect 504508 482984 504514 482996
rect 504634 482984 504640 482996
rect 504508 482956 504640 482984
rect 504508 482944 504514 482956
rect 504634 482944 504640 482956
rect 504692 482944 504698 482996
rect 512822 481692 512828 481704
rect 512783 481664 512828 481692
rect 512822 481652 512828 481664
rect 512880 481652 512886 481704
rect 3786 481584 3792 481636
rect 3844 481624 3850 481636
rect 39390 481624 39396 481636
rect 3844 481596 39396 481624
rect 3844 481584 3850 481596
rect 39390 481584 39396 481596
rect 39448 481584 39454 481636
rect 72786 480224 72792 480276
rect 72844 480264 72850 480276
rect 73062 480264 73068 480276
rect 72844 480236 73068 480264
rect 72844 480224 72850 480236
rect 73062 480224 73068 480236
rect 73120 480224 73126 480276
rect 501598 480224 501604 480276
rect 501656 480264 501662 480276
rect 501690 480264 501696 480276
rect 501656 480236 501696 480264
rect 501656 480224 501662 480236
rect 501690 480224 501696 480236
rect 501748 480224 501754 480276
rect 61562 478864 61568 478916
rect 61620 478904 61626 478916
rect 78674 478904 78680 478916
rect 61620 478876 78680 478904
rect 61620 478864 61626 478876
rect 78674 478864 78680 478876
rect 78732 478864 78738 478916
rect 503898 476076 503904 476128
rect 503956 476116 503962 476128
rect 516502 476116 516508 476128
rect 503956 476088 516508 476116
rect 503956 476076 503962 476088
rect 516502 476076 516508 476088
rect 516560 476076 516566 476128
rect 82909 474963 82967 474969
rect 82909 474929 82921 474963
rect 82955 474960 82967 474963
rect 82998 474960 83004 474972
rect 82955 474932 83004 474960
rect 82955 474929 82967 474932
rect 82909 474923 82967 474929
rect 82998 474920 83004 474932
rect 83056 474920 83062 474972
rect 503898 473356 503904 473408
rect 503956 473396 503962 473408
rect 523310 473396 523316 473408
rect 503956 473368 523316 473396
rect 503956 473356 503962 473368
rect 523310 473356 523316 473368
rect 523368 473356 523374 473408
rect 48958 471928 48964 471980
rect 49016 471968 49022 471980
rect 78674 471968 78680 471980
rect 49016 471940 78680 471968
rect 49016 471928 49022 471940
rect 78674 471928 78680 471940
rect 78732 471928 78738 471980
rect 512822 471968 512828 471980
rect 512783 471940 512828 471968
rect 512822 471928 512828 471940
rect 512880 471928 512886 471980
rect 82909 469251 82967 469257
rect 82909 469217 82921 469251
rect 82955 469248 82967 469251
rect 82998 469248 83004 469260
rect 82955 469220 83004 469248
rect 82955 469217 82967 469220
rect 82909 469211 82967 469217
rect 82998 469208 83004 469220
rect 83056 469208 83062 469260
rect 503898 469208 503904 469260
rect 503956 469248 503962 469260
rect 510798 469248 510804 469260
rect 503956 469220 510804 469248
rect 503956 469208 503962 469220
rect 510798 469208 510804 469220
rect 510856 469208 510862 469260
rect 501598 467780 501604 467832
rect 501656 467820 501662 467832
rect 501690 467820 501696 467832
rect 501656 467792 501696 467820
rect 501656 467780 501662 467792
rect 501690 467780 501696 467792
rect 501748 467780 501754 467832
rect 504358 466420 504364 466472
rect 504416 466420 504422 466472
rect 504376 466392 504404 466420
rect 504450 466392 504456 466404
rect 504376 466364 504456 466392
rect 504450 466352 504456 466364
rect 504508 466352 504514 466404
rect 504174 463632 504180 463684
rect 504232 463672 504238 463684
rect 504450 463672 504456 463684
rect 504232 463644 504456 463672
rect 504232 463632 504238 463644
rect 504450 463632 504456 463644
rect 504508 463632 504514 463684
rect 512822 462380 512828 462392
rect 512783 462352 512828 462380
rect 512822 462340 512828 462352
rect 512880 462340 512886 462392
rect 565078 462340 565084 462392
rect 565136 462380 565142 462392
rect 580166 462380 580172 462392
rect 565136 462352 580172 462380
rect 565136 462340 565142 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 503898 461524 503904 461576
rect 503956 461564 503962 461576
rect 508038 461564 508044 461576
rect 503956 461536 508044 461564
rect 503956 461524 503962 461536
rect 508038 461524 508044 461536
rect 508096 461524 508102 461576
rect 68646 459552 68652 459604
rect 68704 459592 68710 459604
rect 78674 459592 78680 459604
rect 68704 459564 78680 459592
rect 68704 459552 68710 459564
rect 78674 459552 78680 459564
rect 78732 459552 78738 459604
rect 75362 456764 75368 456816
rect 75420 456804 75426 456816
rect 78674 456804 78680 456816
rect 75420 456776 78680 456804
rect 75420 456764 75426 456776
rect 78674 456764 78680 456776
rect 78732 456764 78738 456816
rect 509878 452548 509884 452600
rect 509936 452588 509942 452600
rect 580166 452588 580172 452600
rect 509936 452560 580172 452588
rect 509936 452548 509942 452560
rect 580166 452548 580172 452560
rect 580224 452548 580230 452600
rect 512822 452520 512828 452532
rect 512783 452492 512828 452520
rect 512822 452480 512828 452492
rect 512880 452480 512886 452532
rect 72786 451188 72792 451240
rect 72844 451228 72850 451240
rect 73062 451228 73068 451240
rect 72844 451200 73068 451228
rect 72844 451188 72850 451200
rect 73062 451188 73068 451200
rect 73120 451188 73126 451240
rect 501598 449896 501604 449948
rect 501656 449936 501662 449948
rect 501690 449936 501696 449948
rect 501656 449908 501696 449936
rect 501656 449896 501662 449908
rect 501690 449896 501696 449908
rect 501748 449896 501754 449948
rect 74074 448536 74080 448588
rect 74132 448576 74138 448588
rect 78674 448576 78680 448588
rect 74132 448548 78680 448576
rect 74132 448536 74138 448548
rect 78674 448536 78680 448548
rect 78732 448536 78738 448588
rect 82906 448576 82912 448588
rect 82867 448548 82912 448576
rect 82906 448536 82912 448548
rect 82964 448536 82970 448588
rect 501598 448468 501604 448520
rect 501656 448508 501662 448520
rect 501690 448508 501696 448520
rect 501656 448480 501696 448508
rect 501656 448468 501662 448480
rect 501690 448468 501696 448480
rect 501748 448468 501754 448520
rect 503898 447108 503904 447160
rect 503956 447148 503962 447160
rect 506566 447148 506572 447160
rect 503956 447120 506572 447148
rect 503956 447108 503962 447120
rect 506566 447108 506572 447120
rect 506624 447108 506630 447160
rect 60366 445748 60372 445800
rect 60424 445788 60430 445800
rect 78674 445788 78680 445800
rect 60424 445760 78680 445788
rect 60424 445748 60430 445760
rect 78674 445748 78680 445760
rect 78732 445748 78738 445800
rect 82817 444363 82875 444369
rect 82817 444329 82829 444363
rect 82863 444360 82875 444363
rect 82906 444360 82912 444372
rect 82863 444332 82912 444360
rect 82863 444329 82875 444332
rect 82817 444323 82875 444329
rect 82906 444320 82912 444332
rect 82964 444320 82970 444372
rect 504361 444363 504419 444369
rect 504361 444329 504373 444363
rect 504407 444360 504419 444363
rect 504450 444360 504456 444372
rect 504407 444332 504456 444360
rect 504407 444329 504419 444332
rect 504361 444323 504419 444329
rect 504450 444320 504456 444332
rect 504508 444320 504514 444372
rect 503898 442960 503904 443012
rect 503956 443000 503962 443012
rect 509602 443000 509608 443012
rect 503956 442972 509608 443000
rect 503956 442960 503962 442972
rect 509602 442960 509608 442972
rect 509660 442960 509666 443012
rect 512822 443000 512828 443012
rect 512783 442972 512828 443000
rect 512822 442960 512828 442972
rect 512880 442960 512886 443012
rect 82817 441983 82875 441989
rect 82817 441949 82829 441983
rect 82863 441980 82875 441983
rect 82906 441980 82912 441992
rect 82863 441952 82912 441980
rect 82863 441949 82875 441952
rect 82817 441943 82875 441949
rect 82906 441940 82912 441952
rect 82964 441940 82970 441992
rect 72786 441668 72792 441720
rect 72844 441708 72850 441720
rect 73062 441708 73068 441720
rect 72844 441680 73068 441708
rect 72844 441668 72850 441680
rect 73062 441668 73068 441680
rect 73120 441668 73126 441720
rect 82906 441708 82912 441720
rect 82867 441680 82912 441708
rect 82906 441668 82912 441680
rect 82964 441668 82970 441720
rect 64414 441600 64420 441652
rect 64472 441640 64478 441652
rect 78674 441640 78680 441652
rect 64472 441612 78680 441640
rect 64472 441600 64478 441612
rect 78674 441600 78680 441612
rect 78732 441600 78738 441652
rect 503898 440240 503904 440292
rect 503956 440280 503962 440292
rect 509510 440280 509516 440292
rect 503956 440252 509516 440280
rect 503956 440240 503962 440252
rect 509510 440240 509516 440252
rect 509568 440240 509574 440292
rect 82814 440172 82820 440224
rect 82872 440212 82878 440224
rect 82906 440212 82912 440224
rect 82872 440184 82912 440212
rect 82872 440172 82878 440184
rect 82906 440172 82912 440184
rect 82964 440172 82970 440224
rect 514110 440172 514116 440224
rect 514168 440212 514174 440224
rect 579614 440212 579620 440224
rect 514168 440184 579620 440212
rect 514168 440172 514174 440184
rect 579614 440172 579620 440184
rect 579672 440172 579678 440224
rect 503898 436092 503904 436144
rect 503956 436132 503962 436144
rect 519078 436132 519084 436144
rect 503956 436104 519084 436132
rect 503956 436092 503962 436104
rect 519078 436092 519084 436104
rect 519136 436092 519142 436144
rect 504358 434772 504364 434784
rect 504319 434744 504364 434772
rect 504358 434732 504364 434744
rect 504416 434732 504422 434784
rect 512822 433276 512828 433288
rect 512783 433248 512828 433276
rect 512822 433236 512828 433248
rect 512880 433236 512886 433288
rect 503898 432488 503904 432540
rect 503956 432528 503962 432540
rect 506750 432528 506756 432540
rect 503956 432500 506756 432528
rect 503956 432488 503962 432500
rect 506750 432488 506756 432500
rect 506808 432488 506814 432540
rect 72786 431876 72792 431928
rect 72844 431916 72850 431928
rect 73062 431916 73068 431928
rect 72844 431888 73068 431916
rect 72844 431876 72850 431888
rect 73062 431876 73068 431888
rect 73120 431876 73126 431928
rect 59078 430584 59084 430636
rect 59136 430624 59142 430636
rect 78674 430624 78680 430636
rect 59136 430596 78680 430624
rect 59136 430584 59142 430596
rect 78674 430584 78680 430596
rect 78732 430584 78738 430636
rect 82814 430516 82820 430568
rect 82872 430556 82878 430568
rect 82998 430556 83004 430568
rect 82872 430528 83004 430556
rect 82872 430516 82878 430528
rect 82998 430516 83004 430528
rect 83056 430516 83062 430568
rect 503898 429156 503904 429208
rect 503956 429196 503962 429208
rect 522114 429196 522120 429208
rect 503956 429168 522120 429196
rect 503956 429156 503962 429168
rect 522114 429156 522120 429168
rect 522172 429156 522178 429208
rect 19978 427796 19984 427848
rect 20036 427836 20042 427848
rect 78674 427836 78680 427848
rect 20036 427808 78680 427836
rect 20036 427796 20042 427808
rect 78674 427796 78680 427808
rect 78732 427796 78738 427848
rect 504358 427796 504364 427848
rect 504416 427796 504422 427848
rect 504376 427768 504404 427796
rect 504450 427768 504456 427780
rect 504376 427740 504456 427768
rect 504450 427728 504456 427740
rect 504508 427728 504514 427780
rect 503898 425076 503904 425128
rect 503956 425116 503962 425128
rect 509418 425116 509424 425128
rect 503956 425088 509424 425116
rect 503956 425076 503962 425088
rect 509418 425076 509424 425088
rect 509476 425076 509482 425128
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 69750 425048 69756 425060
rect 3292 425020 69756 425048
rect 3292 425008 3298 425020
rect 69750 425008 69756 425020
rect 69808 425008 69814 425060
rect 504361 425051 504419 425057
rect 504361 425017 504373 425051
rect 504407 425048 504419 425051
rect 504450 425048 504456 425060
rect 504407 425020 504456 425048
rect 504407 425017 504419 425020
rect 504361 425011 504419 425017
rect 504450 425008 504456 425020
rect 504508 425008 504514 425060
rect 501966 423648 501972 423700
rect 502024 423688 502030 423700
rect 502058 423688 502064 423700
rect 502024 423660 502064 423688
rect 502024 423648 502030 423660
rect 502058 423648 502064 423660
rect 502116 423648 502122 423700
rect 512822 423688 512828 423700
rect 512783 423660 512828 423688
rect 512822 423648 512828 423660
rect 512880 423648 512886 423700
rect 72786 422288 72792 422340
rect 72844 422328 72850 422340
rect 73062 422328 73068 422340
rect 72844 422300 73068 422328
rect 72844 422288 72850 422300
rect 73062 422288 73068 422300
rect 73120 422288 73126 422340
rect 503898 420928 503904 420980
rect 503956 420968 503962 420980
rect 506658 420968 506664 420980
rect 503956 420940 506664 420968
rect 503956 420928 503962 420940
rect 506658 420928 506664 420940
rect 506716 420928 506722 420980
rect 46198 419500 46204 419552
rect 46256 419540 46262 419552
rect 78674 419540 78680 419552
rect 46256 419512 78680 419540
rect 46256 419500 46262 419512
rect 78674 419500 78680 419512
rect 78732 419500 78738 419552
rect 3418 417392 3424 417444
rect 3476 417432 3482 417444
rect 69750 417432 69756 417444
rect 3476 417404 69756 417432
rect 3476 417392 3482 417404
rect 69750 417392 69756 417404
rect 69808 417392 69814 417444
rect 76742 416780 76748 416832
rect 76800 416820 76806 416832
rect 78674 416820 78680 416832
rect 76800 416792 78680 416820
rect 76800 416780 76806 416792
rect 78674 416780 78680 416792
rect 78732 416780 78738 416832
rect 504358 415460 504364 415472
rect 504319 415432 504364 415460
rect 504358 415420 504364 415432
rect 504416 415420 504422 415472
rect 512822 413964 512828 413976
rect 512783 413936 512828 413964
rect 512822 413924 512828 413936
rect 512880 413924 512886 413976
rect 65886 412632 65892 412684
rect 65944 412672 65950 412684
rect 78674 412672 78680 412684
rect 65944 412644 78680 412672
rect 65944 412632 65950 412644
rect 78674 412632 78680 412644
rect 78732 412632 78738 412684
rect 72786 412564 72792 412616
rect 72844 412604 72850 412616
rect 73062 412604 73068 412616
rect 72844 412576 73068 412604
rect 72844 412564 72850 412576
rect 73062 412564 73068 412576
rect 73120 412564 73126 412616
rect 501598 411272 501604 411324
rect 501656 411312 501662 411324
rect 501782 411312 501788 411324
rect 501656 411284 501788 411312
rect 501656 411272 501662 411284
rect 501782 411272 501788 411284
rect 501840 411272 501846 411324
rect 504358 408484 504364 408536
rect 504416 408484 504422 408536
rect 504376 408388 504404 408484
rect 504450 408388 504456 408400
rect 504376 408360 504456 408388
rect 504450 408348 504456 408360
rect 504508 408348 504514 408400
rect 503898 407124 503904 407176
rect 503956 407164 503962 407176
rect 508222 407164 508228 407176
rect 503956 407136 508228 407164
rect 503956 407124 503962 407136
rect 508222 407124 508228 407136
rect 508280 407124 508286 407176
rect 63218 405696 63224 405748
rect 63276 405736 63282 405748
rect 78674 405736 78680 405748
rect 63276 405708 78680 405736
rect 63276 405696 63282 405708
rect 78674 405696 78680 405708
rect 78732 405696 78738 405748
rect 512822 404376 512828 404388
rect 512783 404348 512828 404376
rect 512822 404336 512828 404348
rect 512880 404336 512886 404388
rect 516778 404336 516784 404388
rect 516836 404376 516842 404388
rect 580166 404376 580172 404388
rect 516836 404348 580172 404376
rect 516836 404336 516842 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 72786 402976 72792 403028
rect 72844 403016 72850 403028
rect 73062 403016 73068 403028
rect 72844 402988 73068 403016
rect 72844 402976 72850 402988
rect 73062 402976 73068 402988
rect 73120 402976 73126 403028
rect 503898 402976 503904 403028
rect 503956 403016 503962 403028
rect 513742 403016 513748 403028
rect 503956 402988 513748 403016
rect 503956 402976 503962 402988
rect 513742 402976 513748 402988
rect 513800 402976 513806 403028
rect 64322 401616 64328 401668
rect 64380 401656 64386 401668
rect 78674 401656 78680 401668
rect 64380 401628 78680 401656
rect 64380 401616 64386 401628
rect 78674 401616 78680 401628
rect 78732 401616 78738 401668
rect 504450 400868 504456 400920
rect 504508 400908 504514 400920
rect 504634 400908 504640 400920
rect 504508 400880 504640 400908
rect 504508 400868 504514 400880
rect 504634 400868 504640 400880
rect 504692 400868 504698 400920
rect 503898 398828 503904 398880
rect 503956 398868 503962 398880
rect 520826 398868 520832 398880
rect 503956 398840 520832 398868
rect 503956 398828 503962 398840
rect 520826 398828 520832 398840
rect 520884 398828 520890 398880
rect 33778 397468 33784 397520
rect 33836 397508 33842 397520
rect 78674 397508 78680 397520
rect 33836 397480 78680 397508
rect 33836 397468 33842 397480
rect 78674 397468 78680 397480
rect 78732 397468 78738 397520
rect 3326 394680 3332 394732
rect 3384 394720 3390 394732
rect 69842 394720 69848 394732
rect 3384 394692 69848 394720
rect 3384 394680 3390 394692
rect 69842 394680 69848 394692
rect 69900 394680 69906 394732
rect 512822 394652 512828 394664
rect 512783 394624 512828 394652
rect 512822 394612 512828 394624
rect 512880 394612 512886 394664
rect 72786 393252 72792 393304
rect 72844 393292 72850 393304
rect 73062 393292 73068 393304
rect 72844 393264 73068 393292
rect 72844 393252 72850 393264
rect 73062 393252 73068 393264
rect 73120 393252 73126 393304
rect 504358 393252 504364 393304
rect 504416 393292 504422 393304
rect 504450 393292 504456 393304
rect 504416 393264 504456 393292
rect 504416 393252 504422 393264
rect 504450 393252 504456 393264
rect 504508 393252 504514 393304
rect 507118 393252 507124 393304
rect 507176 393292 507182 393304
rect 580166 393292 580172 393304
rect 507176 393264 580172 393292
rect 507176 393252 507182 393264
rect 580166 393252 580172 393264
rect 580224 393252 580230 393304
rect 501690 391892 501696 391944
rect 501748 391932 501754 391944
rect 501782 391932 501788 391944
rect 501748 391904 501788 391932
rect 501748 391892 501754 391904
rect 501782 391892 501788 391904
rect 501840 391892 501846 391944
rect 503898 389172 503904 389224
rect 503956 389212 503962 389224
rect 573450 389212 573456 389224
rect 503956 389184 573456 389212
rect 503956 389172 503962 389184
rect 573450 389172 573456 389184
rect 573508 389172 573514 389224
rect 63126 386384 63132 386436
rect 63184 386424 63190 386436
rect 78674 386424 78680 386436
rect 63184 386396 78680 386424
rect 63184 386384 63190 386396
rect 78674 386384 78680 386396
rect 78732 386384 78738 386436
rect 82817 386291 82875 386297
rect 82817 386257 82829 386291
rect 82863 386288 82875 386291
rect 82906 386288 82912 386300
rect 82863 386260 82912 386288
rect 82863 386257 82875 386260
rect 82817 386251 82875 386257
rect 82906 386248 82912 386260
rect 82964 386248 82970 386300
rect 512822 385132 512828 385144
rect 512783 385104 512828 385132
rect 512822 385092 512828 385104
rect 512880 385092 512886 385144
rect 503898 385024 503904 385076
rect 503956 385064 503962 385076
rect 549898 385064 549904 385076
rect 503956 385036 549904 385064
rect 503956 385024 503962 385036
rect 549898 385024 549904 385036
rect 549956 385024 549962 385076
rect 72786 383732 72792 383784
rect 72844 383772 72850 383784
rect 73062 383772 73068 383784
rect 72844 383744 73068 383772
rect 72844 383732 72850 383744
rect 73062 383732 73068 383744
rect 73120 383732 73126 383784
rect 65794 383664 65800 383716
rect 65852 383704 65858 383716
rect 78674 383704 78680 383716
rect 65852 383676 78680 383704
rect 65852 383664 65858 383676
rect 78674 383664 78680 383676
rect 78732 383664 78738 383716
rect 502978 382916 502984 382968
rect 503036 382956 503042 382968
rect 523402 382956 523408 382968
rect 503036 382928 523408 382956
rect 503036 382916 503042 382928
rect 523402 382916 523408 382928
rect 523460 382916 523466 382968
rect 503898 380876 503904 380928
rect 503956 380916 503962 380928
rect 519170 380916 519176 380928
rect 503956 380888 519176 380916
rect 503956 380876 503962 380888
rect 519170 380876 519176 380888
rect 519228 380876 519234 380928
rect 3418 379516 3424 379568
rect 3476 379556 3482 379568
rect 13170 379556 13176 379568
rect 3476 379528 13176 379556
rect 3476 379516 3482 379528
rect 13170 379516 13176 379528
rect 13228 379516 13234 379568
rect 503898 378156 503904 378208
rect 503956 378196 503962 378208
rect 506934 378196 506940 378208
rect 503956 378168 506940 378196
rect 503956 378156 503962 378168
rect 506934 378156 506940 378168
rect 506992 378156 506998 378208
rect 501690 376660 501696 376712
rect 501748 376700 501754 376712
rect 501782 376700 501788 376712
rect 501748 376672 501788 376700
rect 501748 376660 501754 376672
rect 501782 376660 501788 376672
rect 501840 376660 501846 376712
rect 503898 375300 503904 375352
rect 503956 375340 503962 375352
rect 522298 375340 522304 375352
rect 503956 375312 522304 375340
rect 503956 375300 503962 375312
rect 522298 375300 522304 375312
rect 522356 375300 522362 375352
rect 512822 375272 512828 375284
rect 512783 375244 512828 375272
rect 512822 375232 512828 375244
rect 512880 375232 512886 375284
rect 82814 374796 82820 374808
rect 82775 374768 82820 374796
rect 82814 374756 82820 374768
rect 82872 374756 82878 374808
rect 72786 373940 72792 373992
rect 72844 373980 72850 373992
rect 73062 373980 73068 373992
rect 72844 373952 73068 373980
rect 72844 373940 72850 373952
rect 73062 373940 73068 373952
rect 73120 373940 73126 373992
rect 49602 368500 49608 368552
rect 49660 368540 49666 368552
rect 78674 368540 78680 368552
rect 49660 368512 78680 368540
rect 49660 368500 49666 368512
rect 78674 368500 78680 368512
rect 78732 368500 78738 368552
rect 514110 368500 514116 368552
rect 514168 368540 514174 368552
rect 580166 368540 580172 368552
rect 514168 368512 580172 368540
rect 514168 368500 514174 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 503990 367072 503996 367124
rect 504048 367112 504054 367124
rect 506842 367112 506848 367124
rect 504048 367084 506848 367112
rect 504048 367072 504054 367084
rect 506842 367072 506848 367084
rect 506900 367072 506906 367124
rect 504450 367044 504456 367056
rect 504376 367016 504456 367044
rect 504376 366988 504404 367016
rect 504450 367004 504456 367016
rect 504508 367004 504514 367056
rect 504358 366936 504364 366988
rect 504416 366936 504422 366988
rect 512822 365752 512828 365764
rect 512783 365724 512828 365752
rect 512822 365712 512828 365724
rect 512880 365712 512886 365764
rect 72786 364352 72792 364404
rect 72844 364392 72850 364404
rect 73062 364392 73068 364404
rect 72844 364364 73068 364392
rect 72844 364352 72850 364364
rect 73062 364352 73068 364364
rect 73120 364352 73126 364404
rect 503990 362924 503996 362976
rect 504048 362964 504054 362976
rect 516594 362964 516600 362976
rect 504048 362936 516600 362964
rect 504048 362924 504054 362936
rect 516594 362924 516600 362936
rect 516652 362924 516658 362976
rect 37918 361564 37924 361616
rect 37976 361604 37982 361616
rect 78674 361604 78680 361616
rect 37976 361576 78680 361604
rect 37976 361564 37982 361576
rect 78674 361564 78680 361576
rect 78732 361564 78738 361616
rect 501690 358776 501696 358828
rect 501748 358816 501754 358828
rect 501782 358816 501788 358828
rect 501748 358788 501788 358816
rect 501748 358776 501754 358788
rect 501782 358776 501788 358788
rect 501840 358776 501846 358828
rect 512822 357552 512828 357604
rect 512880 357552 512886 357604
rect 512840 357468 512868 357552
rect 75270 357416 75276 357468
rect 75328 357456 75334 357468
rect 78674 357456 78680 357468
rect 75328 357428 78680 357456
rect 75328 357416 75334 357428
rect 78674 357416 78680 357428
rect 78732 357416 78738 357468
rect 512822 357416 512828 357468
rect 512880 357416 512886 357468
rect 569218 357416 569224 357468
rect 569276 357456 569282 357468
rect 580166 357456 580172 357468
rect 569276 357428 580172 357456
rect 569276 357416 569282 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 501598 357348 501604 357400
rect 501656 357388 501662 357400
rect 501690 357388 501696 357400
rect 501656 357360 501696 357388
rect 501656 357348 501662 357360
rect 501690 357348 501696 357360
rect 501748 357348 501754 357400
rect 512822 356028 512828 356040
rect 512783 356000 512828 356028
rect 512822 355988 512828 356000
rect 512880 355988 512886 356040
rect 505738 355308 505744 355360
rect 505796 355348 505802 355360
rect 519630 355348 519636 355360
rect 505796 355320 519636 355348
rect 505796 355308 505802 355320
rect 519630 355308 519636 355320
rect 519688 355308 519694 355360
rect 13170 351840 13176 351892
rect 13228 351880 13234 351892
rect 78674 351880 78680 351892
rect 13228 351852 78680 351880
rect 13228 351840 13234 351852
rect 78674 351840 78680 351852
rect 78732 351840 78738 351892
rect 15930 346400 15936 346452
rect 15988 346440 15994 346452
rect 78674 346440 78680 346452
rect 15988 346412 78680 346440
rect 15988 346400 15994 346412
rect 78674 346400 78680 346412
rect 78732 346400 78738 346452
rect 512822 346440 512828 346452
rect 512783 346412 512828 346440
rect 512822 346400 512828 346412
rect 512880 346400 512886 346452
rect 504082 345040 504088 345092
rect 504140 345080 504146 345092
rect 513834 345080 513840 345092
rect 504140 345052 513840 345080
rect 504140 345040 504146 345052
rect 513834 345040 513840 345052
rect 513892 345040 513898 345092
rect 82906 342496 82912 342508
rect 82867 342468 82912 342496
rect 82906 342456 82912 342468
rect 82964 342456 82970 342508
rect 504082 340892 504088 340944
rect 504140 340932 504146 340944
rect 527818 340932 527824 340944
rect 504140 340904 527824 340932
rect 504140 340892 504146 340904
rect 527818 340892 527824 340904
rect 527876 340892 527882 340944
rect 501598 339396 501604 339448
rect 501656 339436 501662 339448
rect 501690 339436 501696 339448
rect 501656 339408 501696 339436
rect 501656 339396 501662 339408
rect 501690 339396 501696 339408
rect 501748 339396 501754 339448
rect 504082 338104 504088 338156
rect 504140 338144 504146 338156
rect 519262 338144 519268 338156
rect 504140 338116 519268 338144
rect 504140 338104 504146 338116
rect 519262 338104 519268 338116
rect 519320 338104 519326 338156
rect 82906 336852 82912 336864
rect 82867 336824 82912 336852
rect 82906 336812 82912 336824
rect 82964 336812 82970 336864
rect 3418 336744 3424 336796
rect 3476 336784 3482 336796
rect 72602 336784 72608 336796
rect 3476 336756 72608 336784
rect 3476 336744 3482 336756
rect 72602 336744 72608 336756
rect 72660 336744 72666 336796
rect 512822 336716 512828 336728
rect 512783 336688 512828 336716
rect 512822 336676 512828 336688
rect 512880 336676 512886 336728
rect 57790 335316 57796 335368
rect 57848 335356 57854 335368
rect 78674 335356 78680 335368
rect 57848 335328 78680 335356
rect 57848 335316 57854 335328
rect 78674 335316 78680 335328
rect 78732 335316 78738 335368
rect 504082 335248 504088 335300
rect 504140 335288 504146 335300
rect 569310 335288 569316 335300
rect 504140 335260 569316 335288
rect 504140 335248 504146 335260
rect 569310 335248 569316 335260
rect 569368 335248 569374 335300
rect 63034 332596 63040 332648
rect 63092 332636 63098 332648
rect 78674 332636 78680 332648
rect 63092 332608 78680 332636
rect 63092 332596 63098 332608
rect 78674 332596 78680 332608
rect 78732 332596 78738 332648
rect 17218 329740 17224 329792
rect 17276 329780 17282 329792
rect 78674 329780 78680 329792
rect 17276 329752 78680 329780
rect 17276 329740 17282 329752
rect 78674 329740 78680 329752
rect 78732 329740 78738 329792
rect 512822 327128 512828 327140
rect 512783 327100 512828 327128
rect 512822 327088 512828 327100
rect 512880 327088 512886 327140
rect 76650 324300 76656 324352
rect 76708 324340 76714 324352
rect 78674 324340 78680 324352
rect 76708 324312 78680 324340
rect 76708 324300 76714 324312
rect 78674 324300 78680 324312
rect 78732 324300 78738 324352
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 76558 324272 76564 324284
rect 3292 324244 76564 324272
rect 3292 324232 3298 324244
rect 76558 324232 76564 324244
rect 76616 324232 76622 324284
rect 504082 322940 504088 322992
rect 504140 322980 504146 322992
rect 512178 322980 512184 322992
rect 504140 322952 512184 322980
rect 504140 322940 504146 322952
rect 512178 322940 512184 322952
rect 512236 322940 512242 322992
rect 9122 322872 9128 322924
rect 9180 322912 9186 322924
rect 78674 322912 78680 322924
rect 9180 322884 78680 322912
rect 9180 322872 9186 322884
rect 78674 322872 78680 322884
rect 78732 322872 78738 322924
rect 514018 322872 514024 322924
rect 514076 322912 514082 322924
rect 580166 322912 580172 322924
rect 514076 322884 580172 322912
rect 514076 322872 514082 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 82814 318792 82820 318844
rect 82872 318832 82878 318844
rect 82906 318832 82912 318844
rect 82872 318804 82912 318832
rect 82872 318792 82878 318804
rect 82906 318792 82912 318804
rect 82964 318792 82970 318844
rect 504082 318792 504088 318844
rect 504140 318832 504146 318844
rect 515122 318832 515128 318844
rect 504140 318804 515128 318832
rect 504140 318792 504146 318804
rect 515122 318792 515128 318804
rect 515180 318792 515186 318844
rect 9122 317432 9128 317484
rect 9180 317472 9186 317484
rect 78674 317472 78680 317484
rect 9180 317444 78680 317472
rect 9180 317432 9186 317444
rect 78674 317432 78680 317444
rect 78732 317432 78738 317484
rect 512822 317364 512828 317416
rect 512880 317404 512886 317416
rect 512914 317404 512920 317416
rect 512880 317376 512920 317404
rect 512880 317364 512886 317376
rect 512914 317364 512920 317376
rect 512972 317364 512978 317416
rect 504082 316004 504088 316056
rect 504140 316044 504146 316056
rect 558178 316044 558184 316056
rect 504140 316016 558184 316044
rect 504140 316004 504146 316016
rect 558178 316004 558184 316016
rect 558236 316004 558242 316056
rect 72786 315936 72792 315988
rect 72844 315976 72850 315988
rect 73062 315976 73068 315988
rect 72844 315948 73068 315976
rect 72844 315936 72850 315948
rect 73062 315936 73068 315948
rect 73120 315936 73126 315988
rect 504358 314644 504364 314696
rect 504416 314684 504422 314696
rect 504450 314684 504456 314696
rect 504416 314656 504456 314684
rect 504416 314644 504422 314656
rect 504450 314644 504456 314656
rect 504508 314644 504514 314696
rect 515490 311788 515496 311840
rect 515548 311828 515554 311840
rect 580166 311828 580172 311840
rect 515548 311800 580172 311828
rect 515548 311788 515554 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 71314 310496 71320 310548
rect 71372 310536 71378 310548
rect 78674 310536 78680 310548
rect 71372 310508 78680 310536
rect 71372 310496 71378 310508
rect 78674 310496 78680 310508
rect 78732 310496 78738 310548
rect 3418 308932 3424 308984
rect 3476 308972 3482 308984
rect 9122 308972 9128 308984
rect 3476 308944 9128 308972
rect 3476 308932 3482 308944
rect 9122 308932 9128 308944
rect 9180 308932 9186 308984
rect 72786 306348 72792 306400
rect 72844 306388 72850 306400
rect 73062 306388 73068 306400
rect 72844 306360 73068 306388
rect 72844 306348 72850 306360
rect 73062 306348 73068 306360
rect 73120 306348 73126 306400
rect 504082 306280 504088 306332
rect 504140 306320 504146 306332
rect 567838 306320 567844 306332
rect 504140 306292 567844 306320
rect 504140 306280 504146 306292
rect 567838 306280 567844 306292
rect 567896 306280 567902 306332
rect 76558 299480 76564 299532
rect 76616 299520 76622 299532
rect 79226 299520 79232 299532
rect 76616 299492 79232 299520
rect 76616 299480 76622 299492
rect 79226 299480 79232 299492
rect 79284 299480 79290 299532
rect 82906 299520 82912 299532
rect 82867 299492 82912 299520
rect 82906 299480 82912 299492
rect 82964 299480 82970 299532
rect 540238 299412 540244 299464
rect 540296 299452 540302 299464
rect 579798 299452 579804 299464
rect 540296 299424 579804 299452
rect 540296 299412 540302 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 512822 298052 512828 298104
rect 512880 298092 512886 298104
rect 512914 298092 512920 298104
rect 512880 298064 512920 298092
rect 512880 298052 512886 298064
rect 512914 298052 512920 298064
rect 512972 298052 512978 298104
rect 72786 296624 72792 296676
rect 72844 296664 72850 296676
rect 73062 296664 73068 296676
rect 72844 296636 73068 296664
rect 72844 296624 72850 296636
rect 73062 296624 73068 296636
rect 73120 296624 73126 296676
rect 70118 295332 70124 295384
rect 70176 295372 70182 295384
rect 78674 295372 78680 295384
rect 70176 295344 78680 295372
rect 70176 295332 70182 295344
rect 78674 295332 78680 295344
rect 78732 295332 78738 295384
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 21358 295304 21364 295316
rect 3476 295276 21364 295304
rect 3476 295264 3482 295276
rect 21358 295264 21364 295276
rect 21416 295264 21422 295316
rect 82817 294763 82875 294769
rect 82817 294729 82829 294763
rect 82863 294760 82875 294763
rect 82906 294760 82912 294772
rect 82863 294732 82912 294760
rect 82863 294729 82875 294732
rect 82817 294723 82875 294729
rect 82906 294720 82912 294732
rect 82964 294720 82970 294772
rect 82906 294624 82912 294636
rect 82867 294596 82912 294624
rect 82906 294584 82912 294596
rect 82964 294584 82970 294636
rect 82817 294287 82875 294293
rect 82817 294253 82829 294287
rect 82863 294284 82875 294287
rect 82906 294284 82912 294296
rect 82863 294256 82912 294284
rect 82863 294253 82875 294256
rect 82817 294247 82875 294253
rect 82906 294244 82912 294256
rect 82964 294244 82970 294296
rect 504082 293972 504088 294024
rect 504140 294012 504146 294024
rect 512270 294012 512276 294024
rect 504140 293984 512276 294012
rect 504140 293972 504146 293984
rect 512270 293972 512276 293984
rect 512328 293972 512334 294024
rect 68554 292544 68560 292596
rect 68612 292584 68618 292596
rect 78674 292584 78680 292596
rect 68612 292556 78680 292584
rect 68612 292544 68618 292556
rect 78674 292544 78680 292556
rect 78732 292544 78738 292596
rect 504082 289824 504088 289876
rect 504140 289864 504146 289876
rect 508314 289864 508320 289876
rect 504140 289836 508320 289864
rect 504140 289824 504146 289836
rect 508314 289824 508320 289836
rect 508372 289824 508378 289876
rect 72786 287036 72792 287088
rect 72844 287076 72850 287088
rect 73062 287076 73068 287088
rect 72844 287048 73068 287076
rect 72844 287036 72850 287048
rect 73062 287036 73068 287048
rect 73120 287036 73126 287088
rect 504082 285676 504088 285728
rect 504140 285716 504146 285728
rect 540238 285716 540244 285728
rect 504140 285688 540244 285716
rect 504140 285676 504146 285688
rect 540238 285676 540244 285688
rect 540296 285676 540302 285728
rect 504082 282888 504088 282940
rect 504140 282928 504146 282940
rect 545114 282928 545120 282940
rect 504140 282900 545120 282928
rect 504140 282888 504146 282900
rect 545114 282888 545120 282900
rect 545172 282888 545178 282940
rect 72786 281528 72792 281580
rect 72844 281568 72850 281580
rect 78674 281568 78680 281580
rect 72844 281540 78680 281568
rect 72844 281528 72850 281540
rect 78674 281528 78680 281540
rect 78732 281528 78738 281580
rect 66990 277380 66996 277432
rect 67048 277420 67054 277432
rect 78674 277420 78680 277432
rect 67048 277392 78680 277420
rect 67048 277380 67054 277392
rect 78674 277380 78680 277392
rect 78732 277380 78738 277432
rect 72694 277312 72700 277364
rect 72752 277352 72758 277364
rect 73062 277352 73068 277364
rect 72752 277324 73068 277352
rect 72752 277312 72758 277324
rect 73062 277312 73068 277324
rect 73120 277312 73126 277364
rect 554038 275952 554044 276004
rect 554096 275992 554102 276004
rect 580166 275992 580172 276004
rect 554096 275964 580172 275992
rect 554096 275952 554102 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 504082 274660 504088 274712
rect 504140 274700 504146 274712
rect 519354 274700 519360 274712
rect 504140 274672 519360 274700
rect 504140 274660 504146 274672
rect 519354 274660 519360 274672
rect 519412 274660 519418 274712
rect 82906 273816 82912 273828
rect 82867 273788 82912 273816
rect 82906 273776 82912 273788
rect 82964 273776 82970 273828
rect 70026 273232 70032 273284
rect 70084 273272 70090 273284
rect 78674 273272 78680 273284
rect 70084 273244 78680 273272
rect 70084 273232 70090 273244
rect 78674 273232 78680 273244
rect 78732 273232 78738 273284
rect 512822 269084 512828 269136
rect 512880 269124 512886 269136
rect 513006 269124 513012 269136
rect 512880 269096 513012 269124
rect 512880 269084 512886 269096
rect 513006 269084 513012 269096
rect 513064 269084 513070 269136
rect 72694 267724 72700 267776
rect 72752 267764 72758 267776
rect 73062 267764 73068 267776
rect 72752 267736 73068 267764
rect 72752 267724 72758 267736
rect 73062 267724 73068 267736
rect 73120 267724 73126 267776
rect 504082 267724 504088 267776
rect 504140 267764 504146 267776
rect 515306 267764 515312 267776
rect 504140 267736 515312 267764
rect 504140 267724 504146 267736
rect 515306 267724 515312 267736
rect 515364 267724 515370 267776
rect 57698 266364 57704 266416
rect 57756 266404 57762 266416
rect 78674 266404 78680 266416
rect 57756 266376 78680 266404
rect 57756 266364 57762 266376
rect 78674 266364 78680 266376
rect 78732 266364 78738 266416
rect 3418 264936 3424 264988
rect 3476 264976 3482 264988
rect 68370 264976 68376 264988
rect 3476 264948 68376 264976
rect 3476 264936 3482 264948
rect 68370 264936 68376 264948
rect 68428 264936 68434 264988
rect 55858 263508 55864 263560
rect 55916 263548 55922 263560
rect 78674 263548 78680 263560
rect 55916 263520 78680 263548
rect 55916 263508 55922 263520
rect 78674 263508 78680 263520
rect 78732 263508 78738 263560
rect 504082 260856 504088 260908
rect 504140 260896 504146 260908
rect 507118 260896 507124 260908
rect 504140 260868 507124 260896
rect 504140 260856 504146 260868
rect 507118 260856 507124 260868
rect 507176 260856 507182 260908
rect 82906 259468 82912 259480
rect 82867 259440 82912 259468
rect 82906 259428 82912 259440
rect 82964 259428 82970 259480
rect 82814 259360 82820 259412
rect 82872 259400 82878 259412
rect 82872 259372 82952 259400
rect 82872 259360 82878 259372
rect 82924 259208 82952 259372
rect 82906 259156 82912 259208
rect 82964 259156 82970 259208
rect 72694 258748 72700 258800
rect 72752 258788 72758 258800
rect 73062 258788 73068 258800
rect 72752 258760 73068 258788
rect 72752 258748 72758 258760
rect 73062 258748 73068 258760
rect 73120 258748 73126 258800
rect 504082 256708 504088 256760
rect 504140 256748 504146 256760
rect 508130 256748 508136 256760
rect 504140 256720 508136 256748
rect 504140 256708 504146 256720
rect 508130 256708 508136 256720
rect 508188 256708 508194 256760
rect 66898 251268 66904 251320
rect 66956 251308 66962 251320
rect 78674 251308 78680 251320
rect 66956 251280 78680 251308
rect 66956 251268 66962 251280
rect 78674 251268 78680 251280
rect 78732 251268 78738 251320
rect 3418 251200 3424 251252
rect 3476 251240 3482 251252
rect 68462 251240 68468 251252
rect 3476 251212 68468 251240
rect 3476 251200 3482 251212
rect 68462 251200 68468 251212
rect 68520 251200 68526 251252
rect 567838 251200 567844 251252
rect 567896 251240 567902 251252
rect 580166 251240 580172 251252
rect 567896 251212 580172 251240
rect 567896 251200 567902 251212
rect 580166 251200 580172 251212
rect 580224 251200 580230 251252
rect 512822 249840 512828 249892
rect 512880 249880 512886 249892
rect 513006 249880 513012 249892
rect 512880 249852 513012 249880
rect 512880 249840 512886 249852
rect 513006 249840 513012 249852
rect 513064 249840 513070 249892
rect 504082 249772 504088 249824
rect 504140 249812 504146 249824
rect 518066 249812 518072 249824
rect 504140 249784 518072 249812
rect 504140 249772 504146 249784
rect 518066 249772 518072 249784
rect 518124 249772 518130 249824
rect 67082 249704 67088 249756
rect 67140 249744 67146 249756
rect 78674 249744 78680 249756
rect 67140 249716 78680 249744
rect 67140 249704 67146 249716
rect 78674 249704 78680 249716
rect 78732 249704 78738 249756
rect 72694 249092 72700 249144
rect 72752 249132 72758 249144
rect 73062 249132 73068 249144
rect 72752 249104 73068 249132
rect 72752 249092 72758 249104
rect 73062 249092 73068 249104
rect 73120 249092 73126 249144
rect 504082 245624 504088 245676
rect 504140 245664 504146 245676
rect 547138 245664 547144 245676
rect 504140 245636 547144 245664
rect 504140 245624 504146 245636
rect 547138 245624 547144 245636
rect 547196 245624 547202 245676
rect 78306 245556 78312 245608
rect 78364 245596 78370 245608
rect 79502 245596 79508 245608
rect 78364 245568 79508 245596
rect 78364 245556 78370 245568
rect 79502 245556 79508 245568
rect 79560 245556 79566 245608
rect 504082 242904 504088 242956
rect 504140 242944 504146 242956
rect 507026 242944 507032 242956
rect 504140 242916 507032 242944
rect 504140 242904 504146 242916
rect 507026 242904 507032 242916
rect 507084 242904 507090 242956
rect 73982 241476 73988 241528
rect 74040 241516 74046 241528
rect 78674 241516 78680 241528
rect 74040 241488 78680 241516
rect 74040 241476 74046 241488
rect 78674 241476 78680 241488
rect 78732 241476 78738 241528
rect 72694 239436 72700 239488
rect 72752 239476 72758 239488
rect 73062 239476 73068 239488
rect 72752 239448 73068 239476
rect 72752 239436 72758 239448
rect 73062 239436 73068 239448
rect 73120 239436 73126 239488
rect 69934 237396 69940 237448
rect 69992 237436 69998 237448
rect 78674 237436 78680 237448
rect 69992 237408 78680 237436
rect 69992 237396 69998 237408
rect 78674 237396 78680 237408
rect 78732 237396 78738 237448
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 69658 237368 69664 237380
rect 3476 237340 69664 237368
rect 3476 237328 3482 237340
rect 69658 237328 69664 237340
rect 69716 237328 69722 237380
rect 504082 234608 504088 234660
rect 504140 234648 504146 234660
rect 516686 234648 516692 234660
rect 504140 234620 516692 234648
rect 504140 234608 504146 234620
rect 516686 234608 516692 234620
rect 516744 234608 516750 234660
rect 55858 233248 55864 233300
rect 55916 233288 55922 233300
rect 78674 233288 78680 233300
rect 55916 233260 78680 233288
rect 55916 233248 55922 233260
rect 78674 233248 78680 233260
rect 78732 233248 78738 233300
rect 504082 231820 504088 231872
rect 504140 231860 504146 231872
rect 519538 231860 519544 231872
rect 504140 231832 519544 231860
rect 504140 231820 504146 231832
rect 519538 231820 519544 231832
rect 519596 231820 519602 231872
rect 519630 231412 519636 231464
rect 519688 231452 519694 231464
rect 520918 231452 520924 231464
rect 519688 231424 520924 231452
rect 519688 231412 519694 231424
rect 520918 231412 520924 231424
rect 520976 231412 520982 231464
rect 512822 230460 512828 230512
rect 512880 230500 512886 230512
rect 513006 230500 513012 230512
rect 512880 230472 513012 230500
rect 512880 230460 512886 230472
rect 513006 230460 513012 230472
rect 513064 230460 513070 230512
rect 72694 229712 72700 229764
rect 72752 229752 72758 229764
rect 73062 229752 73068 229764
rect 72752 229724 73068 229752
rect 72752 229712 72758 229724
rect 73062 229712 73068 229724
rect 73120 229712 73126 229764
rect 61470 229100 61476 229152
rect 61528 229140 61534 229152
rect 78674 229140 78680 229152
rect 61528 229112 78680 229140
rect 61528 229100 61534 229112
rect 78674 229100 78680 229112
rect 78732 229100 78738 229152
rect 531958 229032 531964 229084
rect 532016 229072 532022 229084
rect 580166 229072 580172 229084
rect 532016 229044 580172 229072
rect 532016 229032 532022 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 504082 227740 504088 227792
rect 504140 227780 504146 227792
rect 510890 227780 510896 227792
rect 504140 227752 510896 227780
rect 504140 227740 504146 227752
rect 510890 227740 510896 227752
rect 510948 227740 510954 227792
rect 504082 223592 504088 223644
rect 504140 223632 504146 223644
rect 512454 223632 512460 223644
rect 504140 223604 512460 223632
rect 504140 223592 504146 223604
rect 512454 223592 512460 223604
rect 512512 223592 512518 223644
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 72510 223564 72516 223576
rect 3200 223536 72516 223564
rect 3200 223524 3206 223536
rect 72510 223524 72516 223536
rect 72568 223524 72574 223576
rect 68738 223456 68744 223508
rect 68796 223496 68802 223508
rect 78674 223496 78680 223508
rect 68796 223468 78680 223496
rect 68796 223456 68802 223468
rect 78674 223456 78680 223468
rect 78732 223456 78738 223508
rect 504082 220872 504088 220924
rect 504140 220912 504146 220924
rect 509694 220912 509700 220924
rect 504140 220884 509700 220912
rect 504140 220872 504146 220884
rect 509694 220872 509700 220884
rect 509752 220872 509758 220924
rect 82817 219555 82875 219561
rect 82817 219521 82829 219555
rect 82863 219552 82875 219555
rect 82906 219552 82912 219564
rect 82863 219524 82912 219552
rect 82863 219521 82875 219524
rect 82817 219515 82875 219521
rect 82906 219512 82912 219524
rect 82964 219512 82970 219564
rect 82906 219008 82912 219020
rect 82867 218980 82912 219008
rect 82906 218968 82912 218980
rect 82964 218968 82970 219020
rect 540238 217948 540244 218000
rect 540296 217988 540302 218000
rect 580166 217988 580172 218000
rect 540296 217960 580172 217988
rect 540296 217948 540302 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 82817 217447 82875 217453
rect 82817 217413 82829 217447
rect 82863 217444 82875 217447
rect 82998 217444 83004 217456
rect 82863 217416 83004 217444
rect 82863 217413 82875 217416
rect 82817 217407 82875 217413
rect 82998 217404 83004 217416
rect 83056 217404 83062 217456
rect 72694 216928 72700 216980
rect 72752 216968 72758 216980
rect 73062 216968 73068 216980
rect 72752 216940 73068 216968
rect 72752 216928 72758 216940
rect 73062 216928 73068 216940
rect 73120 216928 73126 216980
rect 504082 212508 504088 212560
rect 504140 212548 504146 212560
rect 540238 212548 540244 212560
rect 504140 212520 540244 212548
rect 504140 212508 504146 212520
rect 540238 212508 540244 212520
rect 540296 212508 540302 212560
rect 72510 211148 72516 211200
rect 72568 211188 72574 211200
rect 78674 211188 78680 211200
rect 72568 211160 78680 211188
rect 72568 211148 72574 211160
rect 78674 211148 78680 211160
rect 78732 211148 78738 211200
rect 82725 210715 82783 210721
rect 82725 210681 82737 210715
rect 82771 210712 82783 210715
rect 82906 210712 82912 210724
rect 82771 210684 82912 210712
rect 82771 210681 82783 210684
rect 82725 210675 82783 210681
rect 82906 210672 82912 210684
rect 82964 210672 82970 210724
rect 72694 210400 72700 210452
rect 72752 210440 72758 210452
rect 73062 210440 73068 210452
rect 72752 210412 73068 210440
rect 72752 210400 72758 210412
rect 73062 210400 73068 210412
rect 73120 210400 73126 210452
rect 79502 210400 79508 210452
rect 79560 210440 79566 210452
rect 79686 210440 79692 210452
rect 79560 210412 79692 210440
rect 79560 210400 79566 210412
rect 79686 210400 79692 210412
rect 79744 210400 79750 210452
rect 82817 209967 82875 209973
rect 82817 209933 82829 209967
rect 82863 209964 82875 209967
rect 82906 209964 82912 209976
rect 82863 209936 82912 209964
rect 82863 209933 82875 209936
rect 82817 209927 82875 209933
rect 82906 209924 82912 209936
rect 82964 209924 82970 209976
rect 82725 209831 82783 209837
rect 82725 209797 82737 209831
rect 82771 209828 82783 209831
rect 82906 209828 82912 209840
rect 82771 209800 82912 209828
rect 82771 209797 82783 209800
rect 82725 209791 82783 209797
rect 82906 209788 82912 209800
rect 82964 209788 82970 209840
rect 504082 209788 504088 209840
rect 504140 209828 504146 209840
rect 512546 209828 512552 209840
rect 504140 209800 512552 209828
rect 504140 209788 504146 209800
rect 512546 209788 512552 209800
rect 512604 209788 512610 209840
rect 73890 208360 73896 208412
rect 73948 208400 73954 208412
rect 78674 208400 78680 208412
rect 73948 208372 78680 208400
rect 73948 208360 73954 208372
rect 78674 208360 78680 208372
rect 78732 208360 78738 208412
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 57238 208332 57244 208344
rect 3476 208304 57244 208332
rect 3476 208292 3482 208304
rect 57238 208292 57244 208304
rect 57296 208292 57302 208344
rect 82906 207720 82912 207732
rect 82867 207692 82912 207720
rect 82906 207680 82912 207692
rect 82964 207680 82970 207732
rect 82817 207519 82875 207525
rect 82817 207485 82829 207519
rect 82863 207516 82875 207519
rect 82906 207516 82912 207528
rect 82863 207488 82912 207516
rect 82863 207485 82875 207488
rect 82817 207479 82875 207485
rect 82906 207476 82912 207488
rect 82964 207476 82970 207528
rect 511442 204280 511448 204332
rect 511500 204320 511506 204332
rect 580166 204320 580172 204332
rect 511500 204292 580172 204320
rect 511500 204280 511506 204292
rect 580166 204280 580172 204292
rect 580224 204280 580230 204332
rect 512822 201424 512828 201476
rect 512880 201464 512886 201476
rect 513006 201464 513012 201476
rect 512880 201436 513012 201464
rect 512880 201424 512886 201436
rect 513006 201424 513012 201436
rect 513064 201424 513070 201476
rect 72326 200744 72332 200796
rect 72384 200784 72390 200796
rect 73062 200784 73068 200796
rect 72384 200756 73068 200784
rect 72384 200744 72390 200756
rect 73062 200744 73068 200756
rect 73120 200744 73126 200796
rect 79502 199520 79508 199572
rect 79560 199560 79566 199572
rect 79686 199560 79692 199572
rect 79560 199532 79692 199560
rect 79560 199520 79566 199532
rect 79686 199520 79692 199532
rect 79744 199520 79750 199572
rect 82906 195276 82912 195288
rect 82867 195248 82912 195276
rect 82906 195236 82912 195248
rect 82964 195236 82970 195288
rect 504174 194556 504180 194608
rect 504232 194596 504238 194608
rect 513926 194596 513932 194608
rect 504232 194568 513932 194596
rect 504232 194556 504238 194568
rect 513926 194556 513932 194568
rect 513984 194556 513990 194608
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 71130 194528 71136 194540
rect 3200 194500 71136 194528
rect 3200 194488 3206 194500
rect 71130 194488 71136 194500
rect 71188 194488 71194 194540
rect 504358 193808 504364 193860
rect 504416 193848 504422 193860
rect 515214 193848 515220 193860
rect 504416 193820 515220 193848
rect 504416 193808 504422 193820
rect 515214 193808 515220 193820
rect 515272 193808 515278 193860
rect 72694 193196 72700 193248
rect 72752 193236 72758 193248
rect 78674 193236 78680 193248
rect 72752 193208 78680 193236
rect 72752 193196 72758 193208
rect 78674 193196 78680 193208
rect 78732 193196 78738 193248
rect 68738 190476 68744 190528
rect 68796 190516 68802 190528
rect 78674 190516 78680 190528
rect 68796 190488 78680 190516
rect 68796 190476 68802 190488
rect 78674 190476 78680 190488
rect 78732 190476 78738 190528
rect 79502 190476 79508 190528
rect 79560 190516 79566 190528
rect 79686 190516 79692 190528
rect 79560 190488 79692 190516
rect 79560 190476 79566 190488
rect 79686 190476 79692 190488
rect 79744 190476 79750 190528
rect 504174 187688 504180 187740
rect 504232 187728 504238 187740
rect 554038 187728 554044 187740
rect 504232 187700 554044 187728
rect 504232 187688 504238 187700
rect 554038 187688 554044 187700
rect 554096 187688 554102 187740
rect 82906 182928 82912 182980
rect 82964 182928 82970 182980
rect 82924 182776 82952 182928
rect 82906 182724 82912 182776
rect 82964 182724 82970 182776
rect 71222 182180 71228 182232
rect 71280 182220 71286 182232
rect 78674 182220 78680 182232
rect 71280 182192 78680 182220
rect 71280 182180 71286 182192
rect 78674 182180 78680 182192
rect 78732 182180 78738 182232
rect 512822 182112 512828 182164
rect 512880 182152 512886 182164
rect 513006 182152 513012 182164
rect 512880 182124 513012 182152
rect 512880 182112 512886 182124
rect 513006 182112 513012 182124
rect 513064 182112 513070 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 20070 180792 20076 180804
rect 3292 180764 20076 180792
rect 3292 180752 3298 180764
rect 20070 180752 20076 180764
rect 20128 180752 20134 180804
rect 72326 180752 72332 180804
rect 72384 180792 72390 180804
rect 73062 180792 73068 180804
rect 72384 180764 73068 180792
rect 72384 180752 72390 180764
rect 73062 180752 73068 180764
rect 73120 180752 73126 180804
rect 79502 180752 79508 180804
rect 79560 180792 79566 180804
rect 79686 180792 79692 180804
rect 79560 180764 79692 180792
rect 79560 180752 79566 180764
rect 79686 180752 79692 180764
rect 79744 180752 79750 180804
rect 81066 179324 81072 179376
rect 81124 179364 81130 179376
rect 81894 179364 81900 179376
rect 81124 179336 81900 179364
rect 81124 179324 81130 179336
rect 81894 179324 81900 179336
rect 81952 179324 81958 179376
rect 75178 178100 75184 178152
rect 75236 178140 75242 178152
rect 82262 178140 82268 178152
rect 75236 178112 82268 178140
rect 75236 178100 75242 178112
rect 82262 178100 82268 178112
rect 82320 178100 82326 178152
rect 65702 178032 65708 178084
rect 65760 178072 65766 178084
rect 78674 178072 78680 178084
rect 65760 178044 78680 178072
rect 65760 178032 65766 178044
rect 78674 178032 78680 178044
rect 78732 178032 78738 178084
rect 79962 176672 79968 176724
rect 80020 176712 80026 176724
rect 80698 176712 80704 176724
rect 80020 176684 80704 176712
rect 80020 176672 80026 176684
rect 80698 176672 80704 176684
rect 80756 176672 80762 176724
rect 82725 173519 82783 173525
rect 82725 173485 82737 173519
rect 82771 173516 82783 173519
rect 82906 173516 82912 173528
rect 82771 173488 82912 173516
rect 82771 173485 82783 173488
rect 82725 173479 82783 173485
rect 82906 173476 82912 173488
rect 82964 173476 82970 173528
rect 82817 173383 82875 173389
rect 82817 173349 82829 173383
rect 82863 173380 82875 173383
rect 82906 173380 82912 173392
rect 82863 173352 82912 173380
rect 82863 173349 82875 173352
rect 82817 173343 82875 173349
rect 82906 173340 82912 173352
rect 82964 173340 82970 173392
rect 82725 172295 82783 172301
rect 82725 172261 82737 172295
rect 82771 172292 82783 172295
rect 82906 172292 82912 172304
rect 82771 172264 82912 172292
rect 82771 172261 82783 172264
rect 82725 172255 82783 172261
rect 82906 172252 82912 172264
rect 82964 172252 82970 172304
rect 509234 171776 509240 171828
rect 509292 171816 509298 171828
rect 527174 171816 527180 171828
rect 509292 171788 527180 171816
rect 509292 171776 509298 171788
rect 527174 171776 527180 171788
rect 527232 171776 527238 171828
rect 72326 171164 72332 171216
rect 72384 171204 72390 171216
rect 73062 171204 73068 171216
rect 72384 171176 73068 171204
rect 72384 171164 72390 171176
rect 73062 171164 73068 171176
rect 73120 171164 73126 171216
rect 65610 171096 65616 171148
rect 65668 171136 65674 171148
rect 78674 171136 78680 171148
rect 65668 171108 78680 171136
rect 65668 171096 65674 171108
rect 78674 171096 78680 171108
rect 78732 171096 78738 171148
rect 79502 171096 79508 171148
rect 79560 171136 79566 171148
rect 79686 171136 79692 171148
rect 79560 171108 79692 171136
rect 79560 171096 79566 171108
rect 79686 171096 79692 171108
rect 79744 171096 79750 171148
rect 511350 171028 511356 171080
rect 511408 171068 511414 171080
rect 580166 171068 580172 171080
rect 511408 171040 580172 171068
rect 511408 171028 511414 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 503714 170756 503720 170808
rect 503772 170796 503778 170808
rect 509234 170796 509240 170808
rect 503772 170768 509240 170796
rect 503772 170756 503778 170768
rect 509234 170756 509240 170768
rect 509292 170756 509298 170808
rect 79502 166268 79508 166320
rect 79560 166308 79566 166320
rect 79686 166308 79692 166320
rect 79560 166280 79692 166308
rect 79560 166268 79566 166280
rect 79686 166268 79692 166280
rect 79744 166268 79750 166320
rect 503714 165588 503720 165640
rect 503772 165628 503778 165640
rect 512362 165628 512368 165640
rect 503772 165600 512368 165628
rect 503772 165588 503778 165600
rect 512362 165588 512368 165600
rect 512420 165588 512426 165640
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 72418 165560 72424 165572
rect 3568 165532 72424 165560
rect 3568 165520 3574 165532
rect 72418 165520 72424 165532
rect 72476 165520 72482 165572
rect 68462 165452 68468 165504
rect 68520 165492 68526 165504
rect 78674 165492 78680 165504
rect 68520 165464 78680 165492
rect 68520 165452 68526 165464
rect 78674 165452 78680 165464
rect 78732 165452 78738 165504
rect 512822 162840 512828 162852
rect 512783 162812 512828 162840
rect 512822 162800 512828 162812
rect 512880 162800 512886 162852
rect 72418 161372 72424 161424
rect 72476 161412 72482 161424
rect 73062 161412 73068 161424
rect 72476 161384 73068 161412
rect 72476 161372 72482 161384
rect 73062 161372 73068 161384
rect 73120 161372 73126 161424
rect 14458 158652 14464 158704
rect 14516 158692 14522 158704
rect 78674 158692 78680 158704
rect 14516 158664 78680 158692
rect 14516 158652 14522 158664
rect 78674 158652 78680 158664
rect 78732 158652 78738 158704
rect 82725 158695 82783 158701
rect 82725 158661 82737 158695
rect 82771 158692 82783 158695
rect 82814 158692 82820 158704
rect 82771 158664 82820 158692
rect 82771 158661 82783 158664
rect 82725 158655 82783 158661
rect 82814 158652 82820 158664
rect 82872 158652 82878 158704
rect 573450 158652 573456 158704
rect 573508 158692 573514 158704
rect 579798 158692 579804 158704
rect 573508 158664 579804 158692
rect 573508 158652 573514 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 82817 158423 82875 158429
rect 82817 158389 82829 158423
rect 82863 158420 82875 158423
rect 82906 158420 82912 158432
rect 82863 158392 82912 158420
rect 82863 158389 82875 158392
rect 82817 158383 82875 158389
rect 82906 158380 82912 158392
rect 82964 158380 82970 158432
rect 82906 158012 82912 158024
rect 82867 157984 82912 158012
rect 82906 157972 82912 157984
rect 82964 157972 82970 158024
rect 82814 157836 82820 157888
rect 82872 157876 82878 157888
rect 82909 157879 82967 157885
rect 82909 157876 82921 157879
rect 82872 157848 82921 157876
rect 82872 157836 82878 157848
rect 82909 157845 82921 157848
rect 82955 157845 82967 157879
rect 82909 157839 82967 157845
rect 82722 157400 82728 157412
rect 82683 157372 82728 157400
rect 82722 157360 82728 157372
rect 82780 157360 82786 157412
rect 69658 155184 69664 155236
rect 69716 155224 69722 155236
rect 82170 155224 82176 155236
rect 69716 155196 82176 155224
rect 69716 155184 69722 155196
rect 82170 155184 82176 155196
rect 82228 155184 82234 155236
rect 68462 153212 68468 153264
rect 68520 153252 68526 153264
rect 78674 153252 78680 153264
rect 68520 153224 78680 153252
rect 68520 153212 68526 153224
rect 78674 153212 78680 153224
rect 78732 153212 78738 153264
rect 512822 153252 512828 153264
rect 512783 153224 512828 153252
rect 512822 153212 512828 153224
rect 512880 153212 512886 153264
rect 72418 151784 72424 151836
rect 72476 151824 72482 151836
rect 73062 151824 73068 151836
rect 72476 151796 73068 151824
rect 72476 151784 72482 151796
rect 73062 151784 73068 151796
rect 73120 151784 73126 151836
rect 79502 151784 79508 151836
rect 79560 151824 79566 151836
rect 79686 151824 79692 151836
rect 79560 151796 79692 151824
rect 79560 151784 79566 151796
rect 79686 151784 79692 151796
rect 79744 151784 79750 151836
rect 503714 151784 503720 151836
rect 503772 151824 503778 151836
rect 552750 151824 552756 151836
rect 503772 151796 552756 151824
rect 503772 151784 503778 151796
rect 552750 151784 552756 151796
rect 552808 151784 552814 151836
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 68278 151756 68284 151768
rect 3200 151728 68284 151756
rect 3200 151716 3206 151728
rect 68278 151716 68284 151728
rect 68336 151716 68342 151768
rect 14458 149064 14464 149116
rect 14516 149104 14522 149116
rect 78674 149104 78680 149116
rect 14516 149076 78680 149104
rect 14516 149064 14522 149076
rect 78674 149064 78680 149076
rect 78732 149064 78738 149116
rect 82633 148291 82691 148297
rect 82633 148257 82645 148291
rect 82679 148288 82691 148291
rect 82906 148288 82912 148300
rect 82679 148260 82912 148288
rect 82679 148257 82691 148260
rect 82633 148251 82691 148257
rect 82906 148248 82912 148260
rect 82964 148248 82970 148300
rect 17218 146276 17224 146328
rect 17276 146316 17282 146328
rect 78674 146316 78680 146328
rect 17276 146288 78680 146316
rect 17276 146276 17282 146288
rect 78674 146276 78680 146288
rect 78732 146276 78738 146328
rect 82817 145231 82875 145237
rect 82817 145197 82829 145231
rect 82863 145228 82875 145231
rect 82906 145228 82912 145240
rect 82863 145200 82912 145228
rect 82863 145197 82875 145200
rect 82817 145191 82875 145197
rect 82906 145188 82912 145200
rect 82964 145188 82970 145240
rect 82725 145027 82783 145033
rect 82725 144993 82737 145027
rect 82771 145024 82783 145027
rect 82906 145024 82912 145036
rect 82771 144996 82912 145024
rect 82771 144993 82783 144996
rect 82725 144987 82783 144993
rect 82906 144984 82912 144996
rect 82964 144984 82970 145036
rect 82633 144891 82691 144897
rect 82633 144857 82645 144891
rect 82679 144888 82691 144891
rect 82814 144888 82820 144900
rect 82679 144860 82820 144888
rect 82679 144857 82691 144860
rect 82633 144851 82691 144857
rect 82814 144848 82820 144860
rect 82872 144848 82878 144900
rect 82906 144780 82912 144832
rect 82964 144820 82970 144832
rect 82964 144792 83009 144820
rect 82964 144780 82970 144792
rect 82817 143735 82875 143741
rect 82817 143701 82829 143735
rect 82863 143732 82875 143735
rect 82906 143732 82912 143744
rect 82863 143704 82912 143732
rect 82863 143701 82875 143704
rect 82817 143695 82875 143701
rect 82906 143692 82912 143704
rect 82964 143692 82970 143744
rect 82725 143599 82783 143605
rect 82725 143565 82737 143599
rect 82771 143596 82783 143599
rect 82906 143596 82912 143608
rect 82771 143568 82912 143596
rect 82771 143565 82783 143568
rect 82725 143559 82783 143565
rect 82906 143556 82912 143568
rect 82964 143556 82970 143608
rect 504542 143556 504548 143608
rect 504600 143596 504606 143608
rect 510982 143596 510988 143608
rect 504600 143568 510988 143596
rect 504600 143556 504606 143568
rect 510982 143556 510988 143568
rect 511040 143556 511046 143608
rect 512822 143528 512828 143540
rect 512783 143500 512828 143528
rect 512822 143488 512828 143500
rect 512880 143488 512886 143540
rect 72418 142060 72424 142112
rect 72476 142100 72482 142112
rect 73062 142100 73068 142112
rect 72476 142072 73068 142100
rect 72476 142060 72482 142072
rect 73062 142060 73068 142072
rect 73120 142060 73126 142112
rect 79686 142060 79692 142112
rect 79744 142100 79750 142112
rect 79962 142100 79968 142112
rect 79744 142072 79968 142100
rect 79744 142060 79750 142072
rect 79962 142060 79968 142072
rect 80020 142060 80026 142112
rect 504542 140768 504548 140820
rect 504600 140808 504606 140820
rect 508406 140808 508412 140820
rect 504600 140780 508412 140808
rect 504600 140768 504606 140780
rect 508406 140768 508412 140780
rect 508464 140768 508470 140820
rect 82814 140224 82820 140276
rect 82872 140264 82878 140276
rect 82872 140236 82917 140264
rect 82872 140224 82878 140236
rect 71130 140020 71136 140072
rect 71188 140060 71194 140072
rect 82906 140060 82912 140072
rect 71188 140032 82912 140060
rect 71188 140020 71194 140032
rect 82906 140020 82912 140032
rect 82964 140020 82970 140072
rect 82814 137164 82820 137216
rect 82872 137204 82878 137216
rect 82872 137176 82917 137204
rect 82872 137164 82878 137176
rect 3510 135804 3516 135856
rect 3568 135844 3574 135856
rect 9122 135844 9128 135856
rect 3568 135816 9128 135844
rect 3568 135804 3574 135816
rect 9122 135804 9128 135816
rect 9180 135804 9186 135856
rect 552658 135192 552664 135244
rect 552716 135232 552722 135244
rect 580166 135232 580172 135244
rect 552716 135204 580172 135232
rect 552716 135192 552722 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 82630 134716 82636 134768
rect 82688 134756 82694 134768
rect 82906 134756 82912 134768
rect 82688 134728 82912 134756
rect 82688 134716 82694 134728
rect 82906 134716 82912 134728
rect 82964 134716 82970 134768
rect 512822 133940 512828 133952
rect 512783 133912 512828 133940
rect 512822 133900 512828 133912
rect 512880 133900 512886 133952
rect 503070 133016 503076 133068
rect 503128 133056 503134 133068
rect 508498 133056 508504 133068
rect 503128 133028 508504 133056
rect 503128 133016 503134 133028
rect 508498 133016 508504 133028
rect 508556 133016 508562 133068
rect 82906 132608 82912 132660
rect 82964 132648 82970 132660
rect 82964 132620 83044 132648
rect 82964 132608 82970 132620
rect 72418 132472 72424 132524
rect 72476 132512 72482 132524
rect 73062 132512 73068 132524
rect 72476 132484 73068 132512
rect 72476 132472 72482 132484
rect 73062 132472 73068 132484
rect 73120 132472 73126 132524
rect 79686 132472 79692 132524
rect 79744 132512 79750 132524
rect 79962 132512 79968 132524
rect 79744 132484 79968 132512
rect 79744 132472 79750 132484
rect 79962 132472 79968 132484
rect 80020 132472 80026 132524
rect 82538 132472 82544 132524
rect 82596 132512 82602 132524
rect 83016 132512 83044 132620
rect 82596 132484 83044 132512
rect 82596 132472 82602 132484
rect 57238 131112 57244 131164
rect 57296 131152 57302 131164
rect 78674 131152 78680 131164
rect 57296 131124 78680 131152
rect 57296 131112 57302 131124
rect 78674 131112 78680 131124
rect 78732 131112 78738 131164
rect 72418 126964 72424 127016
rect 72476 127004 72482 127016
rect 78674 127004 78680 127016
rect 72476 126976 78680 127004
rect 72476 126964 72482 126976
rect 78674 126964 78680 126976
rect 78732 126964 78738 127016
rect 73798 126216 73804 126268
rect 73856 126256 73862 126268
rect 79318 126256 79324 126268
rect 73856 126228 79324 126256
rect 73856 126216 73862 126228
rect 79318 126216 79324 126228
rect 79376 126216 79382 126268
rect 504542 125604 504548 125656
rect 504600 125644 504606 125656
rect 509786 125644 509792 125656
rect 504600 125616 509792 125644
rect 504600 125604 504606 125616
rect 509786 125604 509792 125616
rect 509844 125604 509850 125656
rect 82817 124219 82875 124225
rect 82817 124185 82829 124219
rect 82863 124216 82875 124219
rect 82906 124216 82912 124228
rect 82863 124188 82912 124216
rect 82863 124185 82875 124188
rect 82817 124179 82875 124185
rect 82906 124176 82912 124188
rect 82964 124176 82970 124228
rect 512822 124148 512828 124160
rect 512783 124120 512828 124148
rect 512822 124108 512828 124120
rect 512880 124108 512886 124160
rect 538858 124108 538864 124160
rect 538916 124148 538922 124160
rect 580166 124148 580172 124160
rect 538916 124120 580172 124148
rect 538916 124108 538922 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 82906 124080 82912 124092
rect 82867 124052 82912 124080
rect 82906 124040 82912 124052
rect 82964 124040 82970 124092
rect 72326 122748 72332 122800
rect 72384 122788 72390 122800
rect 73062 122788 73068 122800
rect 72384 122760 73068 122788
rect 72384 122748 72390 122760
rect 73062 122748 73068 122760
rect 73120 122748 73126 122800
rect 79686 122748 79692 122800
rect 79744 122788 79750 122800
rect 79962 122788 79968 122800
rect 79744 122760 79968 122788
rect 79744 122748 79750 122760
rect 79962 122748 79968 122760
rect 80020 122748 80026 122800
rect 3418 121456 3424 121508
rect 3476 121496 3482 121508
rect 11698 121496 11704 121508
rect 3476 121468 11704 121496
rect 3476 121456 3482 121468
rect 11698 121456 11704 121468
rect 11756 121456 11762 121508
rect 81066 120028 81072 120080
rect 81124 120068 81130 120080
rect 81894 120068 81900 120080
rect 81124 120040 81900 120068
rect 81124 120028 81130 120040
rect 81894 120028 81900 120040
rect 81952 120028 81958 120080
rect 82906 118708 82912 118720
rect 82867 118680 82912 118708
rect 82906 118668 82912 118680
rect 82964 118668 82970 118720
rect 82906 115240 82912 115252
rect 82867 115212 82912 115240
rect 82906 115200 82912 115212
rect 82964 115200 82970 115252
rect 512822 114560 512828 114572
rect 512783 114532 512828 114560
rect 512822 114520 512828 114532
rect 512880 114520 512886 114572
rect 72326 113160 72332 113212
rect 72384 113200 72390 113212
rect 73062 113200 73068 113212
rect 72384 113172 73068 113200
rect 72384 113160 72390 113172
rect 73062 113160 73068 113172
rect 73120 113160 73126 113212
rect 79686 113160 79692 113212
rect 79744 113200 79750 113212
rect 79962 113200 79968 113212
rect 79744 113172 79968 113200
rect 79744 113160 79750 113172
rect 79962 113160 79968 113172
rect 80020 113160 80026 113212
rect 82817 111027 82875 111033
rect 82817 110993 82829 111027
rect 82863 111024 82875 111027
rect 82906 111024 82912 111036
rect 82863 110996 82912 111024
rect 82863 110993 82875 110996
rect 82817 110987 82875 110993
rect 82906 110984 82912 110996
rect 82964 110984 82970 111036
rect 503254 110440 503260 110492
rect 503312 110480 503318 110492
rect 509234 110480 509240 110492
rect 503312 110452 509240 110480
rect 503312 110440 503318 110452
rect 509234 110440 509240 110452
rect 509292 110440 509298 110492
rect 73062 110372 73068 110424
rect 73120 110412 73126 110424
rect 78674 110412 78680 110424
rect 73120 110384 78680 110412
rect 73120 110372 73126 110384
rect 78674 110372 78680 110384
rect 78732 110372 78738 110424
rect 73062 109012 73068 109064
rect 73120 109052 73126 109064
rect 73798 109052 73804 109064
rect 73120 109024 73804 109052
rect 73120 109012 73126 109024
rect 73798 109012 73804 109024
rect 73856 109012 73862 109064
rect 73798 107856 73804 107908
rect 73856 107896 73862 107908
rect 74166 107896 74172 107908
rect 73856 107868 74172 107896
rect 73856 107856 73862 107868
rect 74166 107856 74172 107868
rect 74224 107856 74230 107908
rect 4062 107652 4068 107704
rect 4120 107692 4126 107704
rect 74258 107692 74264 107704
rect 4120 107664 74264 107692
rect 4120 107652 4126 107664
rect 74258 107652 74264 107664
rect 74316 107652 74322 107704
rect 503346 107652 503352 107704
rect 503404 107692 503410 107704
rect 531958 107692 531964 107704
rect 503404 107664 531964 107692
rect 503404 107652 503410 107664
rect 531958 107652 531964 107664
rect 532016 107652 532022 107704
rect 503898 107516 503904 107568
rect 503956 107556 503962 107568
rect 504358 107556 504364 107568
rect 503956 107528 504364 107556
rect 503956 107516 503962 107528
rect 504358 107516 504364 107528
rect 504416 107516 504422 107568
rect 82630 106700 82636 106752
rect 82688 106740 82694 106752
rect 82906 106740 82912 106752
rect 82688 106712 82912 106740
rect 82688 106700 82694 106712
rect 82906 106700 82912 106712
rect 82964 106700 82970 106752
rect 502978 105476 502984 105528
rect 503036 105516 503042 105528
rect 504450 105516 504456 105528
rect 503036 105488 504456 105516
rect 503036 105476 503042 105488
rect 504450 105476 504456 105488
rect 504508 105476 504514 105528
rect 82998 104836 83004 104848
rect 82924 104808 83004 104836
rect 82924 104780 82952 104808
rect 82998 104796 83004 104808
rect 83056 104796 83062 104848
rect 512641 104839 512699 104845
rect 512641 104805 512653 104839
rect 512687 104836 512699 104839
rect 512822 104836 512828 104848
rect 512687 104808 512828 104836
rect 512687 104805 512699 104808
rect 512641 104799 512699 104805
rect 512822 104796 512828 104808
rect 512880 104796 512886 104848
rect 82906 104728 82912 104780
rect 82964 104728 82970 104780
rect 504542 103504 504548 103556
rect 504600 103544 504606 103556
rect 511350 103544 511356 103556
rect 504600 103516 511356 103544
rect 504600 103504 504606 103516
rect 511350 103504 511356 103516
rect 511408 103504 511414 103556
rect 38657 103139 38715 103145
rect 38657 103105 38669 103139
rect 38703 103136 38715 103139
rect 50985 103139 51043 103145
rect 50985 103136 50997 103139
rect 38703 103108 50997 103136
rect 38703 103105 38715 103108
rect 38657 103099 38715 103105
rect 50985 103105 50997 103108
rect 51031 103105 51043 103139
rect 50985 103099 51043 103105
rect 51077 103071 51135 103077
rect 51077 103037 51089 103071
rect 51123 103068 51135 103071
rect 56597 103071 56655 103077
rect 56597 103068 56609 103071
rect 51123 103040 56609 103068
rect 51123 103037 51135 103040
rect 51077 103031 51135 103037
rect 56597 103037 56609 103040
rect 56643 103037 56655 103071
rect 56597 103031 56655 103037
rect 19337 103003 19395 103009
rect 19337 102969 19349 103003
rect 19383 103000 19395 103003
rect 19383 102972 29868 103000
rect 19383 102969 19395 102972
rect 19337 102963 19395 102969
rect 19337 102867 19395 102873
rect 19337 102864 19349 102867
rect 19260 102836 19349 102864
rect 19260 102805 19288 102836
rect 19337 102833 19349 102836
rect 19383 102833 19395 102867
rect 19337 102827 19395 102833
rect 19245 102799 19303 102805
rect 19245 102765 19257 102799
rect 19291 102765 19303 102799
rect 29840 102796 29868 102972
rect 66165 102935 66223 102941
rect 66165 102901 66177 102935
rect 66211 102932 66223 102935
rect 66211 102904 71268 102932
rect 66211 102901 66223 102904
rect 66165 102895 66223 102901
rect 38657 102799 38715 102805
rect 38657 102796 38669 102799
rect 29840 102768 38669 102796
rect 19245 102759 19303 102765
rect 38657 102765 38669 102768
rect 38703 102765 38715 102799
rect 38657 102759 38715 102765
rect 56597 102799 56655 102805
rect 56597 102765 56609 102799
rect 56643 102796 56655 102799
rect 66165 102799 66223 102805
rect 66165 102796 66177 102799
rect 56643 102768 66177 102796
rect 56643 102765 56655 102768
rect 56597 102759 56655 102765
rect 66165 102765 66177 102768
rect 66211 102765 66223 102799
rect 66165 102759 66223 102765
rect 9122 102688 9128 102740
rect 9180 102728 9186 102740
rect 9677 102731 9735 102737
rect 9677 102728 9689 102731
rect 9180 102700 9689 102728
rect 9180 102688 9186 102700
rect 9677 102697 9689 102700
rect 9723 102697 9735 102731
rect 9677 102691 9735 102697
rect 9677 102595 9735 102601
rect 9677 102561 9689 102595
rect 9723 102592 9735 102595
rect 19245 102595 19303 102601
rect 19245 102592 19257 102595
rect 9723 102564 19257 102592
rect 9723 102561 9735 102564
rect 9677 102555 9735 102561
rect 19245 102561 19257 102564
rect 19291 102561 19303 102595
rect 19245 102555 19303 102561
rect 71240 102456 71268 102904
rect 509234 102864 509240 102876
rect 142724 102836 144960 102864
rect 82722 102756 82728 102808
rect 82780 102796 82786 102808
rect 142724 102805 142752 102836
rect 144932 102805 144960 102836
rect 162780 102836 162900 102864
rect 162780 102805 162808 102836
rect 162872 102805 162900 102836
rect 187436 102836 193260 102864
rect 91281 102799 91339 102805
rect 91281 102796 91293 102799
rect 82780 102768 91293 102796
rect 82780 102756 82786 102768
rect 91281 102765 91293 102768
rect 91327 102765 91339 102799
rect 91281 102759 91339 102765
rect 104161 102799 104219 102805
rect 104161 102765 104173 102799
rect 104207 102796 104219 102799
rect 113821 102799 113879 102805
rect 113821 102796 113833 102799
rect 104207 102768 113833 102796
rect 104207 102765 104219 102768
rect 104161 102759 104219 102765
rect 113821 102765 113833 102768
rect 113867 102765 113879 102799
rect 113821 102759 113879 102765
rect 120721 102799 120779 102805
rect 120721 102765 120733 102799
rect 120767 102796 120779 102799
rect 127345 102799 127403 102805
rect 127345 102796 127357 102799
rect 120767 102768 127357 102796
rect 120767 102765 120779 102768
rect 120721 102759 120779 102765
rect 127345 102765 127357 102768
rect 127391 102765 127403 102799
rect 127345 102759 127403 102765
rect 142709 102799 142767 102805
rect 142709 102765 142721 102799
rect 142755 102765 142767 102799
rect 142709 102759 142767 102765
rect 144917 102799 144975 102805
rect 144917 102765 144929 102799
rect 144963 102765 144975 102799
rect 144917 102759 144975 102765
rect 162765 102799 162823 102805
rect 162765 102765 162777 102799
rect 162811 102765 162823 102799
rect 162765 102759 162823 102765
rect 162857 102799 162915 102805
rect 162857 102765 162869 102799
rect 162903 102765 162915 102799
rect 162857 102759 162915 102765
rect 182085 102799 182143 102805
rect 182085 102765 182097 102799
rect 182131 102796 182143 102799
rect 187436 102796 187464 102836
rect 193232 102805 193260 102836
rect 381556 102836 386368 102864
rect 182131 102768 187464 102796
rect 193217 102799 193275 102805
rect 182131 102765 182143 102768
rect 182085 102759 182143 102765
rect 193217 102765 193229 102799
rect 193263 102765 193275 102799
rect 193217 102759 193275 102765
rect 201696 102768 205588 102796
rect 81066 102688 81072 102740
rect 81124 102728 81130 102740
rect 183557 102731 183615 102737
rect 183557 102728 183569 102731
rect 81124 102700 183569 102728
rect 81124 102688 81130 102700
rect 183557 102697 183569 102700
rect 183603 102697 183615 102731
rect 201494 102728 201500 102740
rect 183557 102691 183615 102697
rect 183848 102700 201500 102728
rect 72970 102620 72976 102672
rect 73028 102660 73034 102672
rect 183649 102663 183707 102669
rect 73028 102632 183600 102660
rect 73028 102620 73034 102632
rect 74166 102552 74172 102604
rect 74224 102592 74230 102604
rect 173986 102592 173992 102604
rect 74224 102564 173992 102592
rect 74224 102552 74230 102564
rect 173986 102552 173992 102564
rect 174044 102552 174050 102604
rect 183572 102601 183600 102632
rect 183649 102629 183661 102663
rect 183695 102660 183707 102663
rect 183848 102660 183876 102700
rect 201494 102688 201500 102700
rect 201552 102688 201558 102740
rect 183695 102632 183876 102660
rect 193217 102663 193275 102669
rect 183695 102629 183707 102632
rect 183649 102623 183707 102629
rect 193217 102629 193229 102663
rect 193263 102660 193275 102663
rect 201696 102660 201724 102768
rect 205560 102728 205588 102768
rect 234632 102768 244320 102796
rect 215205 102731 215263 102737
rect 215205 102728 215217 102731
rect 205560 102700 215217 102728
rect 215205 102697 215217 102700
rect 215251 102697 215263 102731
rect 215205 102691 215263 102697
rect 215297 102731 215355 102737
rect 215297 102697 215309 102731
rect 215343 102728 215355 102731
rect 226981 102731 227039 102737
rect 215343 102700 216536 102728
rect 215343 102697 215355 102700
rect 215297 102691 215355 102697
rect 193263 102632 201724 102660
rect 216508 102660 216536 102700
rect 226981 102697 226993 102731
rect 227027 102728 227039 102731
rect 234632 102728 234660 102768
rect 227027 102700 234660 102728
rect 244292 102728 244320 102768
rect 253952 102768 263640 102796
rect 253952 102728 253980 102768
rect 244292 102700 253980 102728
rect 263612 102728 263640 102768
rect 370608 102768 374040 102796
rect 280525 102731 280583 102737
rect 280525 102728 280537 102731
rect 263612 102700 280537 102728
rect 227027 102697 227039 102700
rect 226981 102691 227039 102697
rect 280525 102697 280537 102700
rect 280571 102697 280583 102731
rect 280525 102691 280583 102697
rect 222197 102663 222255 102669
rect 222197 102660 222209 102663
rect 216508 102632 222209 102660
rect 193263 102629 193275 102632
rect 193217 102623 193275 102629
rect 222197 102629 222209 102632
rect 222243 102629 222255 102663
rect 222197 102623 222255 102629
rect 370498 102620 370504 102672
rect 370556 102660 370562 102672
rect 370608 102660 370636 102768
rect 374012 102728 374040 102768
rect 381556 102728 381584 102836
rect 386340 102805 386368 102836
rect 394620 102836 396028 102864
rect 394620 102805 394648 102836
rect 386325 102799 386383 102805
rect 386325 102765 386337 102799
rect 386371 102765 386383 102799
rect 386325 102759 386383 102765
rect 394605 102799 394663 102805
rect 394605 102765 394617 102799
rect 394651 102765 394663 102799
rect 396000 102796 396028 102836
rect 416700 102836 509240 102864
rect 416700 102805 416728 102836
rect 509234 102824 509240 102836
rect 509292 102824 509298 102876
rect 416593 102799 416651 102805
rect 416593 102796 416605 102799
rect 396000 102768 416605 102796
rect 394605 102759 394663 102765
rect 416593 102765 416605 102768
rect 416639 102765 416651 102799
rect 416593 102759 416651 102765
rect 416685 102799 416743 102805
rect 416685 102765 416697 102799
rect 416731 102765 416743 102799
rect 416685 102759 416743 102765
rect 416777 102799 416835 102805
rect 416777 102765 416789 102799
rect 416823 102796 416835 102799
rect 523402 102796 523408 102808
rect 416823 102768 523408 102796
rect 416823 102765 416835 102768
rect 416777 102759 416835 102765
rect 523402 102756 523408 102768
rect 523460 102756 523466 102808
rect 374012 102700 381584 102728
rect 370556 102632 370636 102660
rect 386325 102663 386383 102669
rect 370556 102620 370562 102632
rect 386325 102629 386337 102663
rect 386371 102660 386383 102663
rect 394605 102663 394663 102669
rect 394605 102660 394617 102663
rect 386371 102632 394617 102660
rect 386371 102629 386383 102632
rect 386325 102623 386383 102629
rect 394605 102629 394617 102632
rect 394651 102629 394663 102663
rect 394605 102623 394663 102629
rect 416682 102620 416688 102672
rect 416740 102660 416746 102672
rect 416740 102632 416785 102660
rect 416740 102620 416746 102632
rect 183557 102595 183615 102601
rect 183557 102561 183569 102595
rect 183603 102561 183615 102595
rect 183557 102555 183615 102561
rect 80149 102527 80207 102533
rect 80149 102493 80161 102527
rect 80195 102524 80207 102527
rect 103517 102527 103575 102533
rect 80195 102496 87000 102524
rect 80195 102493 80207 102496
rect 80149 102487 80207 102493
rect 79965 102459 80023 102465
rect 79965 102456 79977 102459
rect 71240 102428 79977 102456
rect 79965 102425 79977 102428
rect 80011 102425 80023 102459
rect 79965 102419 80023 102425
rect 83090 102416 83096 102468
rect 83148 102456 83154 102468
rect 83642 102456 83648 102468
rect 83148 102428 83648 102456
rect 83148 102416 83154 102428
rect 83642 102416 83648 102428
rect 83700 102416 83706 102468
rect 86972 102465 87000 102496
rect 103517 102493 103529 102527
rect 103563 102524 103575 102527
rect 103563 102496 109080 102524
rect 103563 102493 103575 102496
rect 103517 102487 103575 102493
rect 86957 102459 87015 102465
rect 86957 102425 86969 102459
rect 87003 102425 87015 102459
rect 86957 102419 87015 102425
rect 91281 102459 91339 102465
rect 91281 102425 91293 102459
rect 91327 102456 91339 102459
rect 104161 102459 104219 102465
rect 104161 102456 104173 102459
rect 91327 102428 104173 102456
rect 91327 102425 91339 102428
rect 91281 102419 91339 102425
rect 104161 102425 104173 102428
rect 104207 102425 104219 102459
rect 104161 102419 104219 102425
rect 79870 102348 79876 102400
rect 79928 102388 79934 102400
rect 84838 102388 84844 102400
rect 79928 102360 84844 102388
rect 79928 102348 79934 102360
rect 84838 102348 84844 102360
rect 84896 102348 84902 102400
rect 87049 102391 87107 102397
rect 87049 102357 87061 102391
rect 87095 102388 87107 102391
rect 103517 102391 103575 102397
rect 87095 102360 103468 102388
rect 87095 102357 87107 102360
rect 87049 102351 87107 102357
rect 82909 102323 82967 102329
rect 82909 102289 82921 102323
rect 82955 102320 82967 102323
rect 83366 102320 83372 102332
rect 82955 102292 83372 102320
rect 82955 102289 82967 102292
rect 82909 102283 82967 102289
rect 83366 102280 83372 102292
rect 83424 102280 83430 102332
rect 103440 102320 103468 102360
rect 103517 102357 103529 102391
rect 103563 102357 103575 102391
rect 109052 102388 109080 102496
rect 125502 102484 125508 102536
rect 125560 102524 125566 102536
rect 133690 102524 133696 102536
rect 125560 102496 133696 102524
rect 125560 102484 125566 102496
rect 133690 102484 133696 102496
rect 133748 102484 133754 102536
rect 144917 102527 144975 102533
rect 144917 102493 144929 102527
rect 144963 102524 144975 102527
rect 153197 102527 153255 102533
rect 153197 102524 153209 102527
rect 144963 102496 153209 102524
rect 144963 102493 144975 102496
rect 144917 102487 144975 102493
rect 153197 102493 153209 102496
rect 153243 102493 153255 102527
rect 153197 102487 153255 102493
rect 162857 102527 162915 102533
rect 162857 102493 162869 102527
rect 162903 102524 162915 102527
rect 172517 102527 172575 102533
rect 172517 102524 172529 102527
rect 162903 102496 172529 102524
rect 162903 102493 162915 102496
rect 162857 102487 162915 102493
rect 172517 102493 172529 102496
rect 172563 102493 172575 102527
rect 172517 102487 172575 102493
rect 222197 102527 222255 102533
rect 222197 102493 222209 102527
rect 222243 102524 222255 102527
rect 226981 102527 227039 102533
rect 226981 102524 226993 102527
rect 222243 102496 226993 102524
rect 222243 102493 222255 102496
rect 222197 102487 222255 102493
rect 226981 102493 226993 102496
rect 227027 102493 227039 102527
rect 226981 102487 227039 102493
rect 113821 102459 113879 102465
rect 113821 102425 113833 102459
rect 113867 102456 113879 102459
rect 120721 102459 120779 102465
rect 120721 102456 120733 102459
rect 113867 102428 120733 102456
rect 113867 102425 113879 102428
rect 113821 102419 113879 102425
rect 120721 102425 120733 102428
rect 120767 102425 120779 102459
rect 120721 102419 120779 102425
rect 127345 102459 127403 102465
rect 127345 102425 127357 102459
rect 127391 102456 127403 102459
rect 142709 102459 142767 102465
rect 142709 102456 142721 102459
rect 127391 102428 142721 102456
rect 127391 102425 127403 102428
rect 127345 102419 127403 102425
rect 142709 102425 142721 102428
rect 142755 102425 142767 102459
rect 149054 102456 149060 102468
rect 142709 102419 142767 102425
rect 142816 102428 149060 102456
rect 115937 102391 115995 102397
rect 115937 102388 115949 102391
rect 109052 102360 115949 102388
rect 103517 102351 103575 102357
rect 115937 102357 115949 102360
rect 115983 102357 115995 102391
rect 115937 102351 115995 102357
rect 138017 102391 138075 102397
rect 138017 102357 138029 102391
rect 138063 102388 138075 102391
rect 142816 102388 142844 102428
rect 149054 102416 149060 102428
rect 149112 102416 149118 102468
rect 138063 102360 142844 102388
rect 153197 102391 153255 102397
rect 138063 102357 138075 102360
rect 138017 102351 138075 102357
rect 153197 102357 153209 102391
rect 153243 102388 153255 102391
rect 162765 102391 162823 102397
rect 162765 102388 162777 102391
rect 153243 102360 162777 102388
rect 153243 102357 153255 102360
rect 153197 102351 153255 102357
rect 162765 102357 162777 102360
rect 162811 102357 162823 102391
rect 162765 102351 162823 102357
rect 172517 102391 172575 102397
rect 172517 102357 172529 102391
rect 172563 102388 172575 102391
rect 182085 102391 182143 102397
rect 182085 102388 182097 102391
rect 172563 102360 182097 102388
rect 172563 102357 172575 102360
rect 172517 102351 172575 102357
rect 182085 102357 182097 102360
rect 182131 102357 182143 102391
rect 182085 102351 182143 102357
rect 103532 102320 103560 102351
rect 103440 102292 103560 102320
rect 125597 102323 125655 102329
rect 125597 102289 125609 102323
rect 125643 102320 125655 102323
rect 137925 102323 137983 102329
rect 137925 102320 137937 102323
rect 125643 102292 137937 102320
rect 125643 102289 125655 102292
rect 125597 102283 125655 102289
rect 137925 102289 137937 102292
rect 137971 102289 137983 102323
rect 137925 102283 137983 102289
rect 79686 102212 79692 102264
rect 79744 102252 79750 102264
rect 79870 102252 79876 102264
rect 79744 102224 79876 102252
rect 79744 102212 79750 102224
rect 79870 102212 79876 102224
rect 79928 102212 79934 102264
rect 115937 102187 115995 102193
rect 115937 102153 115949 102187
rect 115983 102184 115995 102187
rect 125597 102187 125655 102193
rect 125597 102184 125609 102187
rect 115983 102156 125609 102184
rect 115983 102153 115995 102156
rect 115937 102147 115995 102153
rect 125597 102153 125609 102156
rect 125643 102153 125655 102187
rect 125597 102147 125655 102153
rect 74258 102076 74264 102128
rect 74316 102116 74322 102128
rect 510890 102116 510896 102128
rect 74316 102088 510896 102116
rect 74316 102076 74322 102088
rect 510890 102076 510896 102088
rect 510948 102076 510954 102128
rect 499482 101940 499488 101992
rect 499540 101980 499546 101992
rect 513834 101980 513840 101992
rect 499540 101952 513840 101980
rect 499540 101940 499546 101952
rect 513834 101940 513840 101952
rect 513892 101940 513898 101992
rect 81986 101872 81992 101924
rect 82044 101912 82050 101924
rect 106458 101912 106464 101924
rect 82044 101884 106464 101912
rect 82044 101872 82050 101884
rect 106458 101872 106464 101884
rect 106516 101872 106522 101924
rect 488442 101872 488448 101924
rect 488500 101912 488506 101924
rect 508498 101912 508504 101924
rect 488500 101884 508504 101912
rect 488500 101872 488506 101884
rect 508498 101872 508504 101884
rect 508556 101872 508562 101924
rect 83642 101804 83648 101856
rect 83700 101844 83706 101856
rect 107654 101844 107660 101856
rect 83700 101816 107660 101844
rect 83700 101804 83706 101816
rect 107654 101804 107660 101816
rect 107712 101804 107718 101856
rect 183557 101847 183615 101853
rect 183557 101813 183569 101847
rect 183603 101844 183615 101847
rect 187786 101844 187792 101856
rect 183603 101816 187792 101844
rect 183603 101813 183615 101816
rect 183557 101807 183615 101813
rect 187786 101804 187792 101816
rect 187844 101804 187850 101856
rect 480070 101804 480076 101856
rect 480128 101844 480134 101856
rect 502518 101844 502524 101856
rect 480128 101816 502524 101844
rect 480128 101804 480134 101816
rect 502518 101804 502524 101816
rect 502576 101804 502582 101856
rect 67174 101736 67180 101788
rect 67232 101776 67238 101788
rect 93946 101776 93952 101788
rect 67232 101748 93952 101776
rect 67232 101736 67238 101748
rect 93946 101736 93952 101748
rect 94004 101736 94010 101788
rect 487062 101736 487068 101788
rect 487120 101776 487126 101788
rect 509786 101776 509792 101788
rect 487120 101748 509792 101776
rect 487120 101736 487126 101748
rect 509786 101736 509792 101748
rect 509844 101736 509850 101788
rect 56502 101668 56508 101720
rect 56560 101708 56566 101720
rect 88518 101708 88524 101720
rect 56560 101680 88524 101708
rect 56560 101668 56566 101680
rect 88518 101668 88524 101680
rect 88576 101668 88582 101720
rect 484302 101668 484308 101720
rect 484360 101708 484366 101720
rect 513926 101708 513932 101720
rect 484360 101680 513932 101708
rect 484360 101668 484366 101680
rect 513926 101668 513932 101680
rect 513984 101668 513990 101720
rect 71590 101600 71596 101652
rect 71648 101640 71654 101652
rect 103606 101640 103612 101652
rect 71648 101612 103612 101640
rect 71648 101600 71654 101612
rect 103606 101600 103612 101612
rect 103664 101600 103670 101652
rect 453942 101600 453948 101652
rect 454000 101640 454006 101652
rect 505646 101640 505652 101652
rect 454000 101612 505652 101640
rect 454000 101600 454006 101612
rect 505646 101600 505652 101612
rect 505704 101600 505710 101652
rect 75546 101532 75552 101584
rect 75604 101572 75610 101584
rect 117314 101572 117320 101584
rect 75604 101544 117320 101572
rect 75604 101532 75610 101544
rect 117314 101532 117320 101544
rect 117372 101532 117378 101584
rect 439498 101532 439504 101584
rect 439556 101572 439562 101584
rect 504358 101572 504364 101584
rect 439556 101544 504364 101572
rect 439556 101532 439562 101544
rect 504358 101532 504364 101544
rect 504416 101532 504422 101584
rect 80974 101464 80980 101516
rect 81032 101504 81038 101516
rect 128354 101504 128360 101516
rect 81032 101476 128360 101504
rect 81032 101464 81038 101476
rect 128354 101464 128360 101476
rect 128412 101464 128418 101516
rect 198734 101464 198740 101516
rect 198792 101504 198798 101516
rect 512454 101504 512460 101516
rect 198792 101476 512460 101504
rect 198792 101464 198798 101476
rect 512454 101464 512460 101476
rect 512512 101464 512518 101516
rect 85574 101396 85580 101448
rect 85632 101436 85638 101448
rect 495250 101436 495256 101448
rect 85632 101408 495256 101436
rect 85632 101396 85638 101408
rect 495250 101396 495256 101408
rect 495308 101396 495314 101448
rect 500862 101396 500868 101448
rect 500920 101436 500926 101448
rect 519170 101436 519176 101448
rect 500920 101408 519176 101436
rect 500920 101396 500926 101408
rect 519170 101396 519176 101408
rect 519228 101396 519234 101448
rect 82170 101260 82176 101312
rect 82228 101300 82234 101312
rect 85574 101300 85580 101312
rect 82228 101272 85580 101300
rect 82228 101260 82234 101272
rect 85574 101260 85580 101272
rect 85632 101260 85638 101312
rect 88334 100852 88340 100904
rect 88392 100892 88398 100904
rect 419442 100892 419448 100904
rect 88392 100864 419448 100892
rect 88392 100852 88398 100864
rect 419442 100852 419448 100864
rect 419500 100852 419506 100904
rect 39298 100784 39304 100836
rect 39356 100824 39362 100836
rect 166442 100824 166448 100836
rect 39356 100796 166448 100824
rect 39356 100784 39362 100796
rect 166442 100784 166448 100796
rect 166500 100784 166506 100836
rect 245562 100784 245568 100836
rect 245620 100824 245626 100836
rect 511442 100824 511448 100836
rect 245620 100796 511448 100824
rect 245620 100784 245626 100796
rect 511442 100784 511448 100796
rect 511500 100784 511506 100836
rect 72602 100716 72608 100768
rect 72660 100756 72666 100768
rect 467834 100756 467840 100768
rect 72660 100728 467840 100756
rect 72660 100716 72666 100728
rect 467834 100716 467840 100728
rect 467892 100716 467898 100768
rect 513282 100716 513288 100768
rect 513340 100756 513346 100768
rect 520918 100756 520924 100768
rect 513340 100728 520924 100756
rect 513340 100716 513346 100728
rect 520918 100716 520924 100728
rect 520976 100716 520982 100768
rect 11698 100648 11704 100700
rect 11756 100688 11762 100700
rect 285122 100688 285128 100700
rect 11756 100660 285128 100688
rect 11756 100648 11762 100660
rect 285122 100648 285128 100660
rect 285180 100648 285186 100700
rect 292482 100648 292488 100700
rect 292540 100688 292546 100700
rect 514110 100688 514116 100700
rect 292540 100660 514116 100688
rect 292540 100648 292546 100660
rect 514110 100648 514116 100660
rect 514168 100648 514174 100700
rect 68370 100580 68376 100632
rect 68428 100620 68434 100632
rect 322106 100620 322112 100632
rect 68428 100592 322112 100620
rect 68428 100580 68434 100592
rect 322106 100580 322112 100592
rect 322164 100580 322170 100632
rect 327074 100580 327080 100632
rect 327132 100620 327138 100632
rect 516778 100620 516784 100632
rect 327132 100592 516784 100620
rect 327132 100580 327138 100592
rect 516778 100580 516784 100592
rect 516836 100580 516842 100632
rect 82538 100512 82544 100564
rect 82596 100552 82602 100564
rect 84930 100552 84936 100564
rect 82596 100524 84936 100552
rect 82596 100512 82602 100524
rect 84930 100512 84936 100524
rect 84988 100512 84994 100564
rect 85025 100555 85083 100561
rect 85025 100521 85037 100555
rect 85071 100552 85083 100555
rect 329466 100552 329472 100564
rect 85071 100524 329472 100552
rect 85071 100521 85083 100524
rect 85025 100515 85083 100521
rect 329466 100512 329472 100524
rect 329524 100512 329530 100564
rect 359090 100512 359096 100564
rect 359148 100552 359154 100564
rect 360102 100552 360108 100564
rect 359148 100524 360108 100552
rect 359148 100512 359154 100524
rect 360102 100512 360108 100524
rect 360160 100512 360166 100564
rect 410978 100512 410984 100564
rect 411036 100552 411042 100564
rect 560938 100552 560944 100564
rect 411036 100524 560944 100552
rect 411036 100512 411042 100524
rect 560938 100512 560944 100524
rect 560996 100512 561002 100564
rect 68830 100444 68836 100496
rect 68888 100484 68894 100496
rect 186130 100484 186136 100496
rect 68888 100456 186136 100484
rect 68888 100444 68894 100456
rect 186130 100444 186136 100456
rect 186188 100444 186194 100496
rect 218330 100444 218336 100496
rect 218388 100484 218394 100496
rect 219342 100484 219348 100496
rect 218388 100456 219348 100484
rect 218388 100444 218394 100456
rect 219342 100444 219348 100456
rect 219400 100444 219406 100496
rect 230658 100444 230664 100496
rect 230716 100484 230722 100496
rect 231762 100484 231768 100496
rect 230716 100456 231768 100484
rect 230716 100444 230722 100456
rect 231762 100444 231768 100456
rect 231820 100444 231826 100496
rect 255314 100444 255320 100496
rect 255372 100484 255378 100496
rect 256602 100484 256608 100496
rect 255372 100456 256608 100484
rect 255372 100444 255378 100456
rect 256602 100444 256608 100456
rect 256660 100444 256666 100496
rect 267826 100444 267832 100496
rect 267884 100484 267890 100496
rect 269022 100484 269028 100496
rect 267884 100456 269028 100484
rect 267884 100444 267890 100456
rect 269022 100444 269028 100456
rect 269080 100444 269086 100496
rect 280154 100444 280160 100496
rect 280212 100484 280218 100496
rect 281442 100484 281448 100496
rect 280212 100456 281448 100484
rect 280212 100444 280218 100456
rect 281442 100444 281448 100456
rect 281500 100444 281506 100496
rect 388898 100444 388904 100496
rect 388956 100484 388962 100496
rect 511258 100484 511264 100496
rect 388956 100456 511264 100484
rect 388956 100444 388962 100456
rect 511258 100444 511264 100456
rect 511316 100444 511322 100496
rect 69750 100376 69756 100428
rect 69808 100416 69814 100428
rect 176378 100416 176384 100428
rect 69808 100388 176384 100416
rect 69808 100376 69814 100388
rect 176378 100376 176384 100388
rect 176436 100376 176442 100428
rect 401226 100376 401232 100428
rect 401284 100416 401290 100428
rect 520458 100416 520464 100428
rect 401284 100388 520464 100416
rect 401284 100376 401290 100388
rect 520458 100376 520464 100388
rect 520516 100376 520522 100428
rect 71498 100308 71504 100360
rect 71556 100348 71562 100360
rect 164050 100348 164056 100360
rect 71556 100320 164056 100348
rect 71556 100308 71562 100320
rect 164050 100308 164056 100320
rect 164108 100308 164114 100360
rect 403618 100308 403624 100360
rect 403676 100348 403682 100360
rect 515398 100348 515404 100360
rect 403676 100320 515404 100348
rect 403676 100308 403682 100320
rect 515398 100308 515404 100320
rect 515456 100308 515462 100360
rect 70302 100240 70308 100292
rect 70360 100280 70366 100292
rect 131850 100280 131856 100292
rect 70360 100252 131856 100280
rect 70360 100240 70366 100252
rect 131850 100240 131856 100252
rect 131908 100240 131914 100292
rect 136818 100240 136824 100292
rect 136876 100280 136882 100292
rect 137922 100280 137928 100292
rect 136876 100252 137928 100280
rect 136876 100240 136882 100252
rect 137922 100240 137928 100252
rect 137980 100240 137986 100292
rect 206002 100240 206008 100292
rect 206060 100280 206066 100292
rect 206922 100280 206928 100292
rect 206060 100252 206928 100280
rect 206060 100240 206066 100252
rect 206922 100240 206928 100252
rect 206980 100240 206986 100292
rect 207658 100240 207664 100292
rect 207716 100280 207722 100292
rect 277578 100280 277584 100292
rect 207716 100252 277584 100280
rect 207716 100240 207722 100252
rect 277578 100240 277584 100252
rect 277636 100240 277642 100292
rect 286318 100240 286324 100292
rect 286376 100280 286382 100292
rect 314746 100280 314752 100292
rect 286376 100252 314752 100280
rect 286376 100240 286382 100252
rect 314746 100240 314752 100252
rect 314804 100240 314810 100292
rect 327718 100240 327724 100292
rect 327776 100280 327782 100292
rect 341794 100280 341800 100292
rect 327776 100252 341800 100280
rect 327776 100240 327782 100252
rect 341794 100240 341800 100252
rect 341852 100240 341858 100292
rect 356517 100283 356575 100289
rect 356517 100249 356529 100283
rect 356563 100280 356575 100283
rect 376386 100280 376392 100292
rect 356563 100252 376392 100280
rect 356563 100249 356575 100252
rect 356517 100243 356575 100249
rect 376386 100240 376392 100252
rect 376444 100240 376450 100292
rect 419442 100240 419448 100292
rect 419500 100280 419506 100292
rect 440786 100280 440792 100292
rect 419500 100252 440792 100280
rect 419500 100240 419506 100252
rect 440786 100240 440792 100252
rect 440844 100240 440850 100292
rect 455506 100240 455512 100292
rect 455564 100280 455570 100292
rect 456702 100280 456708 100292
rect 455564 100252 456708 100280
rect 455564 100240 455570 100252
rect 456702 100240 456708 100252
rect 456760 100240 456766 100292
rect 475378 100240 475384 100292
rect 475436 100280 475442 100292
rect 509970 100280 509976 100292
rect 475436 100252 509976 100280
rect 475436 100240 475442 100252
rect 509970 100240 509976 100252
rect 510028 100240 510034 100292
rect 75822 100172 75828 100224
rect 75880 100212 75886 100224
rect 112162 100212 112168 100224
rect 75880 100184 112168 100212
rect 75880 100172 75886 100184
rect 112162 100172 112168 100184
rect 112220 100172 112226 100224
rect 114554 100172 114560 100224
rect 114612 100212 114618 100224
rect 115842 100212 115848 100224
rect 114612 100184 115848 100212
rect 114612 100172 114618 100184
rect 115842 100172 115848 100184
rect 115900 100172 115906 100224
rect 124858 100172 124864 100224
rect 124916 100212 124922 100224
rect 126882 100212 126888 100224
rect 124916 100184 126888 100212
rect 124916 100172 124922 100184
rect 126882 100172 126888 100184
rect 126940 100172 126946 100224
rect 240778 100172 240784 100224
rect 240836 100212 240842 100224
rect 356698 100212 356704 100224
rect 240836 100184 356704 100212
rect 240836 100172 240842 100184
rect 356698 100172 356704 100184
rect 356756 100172 356762 100224
rect 370590 100172 370596 100224
rect 370648 100212 370654 100224
rect 408586 100212 408592 100224
rect 370648 100184 408592 100212
rect 370648 100172 370654 100184
rect 408586 100172 408592 100184
rect 408644 100172 408650 100224
rect 81342 100104 81348 100156
rect 81400 100144 81406 100156
rect 85025 100147 85083 100153
rect 85025 100144 85037 100147
rect 81400 100116 85037 100144
rect 81400 100104 81406 100116
rect 85025 100113 85037 100116
rect 85071 100113 85083 100147
rect 85025 100107 85083 100113
rect 89898 100104 89904 100156
rect 89956 100144 89962 100156
rect 91002 100144 91008 100156
rect 89956 100116 91008 100144
rect 89956 100104 89962 100116
rect 91002 100104 91008 100116
rect 91060 100104 91066 100156
rect 99650 100104 99656 100156
rect 99708 100144 99714 100156
rect 100662 100144 100668 100156
rect 99708 100116 100668 100144
rect 99708 100104 99714 100116
rect 100662 100104 100668 100116
rect 100720 100104 100726 100156
rect 117958 100104 117964 100156
rect 118016 100144 118022 100156
rect 159082 100144 159088 100156
rect 118016 100116 159088 100144
rect 118016 100104 118022 100116
rect 159082 100104 159088 100116
rect 159140 100104 159146 100156
rect 186958 100104 186964 100156
rect 187016 100144 187022 100156
rect 213362 100144 213368 100156
rect 187016 100116 213368 100144
rect 187016 100104 187022 100116
rect 213362 100104 213368 100116
rect 213420 100104 213426 100156
rect 261478 100104 261484 100156
rect 261536 100144 261542 100156
rect 393682 100144 393688 100156
rect 261536 100116 393688 100144
rect 261536 100104 261542 100116
rect 393682 100104 393688 100116
rect 393740 100104 393746 100156
rect 83550 100036 83556 100088
rect 83608 100076 83614 100088
rect 99466 100076 99472 100088
rect 83608 100048 99472 100076
rect 83608 100036 83614 100048
rect 99466 100036 99472 100048
rect 99524 100036 99530 100088
rect 142798 100036 142804 100088
rect 142856 100076 142862 100088
rect 198642 100076 198648 100088
rect 142856 100048 198648 100076
rect 142856 100036 142862 100048
rect 198642 100036 198648 100048
rect 198700 100036 198706 100088
rect 225598 100036 225604 100088
rect 225656 100076 225662 100088
rect 240594 100076 240600 100088
rect 225656 100048 240600 100076
rect 225656 100036 225662 100048
rect 240594 100036 240600 100048
rect 240652 100036 240658 100088
rect 251818 100036 251824 100088
rect 251876 100076 251882 100088
rect 406194 100076 406200 100088
rect 251876 100048 406200 100076
rect 251876 100036 251882 100048
rect 406194 100036 406200 100048
rect 406252 100036 406258 100088
rect 478782 100036 478788 100088
rect 478840 100076 478846 100088
rect 505738 100076 505744 100088
rect 478840 100048 505744 100076
rect 478840 100036 478846 100048
rect 505738 100036 505744 100048
rect 505796 100036 505802 100088
rect 81434 99968 81440 100020
rect 81492 100008 81498 100020
rect 110414 100008 110420 100020
rect 81492 99980 110420 100008
rect 81492 99968 81498 99980
rect 110414 99968 110420 99980
rect 110472 99968 110478 100020
rect 131758 99968 131764 100020
rect 131816 100008 131822 100020
rect 139210 100008 139216 100020
rect 131816 99980 139216 100008
rect 131816 99968 131822 99980
rect 139210 99968 139216 99980
rect 139268 99968 139274 100020
rect 149698 99968 149704 100020
rect 149756 100008 149762 100020
rect 260282 100008 260288 100020
rect 149756 99980 260288 100008
rect 149756 99968 149762 99980
rect 260282 99968 260288 99980
rect 260340 99968 260346 100020
rect 302142 99968 302148 100020
rect 302200 100008 302206 100020
rect 521838 100008 521844 100020
rect 302200 99980 521844 100008
rect 302200 99968 302206 99980
rect 521838 99968 521844 99980
rect 521896 99968 521902 100020
rect 477770 99900 477776 99952
rect 477828 99940 477834 99952
rect 478690 99940 478696 99952
rect 477828 99912 478696 99940
rect 477828 99900 477834 99912
rect 478690 99900 478696 99912
rect 478748 99900 478754 99952
rect 102226 99832 102232 99884
rect 102284 99872 102290 99884
rect 103422 99872 103428 99884
rect 102284 99844 103428 99872
rect 102284 99832 102290 99844
rect 103422 99832 103428 99844
rect 103480 99832 103486 99884
rect 121914 99696 121920 99748
rect 121972 99736 121978 99748
rect 122742 99736 122748 99748
rect 121972 99708 122748 99736
rect 121972 99696 121978 99708
rect 122742 99696 122748 99708
rect 122800 99696 122806 99748
rect 265250 99628 265256 99680
rect 265308 99668 265314 99680
rect 266262 99668 266268 99680
rect 265308 99640 266268 99668
rect 265308 99628 265314 99640
rect 266262 99628 266268 99640
rect 266320 99628 266326 99680
rect 287514 99356 287520 99408
rect 287572 99396 287578 99408
rect 288342 99396 288348 99408
rect 287572 99368 288348 99396
rect 287572 99356 287578 99368
rect 288342 99356 288348 99368
rect 288400 99356 288406 99408
rect 315298 99356 315304 99408
rect 315356 99396 315362 99408
rect 317138 99396 317144 99408
rect 315356 99368 317144 99396
rect 315356 99356 315362 99368
rect 317138 99356 317144 99368
rect 317196 99356 317202 99408
rect 323578 99356 323584 99408
rect 323636 99396 323642 99408
rect 324498 99396 324504 99408
rect 323636 99368 324504 99396
rect 323636 99356 323642 99368
rect 324498 99356 324504 99368
rect 324556 99356 324562 99408
rect 334434 99356 334440 99408
rect 334492 99396 334498 99408
rect 335262 99396 335268 99408
rect 334492 99368 335268 99396
rect 334492 99356 334498 99368
rect 335262 99356 335268 99368
rect 335320 99356 335326 99408
rect 373994 99356 374000 99408
rect 374052 99396 374058 99408
rect 375282 99396 375288 99408
rect 374052 99368 375288 99396
rect 374052 99356 374058 99368
rect 375282 99356 375288 99368
rect 375340 99356 375346 99408
rect 381354 99356 381360 99408
rect 381412 99396 381418 99408
rect 382182 99396 382188 99408
rect 381412 99368 382188 99396
rect 381412 99356 381418 99368
rect 382182 99356 382188 99368
rect 382240 99356 382246 99408
rect 383930 99356 383936 99408
rect 383988 99396 383994 99408
rect 384942 99396 384948 99408
rect 383988 99368 384948 99396
rect 383988 99356 383994 99368
rect 384942 99356 384948 99368
rect 385000 99356 385006 99408
rect 494698 99356 494704 99408
rect 494756 99396 494762 99408
rect 500034 99396 500040 99408
rect 494756 99368 500040 99396
rect 494756 99356 494762 99368
rect 500034 99356 500040 99368
rect 500092 99356 500098 99408
rect 183738 99288 183744 99340
rect 183796 99328 183802 99340
rect 184842 99328 184848 99340
rect 183796 99300 184848 99328
rect 183796 99288 183802 99300
rect 184842 99288 184848 99300
rect 184900 99288 184906 99340
rect 280522 99328 280528 99340
rect 280483 99300 280528 99328
rect 280522 99288 280528 99300
rect 280580 99288 280586 99340
rect 469122 99288 469128 99340
rect 469180 99328 469186 99340
rect 502886 99328 502892 99340
rect 469180 99300 502892 99328
rect 469180 99288 469186 99300
rect 502886 99288 502892 99300
rect 502944 99288 502950 99340
rect 503070 99288 503076 99340
rect 503128 99328 503134 99340
rect 513282 99328 513288 99340
rect 503128 99300 513288 99328
rect 503128 99288 503134 99300
rect 513282 99288 513288 99300
rect 513340 99288 513346 99340
rect 78398 99220 78404 99272
rect 78456 99260 78462 99272
rect 132586 99260 132592 99272
rect 78456 99232 132592 99260
rect 78456 99220 78462 99232
rect 132586 99220 132592 99232
rect 132644 99220 132650 99272
rect 486970 99220 486976 99272
rect 487028 99260 487034 99272
rect 523310 99260 523316 99272
rect 487028 99232 523316 99260
rect 487028 99220 487034 99232
rect 523310 99220 523316 99232
rect 523368 99220 523374 99272
rect 70210 99152 70216 99204
rect 70268 99192 70274 99204
rect 142154 99192 142160 99204
rect 70268 99164 142160 99192
rect 70268 99152 70274 99164
rect 142154 99152 142160 99164
rect 142212 99152 142218 99204
rect 419442 99152 419448 99204
rect 419500 99192 419506 99204
rect 518986 99192 518992 99204
rect 419500 99164 518992 99192
rect 419500 99152 419506 99164
rect 518986 99152 518992 99164
rect 519044 99152 519050 99204
rect 75638 99084 75644 99136
rect 75696 99124 75702 99136
rect 149054 99124 149060 99136
rect 75696 99096 149060 99124
rect 75696 99084 75702 99096
rect 149054 99084 149060 99096
rect 149112 99084 149118 99136
rect 354582 99084 354588 99136
rect 354640 99124 354646 99136
rect 512270 99124 512276 99136
rect 354640 99096 512276 99124
rect 354640 99084 354646 99096
rect 512270 99084 512276 99096
rect 512328 99084 512334 99136
rect 71406 99016 71412 99068
rect 71464 99056 71470 99068
rect 146294 99056 146300 99068
rect 71464 99028 146300 99056
rect 71464 99016 71470 99028
rect 146294 99016 146300 99028
rect 146352 99016 146358 99068
rect 331122 99016 331128 99068
rect 331180 99056 331186 99068
rect 520642 99056 520648 99068
rect 331180 99028 520648 99056
rect 331180 99016 331186 99028
rect 520642 99016 520648 99028
rect 520700 99016 520706 99068
rect 66162 98948 66168 99000
rect 66220 98988 66226 99000
rect 166994 98988 167000 99000
rect 66220 98960 167000 98988
rect 66220 98948 66226 98960
rect 166994 98948 167000 98960
rect 167052 98948 167058 99000
rect 306282 98948 306288 99000
rect 306340 98988 306346 99000
rect 510798 98988 510804 99000
rect 306340 98960 510804 98988
rect 306340 98948 306346 98960
rect 510798 98948 510804 98960
rect 510856 98948 510862 99000
rect 80698 98880 80704 98932
rect 80756 98920 80762 98932
rect 193214 98920 193220 98932
rect 80756 98892 193220 98920
rect 80756 98880 80762 98892
rect 193214 98880 193220 98892
rect 193272 98880 193278 98932
rect 284202 98880 284208 98932
rect 284260 98920 284266 98932
rect 512546 98920 512552 98932
rect 284260 98892 512552 98920
rect 284260 98880 284266 98892
rect 512546 98880 512552 98892
rect 512604 98880 512610 98932
rect 61746 98812 61752 98864
rect 61804 98852 61810 98864
rect 179414 98852 179420 98864
rect 61804 98824 179420 98852
rect 61804 98812 61810 98824
rect 179414 98812 179420 98824
rect 179472 98812 179478 98864
rect 251082 98812 251088 98864
rect 251140 98852 251146 98864
rect 503990 98852 503996 98864
rect 251140 98824 503996 98852
rect 251140 98812 251146 98824
rect 503990 98812 503996 98824
rect 504048 98812 504054 98864
rect 77938 98744 77944 98796
rect 77996 98784 78002 98796
rect 195974 98784 195980 98796
rect 77996 98756 195980 98784
rect 77996 98744 78002 98756
rect 195974 98744 195980 98756
rect 196032 98744 196038 98796
rect 241422 98744 241428 98796
rect 241480 98784 241486 98796
rect 515122 98784 515128 98796
rect 241480 98756 515128 98784
rect 241480 98744 241486 98756
rect 515122 98744 515128 98756
rect 515180 98744 515186 98796
rect 67266 98676 67272 98728
rect 67324 98716 67330 98728
rect 218054 98716 218060 98728
rect 67324 98688 218060 98716
rect 67324 98676 67330 98688
rect 218054 98676 218060 98688
rect 218112 98676 218118 98728
rect 227622 98676 227628 98728
rect 227680 98716 227686 98728
rect 509694 98716 509700 98728
rect 227680 98688 509700 98716
rect 227680 98676 227686 98688
rect 509694 98676 509700 98688
rect 509752 98676 509758 98728
rect 81158 98608 81164 98660
rect 81216 98648 81222 98660
rect 207014 98648 207020 98660
rect 81216 98620 207020 98648
rect 81216 98608 81222 98620
rect 207014 98608 207020 98620
rect 207072 98608 207078 98660
rect 216582 98608 216588 98660
rect 216640 98648 216646 98660
rect 519078 98648 519084 98660
rect 216640 98620 519084 98648
rect 216640 98608 216646 98620
rect 519078 98608 519084 98620
rect 519136 98608 519142 98660
rect 187694 97996 187700 98048
rect 187752 98036 187758 98048
rect 188430 98036 188436 98048
rect 187752 98008 188436 98036
rect 187752 97996 187758 98008
rect 188430 97996 188436 98008
rect 188488 97996 188494 98048
rect 25498 97928 25504 97980
rect 25556 97968 25562 97980
rect 129458 97968 129464 97980
rect 25556 97940 129464 97968
rect 25556 97928 25562 97940
rect 129458 97928 129464 97940
rect 129516 97928 129522 97980
rect 146754 97928 146760 97980
rect 146812 97968 146818 97980
rect 567838 97968 567844 97980
rect 146812 97940 567844 97968
rect 146812 97928 146818 97940
rect 567838 97928 567844 97940
rect 567896 97928 567902 97980
rect 43438 97860 43444 97912
rect 43496 97900 43502 97912
rect 346762 97900 346768 97912
rect 43496 97872 346768 97900
rect 43496 97860 43502 97872
rect 346762 97860 346768 97872
rect 346820 97860 346826 97912
rect 69842 97792 69848 97844
rect 69900 97832 69906 97844
rect 178770 97832 178776 97844
rect 69900 97804 178776 97832
rect 69900 97792 69906 97804
rect 178770 97792 178776 97804
rect 178828 97792 178834 97844
rect 491294 97588 491300 97640
rect 491352 97628 491358 97640
rect 503070 97628 503076 97640
rect 491352 97600 503076 97628
rect 491352 97588 491358 97600
rect 503070 97588 503076 97600
rect 503128 97588 503134 97640
rect 487798 97520 487804 97572
rect 487856 97560 487862 97572
rect 523218 97560 523224 97572
rect 487856 97532 523224 97560
rect 487856 97520 487862 97532
rect 523218 97520 523224 97532
rect 523276 97520 523282 97572
rect 463602 97452 463608 97504
rect 463660 97492 463666 97504
rect 505370 97492 505376 97504
rect 463660 97464 505376 97492
rect 463660 97452 463666 97464
rect 505370 97452 505376 97464
rect 505428 97452 505434 97504
rect 61838 97384 61844 97436
rect 61896 97424 61902 97436
rect 81894 97424 81900 97436
rect 61896 97396 81900 97424
rect 61896 97384 61902 97396
rect 81894 97384 81900 97396
rect 81952 97384 81958 97436
rect 365622 97384 365628 97436
rect 365680 97424 365686 97436
rect 517790 97424 517796 97436
rect 365680 97396 517796 97424
rect 365680 97384 365686 97396
rect 517790 97384 517796 97396
rect 517848 97384 517854 97436
rect 57882 97316 57888 97368
rect 57940 97356 57946 97368
rect 81434 97356 81440 97368
rect 57940 97328 81440 97356
rect 57940 97316 57946 97328
rect 81434 97316 81440 97328
rect 81492 97316 81498 97368
rect 355962 97316 355968 97368
rect 356020 97356 356026 97368
rect 520550 97356 520556 97368
rect 356020 97328 520556 97356
rect 356020 97316 356026 97328
rect 520550 97316 520556 97328
rect 520608 97316 520614 97368
rect 79778 97248 79784 97300
rect 79836 97288 79842 97300
rect 212534 97288 212540 97300
rect 79836 97260 212540 97288
rect 79836 97248 79842 97260
rect 212534 97248 212540 97260
rect 212592 97248 212598 97300
rect 329742 97248 329748 97300
rect 329800 97288 329806 97300
rect 516410 97288 516416 97300
rect 329800 97260 516416 97288
rect 329800 97248 329806 97260
rect 516410 97248 516416 97260
rect 516468 97248 516474 97300
rect 212258 96636 212264 96688
rect 212316 96676 212322 96688
rect 212350 96676 212356 96688
rect 212316 96648 212356 96676
rect 212316 96636 212322 96648
rect 212350 96636 212356 96648
rect 212408 96636 212414 96688
rect 356514 96676 356520 96688
rect 356475 96648 356520 96676
rect 356514 96636 356520 96648
rect 356572 96636 356578 96688
rect 168834 96568 168840 96620
rect 168892 96608 168898 96620
rect 176657 96611 176715 96617
rect 176657 96608 176669 96611
rect 168892 96580 176669 96608
rect 168892 96568 168898 96580
rect 176657 96577 176669 96580
rect 176703 96577 176715 96611
rect 176657 96571 176715 96577
rect 176746 96568 176752 96620
rect 176804 96568 176810 96620
rect 176841 96611 176899 96617
rect 176841 96577 176853 96611
rect 176887 96608 176899 96611
rect 212169 96611 212227 96617
rect 212169 96608 212181 96611
rect 176887 96580 212181 96608
rect 176887 96577 176899 96580
rect 176841 96571 176899 96577
rect 212169 96577 212181 96580
rect 212215 96577 212227 96611
rect 212169 96571 212227 96577
rect 212445 96611 212503 96617
rect 212445 96577 212457 96611
rect 212491 96608 212503 96611
rect 356425 96611 356483 96617
rect 356425 96608 356437 96611
rect 212491 96580 356437 96608
rect 212491 96577 212503 96580
rect 212445 96571 212503 96577
rect 356425 96577 356437 96580
rect 356471 96577 356483 96611
rect 356425 96571 356483 96577
rect 356609 96611 356667 96617
rect 356609 96577 356621 96611
rect 356655 96608 356667 96611
rect 512733 96611 512791 96617
rect 512733 96608 512745 96611
rect 356655 96580 512745 96608
rect 356655 96577 356667 96580
rect 356609 96571 356667 96577
rect 512733 96577 512745 96580
rect 512779 96577 512791 96611
rect 512733 96571 512791 96577
rect 512917 96611 512975 96617
rect 512917 96577 512929 96611
rect 512963 96608 512975 96611
rect 565078 96608 565084 96620
rect 512963 96580 565084 96608
rect 512963 96577 512975 96580
rect 512917 96571 512975 96577
rect 565078 96568 565084 96580
rect 565136 96568 565142 96620
rect 32398 96500 32404 96552
rect 32456 96540 32462 96552
rect 176565 96543 176623 96549
rect 176565 96540 176577 96543
rect 32456 96512 176577 96540
rect 32456 96500 32462 96512
rect 176565 96509 176577 96512
rect 176611 96509 176623 96543
rect 176565 96503 176623 96509
rect 176764 96481 176792 96568
rect 176933 96543 176991 96549
rect 176933 96509 176945 96543
rect 176979 96540 176991 96543
rect 356333 96543 356391 96549
rect 356333 96540 356345 96543
rect 176979 96512 356345 96540
rect 176979 96509 176991 96512
rect 176933 96503 176991 96509
rect 356333 96509 356345 96512
rect 356379 96509 356391 96543
rect 356333 96503 356391 96509
rect 356701 96543 356759 96549
rect 356701 96509 356713 96543
rect 356747 96540 356759 96543
rect 413554 96540 413560 96552
rect 356747 96512 413560 96540
rect 356747 96509 356759 96512
rect 356701 96503 356759 96509
rect 413554 96500 413560 96512
rect 413612 96500 413618 96552
rect 456610 96500 456616 96552
rect 456668 96540 456674 96552
rect 512549 96543 512607 96549
rect 512549 96540 512561 96543
rect 456668 96512 512561 96540
rect 456668 96500 456674 96512
rect 512549 96509 512561 96512
rect 512595 96509 512607 96543
rect 512549 96503 512607 96509
rect 176749 96475 176807 96481
rect 176749 96441 176761 96475
rect 176795 96441 176807 96475
rect 176749 96435 176807 96441
rect 191098 96432 191104 96484
rect 191156 96472 191162 96484
rect 212353 96475 212411 96481
rect 212353 96472 212365 96475
rect 191156 96444 212365 96472
rect 191156 96432 191162 96444
rect 212353 96441 212365 96444
rect 212399 96441 212411 96475
rect 212353 96435 212411 96441
rect 212445 96475 212503 96481
rect 212445 96441 212457 96475
rect 212491 96472 212503 96475
rect 512638 96472 512644 96484
rect 212491 96444 347820 96472
rect 212491 96441 212503 96444
rect 212445 96435 212503 96441
rect 347792 96404 347820 96444
rect 356624 96444 512644 96472
rect 356624 96404 356652 96444
rect 512638 96432 512644 96444
rect 512696 96432 512702 96484
rect 347792 96376 356652 96404
rect 440142 96364 440148 96416
rect 440200 96404 440206 96416
rect 516318 96404 516324 96416
rect 440200 96376 516324 96404
rect 440200 96364 440206 96376
rect 516318 96364 516324 96376
rect 516376 96364 516382 96416
rect 398742 96296 398748 96348
rect 398800 96336 398806 96348
rect 501782 96336 501788 96348
rect 398800 96308 501788 96336
rect 398800 96296 398806 96308
rect 501782 96296 501788 96308
rect 501840 96296 501846 96348
rect 512549 96339 512607 96345
rect 512549 96305 512561 96339
rect 512595 96336 512607 96339
rect 519262 96336 519268 96348
rect 512595 96308 519268 96336
rect 512595 96305 512607 96308
rect 512549 96299 512607 96305
rect 519262 96296 519268 96308
rect 519320 96296 519326 96348
rect 389082 96228 389088 96280
rect 389140 96268 389146 96280
rect 510982 96268 510988 96280
rect 389140 96240 510988 96268
rect 389140 96228 389146 96240
rect 510982 96228 510988 96240
rect 511040 96228 511046 96280
rect 349062 96160 349068 96212
rect 349120 96200 349126 96212
rect 508406 96200 508412 96212
rect 349120 96172 508412 96200
rect 349120 96160 349126 96172
rect 508406 96160 508412 96172
rect 508464 96160 508470 96212
rect 326982 96092 326988 96144
rect 327040 96132 327046 96144
rect 515030 96132 515036 96144
rect 327040 96104 515036 96132
rect 327040 96092 327046 96104
rect 515030 96092 515036 96104
rect 515088 96092 515094 96144
rect 275922 96024 275928 96076
rect 275980 96064 275986 96076
rect 510706 96064 510712 96076
rect 275980 96036 510712 96064
rect 275980 96024 275986 96036
rect 510706 96024 510712 96036
rect 510764 96024 510770 96076
rect 195882 95956 195888 96008
rect 195940 95996 195946 96008
rect 516502 95996 516508 96008
rect 195940 95968 516508 95996
rect 195940 95956 195946 95968
rect 516502 95956 516508 95968
rect 516560 95956 516566 96008
rect 83277 95931 83335 95937
rect 83277 95897 83289 95931
rect 83323 95928 83335 95931
rect 83366 95928 83372 95940
rect 83323 95900 83372 95928
rect 83323 95897 83335 95900
rect 83277 95891 83335 95897
rect 83366 95888 83372 95900
rect 83424 95888 83430 95940
rect 151722 95888 151728 95940
rect 151780 95928 151786 95940
rect 520826 95928 520832 95940
rect 151780 95900 520832 95928
rect 151780 95888 151786 95900
rect 520826 95888 520832 95900
rect 520884 95888 520890 95940
rect 512641 95251 512699 95257
rect 512641 95217 512653 95251
rect 512687 95248 512699 95251
rect 512730 95248 512736 95260
rect 512687 95220 512736 95248
rect 512687 95217 512699 95220
rect 512641 95211 512699 95217
rect 512730 95208 512736 95220
rect 512788 95208 512794 95260
rect 484210 95004 484216 95056
rect 484268 95044 484274 95056
rect 487798 95044 487804 95056
rect 484268 95016 487804 95044
rect 484268 95004 484274 95016
rect 487798 95004 487804 95016
rect 487856 95004 487862 95056
rect 481726 94936 481732 94988
rect 481784 94976 481790 94988
rect 484486 94976 484492 94988
rect 481784 94948 484492 94976
rect 481784 94936 481790 94948
rect 484486 94936 484492 94948
rect 484544 94936 484550 94988
rect 86957 94843 87015 94849
rect 86957 94809 86969 94843
rect 87003 94840 87015 94843
rect 96525 94843 96583 94849
rect 96525 94840 96537 94843
rect 87003 94812 96537 94840
rect 87003 94809 87015 94812
rect 86957 94803 87015 94809
rect 96525 94809 96537 94812
rect 96571 94809 96583 94843
rect 96525 94803 96583 94809
rect 83458 94664 83464 94716
rect 83516 94704 83522 94716
rect 86957 94707 87015 94713
rect 86957 94704 86969 94707
rect 83516 94676 86969 94704
rect 83516 94664 83522 94676
rect 86957 94673 86969 94676
rect 87003 94673 87015 94707
rect 86957 94667 87015 94673
rect 492766 94664 492772 94716
rect 492824 94704 492830 94716
rect 523126 94704 523132 94716
rect 492824 94676 523132 94704
rect 492824 94664 492830 94676
rect 523126 94664 523132 94676
rect 523184 94664 523190 94716
rect 115937 94639 115995 94645
rect 115937 94605 115949 94639
rect 115983 94605 115995 94639
rect 115937 94599 115995 94605
rect 83090 94528 83096 94580
rect 83148 94568 83154 94580
rect 83458 94568 83464 94580
rect 83148 94540 83464 94568
rect 83148 94528 83154 94540
rect 83458 94528 83464 94540
rect 83516 94528 83522 94580
rect 96525 94571 96583 94577
rect 96525 94537 96537 94571
rect 96571 94568 96583 94571
rect 115952 94568 115980 94599
rect 393222 94596 393228 94648
rect 393280 94636 393286 94648
rect 505554 94636 505560 94648
rect 393280 94608 505560 94636
rect 393280 94596 393286 94608
rect 505554 94596 505560 94608
rect 505612 94596 505618 94648
rect 96571 94540 115980 94568
rect 96571 94537 96583 94540
rect 96525 94531 96583 94537
rect 367002 94528 367008 94580
rect 367060 94568 367066 94580
rect 501598 94568 501604 94580
rect 367060 94540 501604 94568
rect 367060 94528 367066 94540
rect 501598 94528 501604 94540
rect 501656 94528 501662 94580
rect 79134 94460 79140 94512
rect 79192 94500 79198 94512
rect 567194 94500 567200 94512
rect 79192 94472 567200 94500
rect 79192 94460 79198 94472
rect 567194 94460 567200 94472
rect 567252 94460 567258 94512
rect 487798 93848 487804 93900
rect 487856 93888 487862 93900
rect 491294 93888 491300 93900
rect 487856 93860 491300 93888
rect 487856 93848 487862 93860
rect 491294 93848 491300 93860
rect 491352 93848 491358 93900
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 15930 93820 15936 93832
rect 3476 93792 15936 93820
rect 3476 93780 3482 93792
rect 15930 93780 15936 93792
rect 15988 93780 15994 93832
rect 433242 93712 433248 93764
rect 433300 93752 433306 93764
rect 507118 93752 507124 93764
rect 433300 93724 507124 93752
rect 433300 93712 433306 93724
rect 507118 93712 507124 93724
rect 507176 93712 507182 93764
rect 411165 93687 411223 93693
rect 411165 93653 411177 93687
rect 411211 93684 411223 93687
rect 522114 93684 522120 93696
rect 411211 93656 522120 93684
rect 411211 93653 411223 93656
rect 411165 93647 411223 93653
rect 522114 93644 522120 93656
rect 522172 93644 522178 93696
rect 386322 93576 386328 93628
rect 386380 93616 386386 93628
rect 521746 93616 521752 93628
rect 386380 93588 521752 93616
rect 386380 93576 386386 93588
rect 521746 93576 521752 93588
rect 521804 93576 521810 93628
rect 249702 93508 249708 93560
rect 249760 93548 249766 93560
rect 516686 93548 516692 93560
rect 249760 93520 516692 93548
rect 249760 93508 249766 93520
rect 516686 93508 516692 93520
rect 516744 93508 516750 93560
rect 220722 93440 220728 93492
rect 220780 93480 220786 93492
rect 505186 93480 505192 93492
rect 220780 93452 505192 93480
rect 220780 93440 220786 93452
rect 505186 93440 505192 93452
rect 505244 93440 505250 93492
rect 217962 93372 217968 93424
rect 218020 93412 218026 93424
rect 521930 93412 521936 93424
rect 218020 93384 521936 93412
rect 218020 93372 218026 93384
rect 521930 93372 521936 93384
rect 521988 93372 521994 93424
rect 173802 93304 173808 93356
rect 173860 93344 173866 93356
rect 196066 93344 196072 93356
rect 173860 93316 196072 93344
rect 173860 93304 173866 93316
rect 196066 93304 196072 93316
rect 196124 93304 196130 93356
rect 200022 93304 200028 93356
rect 200080 93344 200086 93356
rect 520734 93344 520740 93356
rect 200080 93316 520740 93344
rect 200080 93304 200086 93316
rect 520734 93304 520740 93316
rect 520792 93304 520798 93356
rect 115937 93279 115995 93285
rect 115937 93245 115949 93279
rect 115983 93276 115995 93279
rect 122834 93276 122840 93288
rect 115983 93248 122840 93276
rect 115983 93245 115995 93248
rect 115937 93239 115995 93245
rect 122834 93236 122840 93248
rect 122892 93236 122898 93288
rect 186222 93236 186228 93288
rect 186280 93276 186286 93288
rect 515306 93276 515312 93288
rect 186280 93248 515312 93276
rect 186280 93236 186286 93248
rect 515306 93236 515312 93248
rect 515364 93236 515370 93288
rect 183462 93168 183468 93220
rect 183520 93208 183526 93220
rect 518066 93208 518072 93220
rect 183520 93180 518072 93208
rect 183520 93168 183526 93180
rect 518066 93168 518072 93180
rect 518124 93168 518130 93220
rect 59262 93100 59268 93152
rect 59320 93140 59326 93152
rect 78674 93140 78680 93152
rect 59320 93112 78680 93140
rect 59320 93100 59326 93112
rect 78674 93100 78680 93112
rect 78732 93100 78738 93152
rect 146202 93100 146208 93152
rect 146260 93140 146266 93152
rect 522022 93140 522028 93152
rect 146260 93112 522028 93140
rect 146260 93100 146266 93112
rect 522022 93100 522028 93112
rect 522080 93100 522086 93152
rect 488534 91944 488540 91996
rect 488592 91984 488598 91996
rect 492766 91984 492772 91996
rect 488592 91956 492772 91984
rect 488592 91944 488598 91956
rect 492766 91944 492772 91956
rect 492824 91944 492830 91996
rect 436002 91876 436008 91928
rect 436060 91916 436066 91928
rect 507946 91916 507952 91928
rect 436060 91888 507952 91916
rect 436060 91876 436066 91888
rect 507946 91876 507952 91888
rect 508004 91876 508010 91928
rect 278682 91808 278688 91860
rect 278740 91848 278746 91860
rect 505094 91848 505100 91860
rect 278740 91820 505100 91848
rect 278740 91808 278746 91820
rect 505094 91808 505100 91820
rect 505152 91808 505158 91860
rect 79410 91740 79416 91792
rect 79468 91780 79474 91792
rect 444374 91780 444380 91792
rect 79468 91752 444380 91780
rect 79468 91740 79474 91752
rect 444374 91740 444380 91752
rect 444432 91740 444438 91792
rect 480714 91060 480720 91112
rect 480772 91100 480778 91112
rect 481726 91100 481732 91112
rect 480772 91072 481732 91100
rect 480772 91060 480778 91072
rect 481726 91060 481732 91072
rect 481784 91060 481790 91112
rect 483014 91060 483020 91112
rect 483072 91100 483078 91112
rect 488626 91100 488632 91112
rect 483072 91072 488632 91100
rect 483072 91060 483078 91072
rect 488626 91060 488632 91072
rect 488684 91060 488690 91112
rect 298002 90380 298008 90432
rect 298060 90420 298066 90432
rect 519354 90420 519360 90432
rect 298060 90392 519360 90420
rect 298060 90380 298066 90392
rect 519354 90380 519360 90392
rect 519412 90380 519418 90432
rect 76650 90312 76656 90364
rect 76708 90352 76714 90364
rect 335354 90352 335360 90364
rect 76708 90324 335360 90352
rect 76708 90312 76714 90324
rect 335354 90312 335360 90324
rect 335412 90312 335418 90364
rect 356514 89700 356520 89752
rect 356572 89700 356578 89752
rect 176746 89672 176752 89684
rect 176707 89644 176752 89672
rect 176746 89632 176752 89644
rect 176804 89632 176810 89684
rect 356532 89604 356560 89700
rect 356606 89604 356612 89616
rect 356532 89576 356612 89604
rect 356606 89564 356612 89576
rect 356664 89564 356670 89616
rect 83274 89400 83280 89412
rect 83235 89372 83280 89400
rect 83274 89360 83280 89372
rect 83332 89360 83338 89412
rect 78122 89020 78128 89072
rect 78180 89060 78186 89072
rect 304994 89060 305000 89072
rect 78180 89032 305000 89060
rect 78180 89020 78186 89032
rect 304994 89020 305000 89032
rect 305052 89020 305058 89072
rect 280062 88952 280068 89004
rect 280120 88992 280126 89004
rect 508038 88992 508044 89004
rect 280120 88964 508044 88992
rect 280120 88952 280126 88964
rect 508038 88952 508044 88964
rect 508096 88952 508102 89004
rect 484486 88612 484492 88664
rect 484544 88652 484550 88664
rect 487798 88652 487804 88664
rect 484544 88624 487804 88652
rect 484544 88612 484550 88624
rect 487798 88612 487804 88624
rect 487856 88612 487862 88664
rect 482278 88476 482284 88528
rect 482336 88516 482342 88528
rect 484210 88516 484216 88528
rect 482336 88488 484216 88516
rect 482336 88476 482342 88488
rect 484210 88476 484216 88488
rect 484268 88476 484274 88528
rect 84930 87592 84936 87644
rect 84988 87632 84994 87644
rect 138014 87632 138020 87644
rect 84988 87604 138020 87632
rect 84988 87592 84994 87604
rect 138014 87592 138020 87604
rect 138072 87592 138078 87644
rect 176470 87592 176476 87644
rect 176528 87632 176534 87644
rect 187694 87632 187700 87644
rect 176528 87604 187700 87632
rect 176528 87592 176534 87604
rect 187694 87592 187700 87604
rect 187752 87592 187758 87644
rect 293862 87592 293868 87644
rect 293920 87632 293926 87644
rect 506750 87632 506756 87644
rect 293920 87604 506756 87632
rect 293920 87592 293926 87604
rect 506750 87592 506756 87604
rect 506808 87592 506814 87644
rect 151538 86980 151544 87032
rect 151596 87020 151602 87032
rect 151630 87020 151636 87032
rect 151596 86992 151636 87020
rect 151596 86980 151602 86992
rect 151630 86980 151636 86992
rect 151688 86980 151694 87032
rect 411162 87020 411168 87032
rect 411123 86992 411168 87020
rect 411162 86980 411168 86992
rect 411220 86980 411226 87032
rect 512730 86980 512736 87032
rect 512788 87020 512794 87032
rect 512822 87020 512828 87032
rect 512788 86992 512828 87020
rect 512788 86980 512794 86992
rect 512822 86980 512828 86992
rect 512880 86980 512886 87032
rect 176654 86912 176660 86964
rect 176712 86952 176718 86964
rect 176746 86952 176752 86964
rect 176712 86924 176752 86952
rect 176712 86912 176718 86924
rect 176746 86912 176752 86924
rect 176804 86912 176810 86964
rect 198461 86955 198519 86961
rect 198461 86921 198473 86955
rect 198507 86952 198519 86955
rect 198550 86952 198556 86964
rect 198507 86924 198556 86952
rect 198507 86921 198519 86924
rect 198461 86915 198519 86921
rect 198550 86912 198556 86924
rect 198608 86912 198614 86964
rect 280433 86955 280491 86961
rect 280433 86921 280445 86955
rect 280479 86952 280491 86955
rect 280522 86952 280528 86964
rect 280479 86924 280528 86952
rect 280479 86921 280491 86924
rect 280433 86915 280491 86921
rect 280522 86912 280528 86924
rect 280580 86912 280586 86964
rect 483750 86912 483756 86964
rect 483808 86952 483814 86964
rect 484486 86952 484492 86964
rect 483808 86924 484492 86952
rect 483808 86912 483814 86924
rect 484486 86912 484492 86924
rect 484544 86912 484550 86964
rect 487246 86640 487252 86692
rect 487304 86680 487310 86692
rect 488534 86680 488540 86692
rect 487304 86652 488540 86680
rect 487304 86640 487310 86652
rect 488534 86640 488540 86652
rect 488592 86640 488598 86692
rect 201402 86368 201408 86420
rect 201460 86408 201466 86420
rect 274634 86408 274640 86420
rect 201460 86380 274640 86408
rect 201460 86368 201466 86380
rect 274634 86368 274640 86380
rect 274692 86368 274698 86420
rect 253842 86300 253848 86352
rect 253900 86340 253906 86352
rect 504266 86340 504272 86352
rect 253900 86312 504272 86340
rect 253900 86300 253906 86312
rect 504266 86300 504272 86312
rect 504324 86300 504330 86352
rect 75454 86232 75460 86284
rect 75512 86272 75518 86284
rect 342254 86272 342260 86284
rect 75512 86244 342260 86272
rect 75512 86232 75518 86244
rect 342254 86232 342260 86244
rect 342312 86232 342318 86284
rect 473262 86232 473268 86284
rect 473320 86272 473326 86284
rect 528554 86272 528560 86284
rect 473320 86244 528560 86272
rect 473320 86232 473326 86244
rect 528554 86232 528560 86244
rect 528612 86232 528618 86284
rect 477494 85552 477500 85604
rect 477552 85592 477558 85604
rect 480714 85592 480720 85604
rect 477552 85564 480720 85592
rect 477552 85552 477558 85564
rect 480714 85552 480720 85564
rect 480772 85552 480778 85604
rect 79778 85524 79784 85536
rect 79739 85496 79784 85524
rect 79778 85484 79784 85496
rect 79836 85484 79842 85536
rect 512822 85524 512828 85536
rect 512783 85496 512828 85524
rect 512822 85484 512828 85496
rect 512880 85484 512886 85536
rect 558178 85484 558184 85536
rect 558236 85524 558242 85536
rect 564434 85524 564440 85536
rect 558236 85496 564440 85524
rect 558236 85484 558242 85496
rect 564434 85484 564440 85496
rect 564492 85484 564498 85536
rect 77018 84872 77024 84924
rect 77076 84912 77082 84924
rect 155954 84912 155960 84924
rect 77076 84884 155960 84912
rect 77076 84872 77082 84884
rect 155954 84872 155960 84884
rect 156012 84872 156018 84924
rect 102042 84804 102048 84856
rect 102100 84844 102106 84856
rect 261478 84844 261484 84856
rect 102100 84816 261484 84844
rect 102100 84804 102106 84816
rect 261478 84804 261484 84816
rect 261536 84804 261542 84856
rect 314562 84804 314568 84856
rect 314620 84844 314626 84856
rect 508222 84844 508228 84856
rect 314620 84816 508228 84844
rect 314620 84804 314626 84816
rect 508222 84804 508228 84816
rect 508280 84804 508286 84856
rect 482922 84232 482928 84244
rect 478892 84204 482928 84232
rect 476114 84124 476120 84176
rect 476172 84164 476178 84176
rect 478892 84164 478920 84204
rect 482922 84192 482928 84204
rect 482980 84192 482986 84244
rect 476172 84136 478920 84164
rect 476172 84124 476178 84136
rect 78214 83580 78220 83632
rect 78272 83620 78278 83632
rect 287054 83620 287060 83632
rect 78272 83592 287060 83620
rect 78272 83580 78278 83592
rect 287054 83580 287060 83592
rect 287112 83580 287118 83632
rect 210878 83512 210884 83564
rect 210936 83552 210942 83564
rect 502702 83552 502708 83564
rect 210936 83524 502708 83552
rect 210936 83512 210942 83524
rect 502702 83512 502708 83524
rect 502760 83512 502766 83564
rect 79226 83444 79232 83496
rect 79284 83484 79290 83496
rect 451274 83484 451280 83496
rect 79284 83456 451280 83484
rect 79284 83444 79290 83456
rect 451274 83444 451280 83456
rect 451332 83444 451338 83496
rect 481082 82832 481088 82884
rect 481140 82872 481146 82884
rect 483750 82872 483756 82884
rect 481140 82844 483756 82872
rect 481140 82832 481146 82844
rect 483750 82832 483756 82844
rect 483808 82832 483814 82884
rect 485498 82832 485504 82884
rect 485556 82872 485562 82884
rect 487246 82872 487252 82884
rect 485556 82844 487252 82872
rect 485556 82832 485562 82844
rect 487246 82832 487252 82844
rect 487304 82832 487310 82884
rect 89898 82084 89904 82136
rect 89956 82124 89962 82136
rect 90082 82124 90088 82136
rect 89956 82096 90088 82124
rect 89956 82084 89962 82096
rect 90082 82084 90088 82096
rect 90140 82084 90146 82136
rect 211062 82084 211068 82136
rect 211120 82124 211126 82136
rect 396074 82124 396080 82136
rect 211120 82096 396080 82124
rect 211120 82084 211126 82096
rect 396074 82084 396080 82096
rect 396132 82084 396138 82136
rect 478874 81404 478880 81456
rect 478932 81444 478938 81456
rect 481082 81444 481088 81456
rect 478932 81416 481088 81444
rect 478932 81404 478938 81416
rect 481082 81404 481088 81416
rect 481140 81404 481146 81456
rect 151538 81104 151544 81116
rect 151499 81076 151544 81104
rect 151538 81064 151544 81076
rect 151596 81064 151602 81116
rect 228910 80656 228916 80708
rect 228968 80696 228974 80708
rect 505462 80696 505468 80708
rect 228968 80668 505468 80696
rect 228968 80656 228974 80668
rect 505462 80656 505468 80668
rect 505520 80656 505526 80708
rect 356606 80044 356612 80096
rect 356664 80044 356670 80096
rect 474642 80044 474648 80096
rect 474700 80084 474706 80096
rect 476114 80084 476120 80096
rect 474700 80056 476120 80084
rect 474700 80044 474706 80056
rect 476114 80044 476120 80056
rect 476172 80044 476178 80096
rect 356624 79948 356652 80044
rect 356698 79948 356704 79960
rect 356624 79920 356704 79948
rect 356698 79908 356704 79920
rect 356756 79908 356762 79960
rect 271782 79364 271788 79416
rect 271840 79404 271846 79416
rect 506474 79404 506480 79416
rect 271840 79376 506480 79404
rect 271840 79364 271846 79376
rect 506474 79364 506480 79376
rect 506532 79364 506538 79416
rect 76834 79296 76840 79348
rect 76892 79336 76898 79348
rect 378134 79336 378140 79348
rect 76892 79308 378140 79336
rect 76892 79296 76898 79308
rect 378134 79296 378140 79308
rect 378192 79296 378198 79348
rect 473262 79296 473268 79348
rect 473320 79336 473326 79348
rect 477402 79336 477408 79348
rect 473320 79308 477408 79336
rect 473320 79296 473326 79308
rect 477402 79296 477408 79308
rect 477460 79296 477466 79348
rect 483658 78208 483664 78260
rect 483716 78248 483722 78260
rect 485498 78248 485504 78260
rect 483716 78220 485504 78248
rect 483716 78208 483722 78220
rect 485498 78208 485504 78220
rect 485556 78208 485562 78260
rect 75362 78072 75368 78124
rect 75420 78112 75426 78124
rect 263594 78112 263600 78124
rect 75420 78084 263600 78112
rect 75420 78072 75426 78084
rect 263594 78072 263600 78084
rect 263652 78072 263658 78124
rect 471238 78072 471244 78124
rect 471296 78112 471302 78124
rect 474642 78112 474648 78124
rect 471296 78084 474648 78112
rect 471296 78072 471302 78084
rect 474642 78072 474648 78084
rect 474700 78072 474706 78124
rect 157242 78004 157248 78056
rect 157300 78044 157306 78056
rect 230474 78044 230480 78056
rect 157300 78016 230480 78044
rect 157300 78004 157306 78016
rect 230474 78004 230480 78016
rect 230532 78004 230538 78056
rect 245562 78004 245568 78056
rect 245620 78044 245626 78056
rect 501874 78044 501880 78056
rect 245620 78016 501880 78044
rect 245620 78004 245626 78016
rect 501874 78004 501880 78016
rect 501932 78004 501938 78056
rect 194502 77936 194508 77988
rect 194560 77976 194566 77988
rect 481634 77976 481640 77988
rect 194560 77948 481640 77976
rect 194560 77936 194566 77948
rect 481634 77936 481640 77948
rect 481692 77936 481698 77988
rect 475378 77528 475384 77580
rect 475436 77568 475442 77580
rect 478874 77568 478880 77580
rect 475436 77540 478880 77568
rect 475436 77528 475442 77540
rect 478874 77528 478880 77540
rect 478932 77528 478938 77580
rect 151538 77364 151544 77376
rect 151499 77336 151544 77364
rect 151538 77324 151544 77336
rect 151596 77324 151602 77376
rect 198458 77296 198464 77308
rect 198419 77268 198464 77296
rect 198458 77256 198464 77268
rect 198516 77256 198522 77308
rect 280430 77296 280436 77308
rect 280391 77268 280436 77296
rect 280430 77256 280436 77268
rect 280488 77256 280494 77308
rect 72510 77188 72516 77240
rect 72568 77228 72574 77240
rect 212353 77231 212411 77237
rect 212353 77228 212365 77231
rect 72568 77200 212365 77228
rect 72568 77188 72574 77200
rect 212353 77197 212365 77200
rect 212399 77197 212411 77231
rect 212353 77191 212411 77197
rect 212445 77231 212503 77237
rect 212445 77197 212457 77231
rect 212491 77228 212503 77231
rect 580166 77228 580172 77240
rect 212491 77200 580172 77228
rect 212491 77197 212503 77200
rect 212445 77191 212503 77197
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 151446 77160 151452 77172
rect 151407 77132 151452 77160
rect 151446 77120 151452 77132
rect 151504 77120 151510 77172
rect 176749 77163 176807 77169
rect 176749 77129 176761 77163
rect 176795 77160 176807 77163
rect 176838 77160 176844 77172
rect 176795 77132 176844 77160
rect 176795 77129 176807 77132
rect 176749 77123 176807 77129
rect 176838 77120 176844 77132
rect 176896 77120 176902 77172
rect 198458 77160 198464 77172
rect 198419 77132 198464 77160
rect 198458 77120 198464 77132
rect 198516 77120 198522 77172
rect 356698 77160 356704 77172
rect 356659 77132 356704 77160
rect 356698 77120 356704 77132
rect 356756 77120 356762 77172
rect 411162 77160 411168 77172
rect 411123 77132 411168 77160
rect 411162 77120 411168 77132
rect 411220 77120 411226 77172
rect 470594 76712 470600 76764
rect 470652 76752 470658 76764
rect 473262 76752 473268 76764
rect 470652 76724 473268 76752
rect 470652 76712 470658 76724
rect 473262 76712 473268 76724
rect 473320 76712 473326 76764
rect 85482 76576 85488 76628
rect 85540 76616 85546 76628
rect 242894 76616 242900 76628
rect 85540 76588 242900 76616
rect 85540 76576 85546 76588
rect 242894 76576 242900 76588
rect 242952 76576 242958 76628
rect 184842 76508 184848 76560
rect 184900 76548 184906 76560
rect 360194 76548 360200 76560
rect 184900 76520 360200 76548
rect 184900 76508 184906 76520
rect 360194 76508 360200 76520
rect 360252 76508 360258 76560
rect 79781 75939 79839 75945
rect 79781 75905 79793 75939
rect 79827 75936 79839 75939
rect 79962 75936 79968 75948
rect 79827 75908 79968 75936
rect 79827 75905 79839 75908
rect 79781 75899 79839 75905
rect 79962 75896 79968 75908
rect 80020 75896 80026 75948
rect 512822 75936 512828 75948
rect 512783 75908 512828 75936
rect 512822 75896 512828 75908
rect 512880 75896 512886 75948
rect 480898 75828 480904 75880
rect 480956 75868 480962 75880
rect 482278 75868 482284 75880
rect 480956 75840 482284 75868
rect 480956 75828 480962 75840
rect 482278 75828 482284 75840
rect 482336 75828 482342 75880
rect 119982 75148 119988 75200
rect 120040 75188 120046 75200
rect 204254 75188 204260 75200
rect 120040 75160 204260 75188
rect 120040 75148 120046 75160
rect 204254 75148 204260 75160
rect 204312 75148 204318 75200
rect 233142 75148 233148 75200
rect 233200 75188 233206 75200
rect 309226 75188 309232 75200
rect 233200 75160 309232 75188
rect 233200 75148 233206 75160
rect 309226 75148 309232 75160
rect 309284 75148 309290 75200
rect 107562 73924 107568 73976
rect 107620 73964 107626 73976
rect 133874 73964 133880 73976
rect 107620 73936 133880 73964
rect 107620 73924 107626 73936
rect 133874 73924 133880 73936
rect 133932 73924 133938 73976
rect 240042 73924 240048 73976
rect 240100 73964 240106 73976
rect 385034 73964 385040 73976
rect 240100 73936 385040 73964
rect 240100 73924 240106 73936
rect 385034 73924 385040 73936
rect 385092 73924 385098 73976
rect 76558 73856 76564 73908
rect 76616 73896 76622 73908
rect 171134 73896 171140 73908
rect 76616 73868 171140 73896
rect 76616 73856 76622 73868
rect 171134 73856 171140 73868
rect 171192 73856 171198 73908
rect 332502 73856 332508 73908
rect 332560 73896 332566 73908
rect 501690 73896 501696 73908
rect 332560 73868 501696 73896
rect 332560 73856 332566 73868
rect 501690 73856 501696 73868
rect 501748 73856 501754 73908
rect 19242 73788 19248 73840
rect 19300 73828 19306 73840
rect 338114 73828 338120 73840
rect 19300 73800 338120 73828
rect 19300 73788 19306 73800
rect 338114 73788 338120 73800
rect 338172 73788 338178 73840
rect 342162 72496 342168 72548
rect 342220 72536 342226 72548
rect 489914 72536 489920 72548
rect 342220 72508 489920 72536
rect 342220 72496 342226 72508
rect 489914 72496 489920 72508
rect 489972 72496 489978 72548
rect 84010 72428 84016 72480
rect 84068 72468 84074 72480
rect 553394 72468 553400 72480
rect 84068 72440 553400 72468
rect 84068 72428 84074 72440
rect 553394 72428 553400 72440
rect 553452 72428 553458 72480
rect 469306 71952 469312 72004
rect 469364 71992 469370 72004
rect 471238 71992 471244 72004
rect 469364 71964 471244 71992
rect 469364 71952 469370 71964
rect 471238 71952 471244 71964
rect 471296 71952 471302 72004
rect 226242 71068 226248 71120
rect 226300 71108 226306 71120
rect 284294 71108 284300 71120
rect 226300 71080 284300 71108
rect 226300 71068 226306 71080
rect 284294 71068 284300 71080
rect 284352 71068 284358 71120
rect 364150 71068 364156 71120
rect 364208 71108 364214 71120
rect 371234 71108 371240 71120
rect 364208 71080 371240 71108
rect 364208 71068 364214 71080
rect 371234 71068 371240 71080
rect 371292 71068 371298 71120
rect 93762 71000 93768 71052
rect 93820 71040 93826 71052
rect 365714 71040 365720 71052
rect 93820 71012 365720 71040
rect 93820 71000 93826 71012
rect 365714 71000 365720 71012
rect 365772 71000 365778 71052
rect 375190 71000 375196 71052
rect 375248 71040 375254 71052
rect 418154 71040 418160 71052
rect 375248 71012 418160 71040
rect 375248 71000 375254 71012
rect 418154 71000 418160 71012
rect 418212 71000 418218 71052
rect 472434 70592 472440 70644
rect 472492 70632 472498 70644
rect 475378 70632 475384 70644
rect 472492 70604 475384 70632
rect 472492 70592 472498 70604
rect 475378 70592 475384 70604
rect 475436 70592 475442 70644
rect 83642 70456 83648 70508
rect 83700 70456 83706 70508
rect 83660 70372 83688 70456
rect 89898 70428 89904 70440
rect 89824 70400 89904 70428
rect 83642 70320 83648 70372
rect 83700 70320 83706 70372
rect 89824 70236 89852 70400
rect 89898 70388 89904 70400
rect 89956 70388 89962 70440
rect 280246 70388 280252 70440
rect 280304 70428 280310 70440
rect 280304 70400 280384 70428
rect 280304 70388 280310 70400
rect 280356 70372 280384 70400
rect 280338 70320 280344 70372
rect 280396 70320 280402 70372
rect 356701 70295 356759 70301
rect 356701 70261 356713 70295
rect 356747 70292 356759 70295
rect 356790 70292 356796 70304
rect 356747 70264 356796 70292
rect 356747 70261 356759 70264
rect 356701 70255 356759 70261
rect 356790 70252 356796 70264
rect 356848 70252 356854 70304
rect 89806 70184 89812 70236
rect 89864 70184 89870 70236
rect 338022 69708 338028 69760
rect 338080 69748 338086 69760
rect 496814 69748 496820 69760
rect 338080 69720 496820 69748
rect 338080 69708 338086 69720
rect 496814 69708 496820 69720
rect 496872 69708 496878 69760
rect 74074 69640 74080 69692
rect 74132 69680 74138 69692
rect 445754 69680 445760 69692
rect 74132 69652 445760 69680
rect 74132 69640 74138 69652
rect 445754 69640 445760 69652
rect 445812 69640 445818 69692
rect 469858 69232 469864 69284
rect 469916 69272 469922 69284
rect 472434 69272 472440 69284
rect 469916 69244 472440 69272
rect 469916 69232 469922 69244
rect 472434 69232 472440 69244
rect 472492 69232 472498 69284
rect 468938 69028 468944 69080
rect 468996 69068 469002 69080
rect 470502 69068 470508 69080
rect 468996 69040 470508 69068
rect 468996 69028 469002 69040
rect 470502 69028 470508 69040
rect 470560 69028 470566 69080
rect 128262 68416 128268 68468
rect 128320 68456 128326 68468
rect 289814 68456 289820 68468
rect 128320 68428 289820 68456
rect 128320 68416 128326 68428
rect 289814 68416 289820 68428
rect 289872 68416 289878 68468
rect 81710 68348 81716 68400
rect 81768 68388 81774 68400
rect 320174 68388 320180 68400
rect 81768 68360 320180 68388
rect 81768 68348 81774 68360
rect 320174 68348 320180 68360
rect 320232 68348 320238 68400
rect 348970 68348 348976 68400
rect 349028 68388 349034 68400
rect 502610 68388 502616 68400
rect 349028 68360 502616 68388
rect 349028 68348 349034 68360
rect 502610 68348 502616 68360
rect 502668 68348 502674 68400
rect 96522 68280 96528 68332
rect 96580 68320 96586 68332
rect 504174 68320 504180 68332
rect 96580 68292 504180 68320
rect 96580 68280 96586 68292
rect 504174 68280 504180 68292
rect 504232 68280 504238 68332
rect 79778 67600 79784 67652
rect 79836 67640 79842 67652
rect 79962 67640 79968 67652
rect 79836 67612 79968 67640
rect 79836 67600 79842 67612
rect 79962 67600 79968 67612
rect 80020 67600 80026 67652
rect 151449 67643 151507 67649
rect 151449 67609 151461 67643
rect 151495 67640 151507 67643
rect 151538 67640 151544 67652
rect 151495 67612 151544 67640
rect 151495 67609 151507 67612
rect 151449 67603 151507 67609
rect 151538 67600 151544 67612
rect 151596 67600 151602 67652
rect 176746 67640 176752 67652
rect 176707 67612 176752 67640
rect 176746 67600 176752 67612
rect 176804 67600 176810 67652
rect 198461 67643 198519 67649
rect 198461 67609 198473 67643
rect 198507 67640 198519 67643
rect 198550 67640 198556 67652
rect 198507 67612 198556 67640
rect 198507 67609 198519 67612
rect 198461 67603 198519 67609
rect 198550 67600 198556 67612
rect 198608 67600 198614 67652
rect 411162 67640 411168 67652
rect 411123 67612 411168 67640
rect 411162 67600 411168 67612
rect 411220 67600 411226 67652
rect 140774 67532 140780 67584
rect 140832 67572 140838 67584
rect 140866 67572 140872 67584
rect 140832 67544 140872 67572
rect 140832 67532 140838 67544
rect 140866 67532 140872 67544
rect 140924 67532 140930 67584
rect 467098 67464 467104 67516
rect 467156 67504 467162 67516
rect 469306 67504 469312 67516
rect 467156 67476 469312 67504
rect 467156 67464 467162 67476
rect 469306 67464 469312 67476
rect 469364 67464 469370 67516
rect 467190 67192 467196 67244
rect 467248 67232 467254 67244
rect 468938 67232 468944 67244
rect 467248 67204 468944 67232
rect 467248 67192 467254 67204
rect 468938 67192 468944 67204
rect 468996 67192 469002 67244
rect 256510 66920 256516 66972
rect 256568 66960 256574 66972
rect 303614 66960 303620 66972
rect 256568 66932 303620 66960
rect 256568 66920 256574 66932
rect 303614 66920 303620 66932
rect 303672 66920 303678 66972
rect 371142 66920 371148 66972
rect 371200 66960 371206 66972
rect 378226 66960 378232 66972
rect 371200 66932 378232 66960
rect 371200 66920 371206 66932
rect 378226 66920 378232 66932
rect 378284 66920 378290 66972
rect 119982 66852 119988 66904
rect 120040 66892 120046 66904
rect 508314 66892 508320 66904
rect 120040 66864 508320 66892
rect 120040 66852 120046 66864
rect 508314 66852 508320 66864
rect 508372 66852 508378 66904
rect 83366 66212 83372 66224
rect 83327 66184 83372 66212
rect 83366 66172 83372 66184
rect 83424 66172 83430 66224
rect 512822 66212 512828 66224
rect 512783 66184 512828 66212
rect 512822 66172 512828 66184
rect 512880 66172 512886 66224
rect 360102 65628 360108 65680
rect 360160 65668 360166 65680
rect 433334 65668 433340 65680
rect 360160 65640 433340 65668
rect 360160 65628 360166 65640
rect 433334 65628 433340 65640
rect 433392 65628 433398 65680
rect 315942 65560 315948 65612
rect 316000 65600 316006 65612
rect 505278 65600 505284 65612
rect 316000 65572 505284 65600
rect 316000 65560 316006 65572
rect 505278 65560 505284 65572
rect 505336 65560 505342 65612
rect 106182 65492 106188 65544
rect 106240 65532 106246 65544
rect 208394 65532 208400 65544
rect 106240 65504 208400 65532
rect 106240 65492 106246 65504
rect 208394 65492 208400 65504
rect 208452 65492 208458 65544
rect 210970 65492 210976 65544
rect 211028 65532 211034 65544
rect 504082 65532 504088 65544
rect 211028 65504 504088 65532
rect 211028 65492 211034 65504
rect 504082 65492 504088 65504
rect 504140 65492 504146 65544
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 33778 64852 33784 64864
rect 3384 64824 33784 64852
rect 3384 64812 3390 64824
rect 33778 64812 33784 64824
rect 33836 64812 33842 64864
rect 519538 64812 519544 64864
rect 519596 64852 519602 64864
rect 579798 64852 579804 64864
rect 519596 64824 579804 64852
rect 519596 64812 519602 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 88242 64132 88248 64184
rect 88300 64172 88306 64184
rect 509602 64172 509608 64184
rect 88300 64144 509608 64172
rect 88300 64132 88306 64144
rect 509602 64132 509608 64144
rect 509660 64132 509666 64184
rect 22002 62840 22008 62892
rect 22060 62880 22066 62892
rect 240778 62880 240784 62892
rect 22060 62852 240784 62880
rect 22060 62840 22066 62852
rect 240778 62840 240784 62852
rect 240836 62840 240842 62892
rect 165522 62772 165528 62824
rect 165580 62812 165586 62824
rect 506658 62812 506664 62824
rect 165580 62784 506664 62812
rect 165580 62772 165586 62784
rect 506658 62772 506664 62784
rect 506716 62772 506722 62824
rect 476758 62636 476764 62688
rect 476816 62676 476822 62688
rect 480898 62676 480904 62688
rect 476816 62648 480904 62676
rect 476816 62636 476822 62648
rect 480898 62636 480904 62648
rect 480956 62636 480962 62688
rect 465166 62092 465172 62144
rect 465224 62132 465230 62144
rect 467190 62132 467196 62144
rect 465224 62104 467196 62132
rect 465224 62092 465230 62104
rect 467190 62092 467196 62104
rect 467248 62092 467254 62144
rect 222102 61616 222108 61668
rect 222160 61656 222166 61668
rect 269114 61656 269120 61668
rect 222160 61628 269120 61656
rect 222160 61616 222166 61628
rect 269114 61616 269120 61628
rect 269172 61616 269178 61668
rect 75270 61548 75276 61600
rect 75328 61588 75334 61600
rect 267734 61588 267740 61600
rect 75328 61560 267740 61588
rect 75328 61548 75334 61560
rect 267734 61548 267740 61560
rect 267792 61548 267798 61600
rect 107470 61480 107476 61532
rect 107528 61520 107534 61532
rect 311986 61520 311992 61532
rect 107528 61492 311992 61520
rect 107528 61480 107534 61492
rect 311986 61480 311992 61492
rect 312044 61480 312050 61532
rect 260742 61412 260748 61464
rect 260800 61452 260806 61464
rect 502334 61452 502340 61464
rect 260800 61424 502340 61452
rect 260800 61412 260806 61424
rect 502334 61412 502340 61424
rect 502392 61412 502398 61464
rect 99282 61344 99288 61396
rect 99340 61384 99346 61396
rect 509510 61384 509516 61396
rect 99340 61356 509516 61384
rect 99340 61344 99346 61356
rect 509510 61344 509516 61356
rect 509568 61344 509574 61396
rect 151538 60840 151544 60852
rect 151464 60812 151544 60840
rect 89806 60732 89812 60784
rect 89864 60732 89870 60784
rect 79686 60664 79692 60716
rect 79744 60704 79750 60716
rect 79870 60704 79876 60716
rect 79744 60676 79876 60704
rect 79744 60664 79750 60676
rect 79870 60664 79876 60676
rect 79928 60664 79934 60716
rect 89824 60704 89852 60732
rect 151464 60716 151492 60812
rect 151538 60800 151544 60812
rect 151596 60800 151602 60852
rect 198550 60840 198556 60852
rect 198476 60812 198556 60840
rect 198476 60716 198504 60812
rect 198550 60800 198556 60812
rect 198608 60800 198614 60852
rect 482002 60732 482008 60784
rect 482060 60772 482066 60784
rect 483658 60772 483664 60784
rect 482060 60744 483664 60772
rect 482060 60732 482066 60744
rect 483658 60732 483664 60744
rect 483716 60732 483722 60784
rect 89990 60704 89996 60716
rect 89824 60676 89996 60704
rect 89990 60664 89996 60676
rect 90048 60664 90054 60716
rect 151446 60664 151452 60716
rect 151504 60664 151510 60716
rect 198458 60664 198464 60716
rect 198516 60664 198522 60716
rect 333882 60120 333888 60172
rect 333940 60160 333946 60172
rect 456794 60160 456800 60172
rect 333940 60132 456800 60160
rect 333940 60120 333946 60132
rect 456794 60120 456800 60132
rect 456852 60120 456858 60172
rect 45462 60052 45468 60104
rect 45520 60092 45526 60104
rect 370590 60092 370596 60104
rect 45520 60064 370596 60092
rect 45520 60052 45526 60064
rect 370590 60052 370596 60064
rect 370648 60052 370654 60104
rect 467742 60052 467748 60104
rect 467800 60092 467806 60104
rect 494054 60092 494060 60104
rect 467800 60064 494060 60092
rect 467800 60052 467806 60064
rect 494054 60052 494060 60064
rect 494112 60052 494118 60104
rect 97902 59984 97908 60036
rect 97960 60024 97966 60036
rect 504358 60024 504364 60036
rect 97960 59996 504364 60024
rect 97960 59984 97966 59996
rect 504358 59984 504364 59996
rect 504416 59984 504422 60036
rect 144638 58760 144644 58812
rect 144696 58800 144702 58812
rect 396166 58800 396172 58812
rect 144696 58772 396172 58800
rect 144696 58760 144702 58772
rect 396166 58760 396172 58772
rect 396224 58760 396230 58812
rect 68830 58692 68836 58744
rect 68888 58732 68894 58744
rect 323578 58732 323584 58744
rect 68888 58704 323584 58732
rect 68888 58692 68894 58704
rect 323578 58692 323584 58704
rect 323636 58692 323642 58744
rect 219250 58624 219256 58676
rect 219308 58664 219314 58676
rect 506566 58664 506572 58676
rect 219308 58636 506572 58664
rect 219308 58624 219314 58636
rect 506566 58624 506572 58636
rect 506624 58624 506630 58676
rect 445570 57944 445576 57996
rect 445628 57984 445634 57996
rect 445662 57984 445668 57996
rect 445628 57956 445668 57984
rect 445628 57944 445634 57956
rect 445662 57944 445668 57956
rect 445720 57944 445726 57996
rect 79870 57916 79876 57928
rect 79831 57888 79876 57916
rect 79870 57876 79876 57888
rect 79928 57876 79934 57928
rect 89901 57919 89959 57925
rect 89901 57885 89913 57919
rect 89947 57916 89959 57919
rect 89990 57916 89996 57928
rect 89947 57888 89996 57916
rect 89947 57885 89959 57888
rect 89901 57879 89959 57885
rect 89990 57876 89996 57888
rect 90048 57876 90054 57928
rect 140682 57876 140688 57928
rect 140740 57916 140746 57928
rect 140774 57916 140780 57928
rect 140740 57888 140780 57916
rect 140740 57876 140746 57888
rect 140774 57876 140780 57888
rect 140832 57876 140838 57928
rect 144730 57916 144736 57928
rect 144691 57888 144736 57916
rect 144730 57876 144736 57888
rect 144788 57876 144794 57928
rect 176749 57919 176807 57925
rect 176749 57885 176761 57919
rect 176795 57916 176807 57919
rect 176838 57916 176844 57928
rect 176795 57888 176844 57916
rect 176795 57885 176807 57888
rect 176749 57879 176807 57885
rect 176838 57876 176844 57888
rect 176896 57876 176902 57928
rect 198458 57916 198464 57928
rect 198419 57888 198464 57916
rect 198458 57876 198464 57888
rect 198516 57876 198522 57928
rect 212442 57916 212448 57928
rect 212403 57888 212448 57916
rect 212442 57876 212448 57888
rect 212500 57876 212506 57928
rect 280341 57919 280399 57925
rect 280341 57885 280353 57919
rect 280387 57916 280399 57919
rect 280430 57916 280436 57928
rect 280387 57888 280436 57916
rect 280387 57885 280399 57888
rect 280341 57879 280399 57885
rect 280430 57876 280436 57888
rect 280488 57876 280494 57928
rect 333882 57916 333888 57928
rect 333843 57888 333888 57916
rect 333882 57876 333888 57888
rect 333940 57876 333946 57928
rect 356606 57916 356612 57928
rect 356567 57888 356612 57916
rect 356606 57876 356612 57888
rect 356664 57876 356670 57928
rect 411162 57916 411168 57928
rect 411123 57888 411168 57916
rect 411162 57876 411168 57888
rect 411220 57876 411226 57928
rect 83369 57851 83427 57857
rect 83369 57817 83381 57851
rect 83415 57848 83427 57851
rect 83550 57848 83556 57860
rect 83415 57820 83556 57848
rect 83415 57817 83427 57820
rect 83369 57811 83427 57817
rect 83550 57808 83556 57820
rect 83608 57808 83614 57860
rect 462406 57808 462412 57860
rect 462464 57848 462470 57860
rect 465166 57848 465172 57860
rect 462464 57820 465172 57848
rect 462464 57808 462470 57820
rect 465166 57808 465172 57820
rect 465224 57808 465230 57860
rect 467834 57740 467840 57792
rect 467892 57780 467898 57792
rect 469858 57780 469864 57792
rect 467892 57752 469864 57780
rect 467892 57740 467898 57752
rect 469858 57740 469864 57752
rect 469916 57740 469922 57792
rect 344830 57264 344836 57316
rect 344888 57304 344894 57316
rect 527174 57304 527180 57316
rect 344888 57276 527180 57304
rect 344888 57264 344894 57276
rect 527174 57264 527180 57276
rect 527232 57264 527238 57316
rect 83642 57196 83648 57248
rect 83700 57236 83706 57248
rect 376754 57236 376760 57248
rect 83700 57208 376760 57236
rect 83700 57196 83706 57208
rect 376754 57196 376760 57208
rect 376812 57196 376818 57248
rect 380802 57196 380808 57248
rect 380860 57236 380866 57248
rect 431954 57236 431960 57248
rect 380860 57208 431960 57236
rect 380860 57196 380866 57208
rect 431954 57196 431960 57208
rect 432012 57196 432018 57248
rect 512822 56624 512828 56636
rect 512783 56596 512828 56624
rect 512822 56584 512828 56596
rect 512880 56584 512886 56636
rect 140682 56556 140688 56568
rect 140643 56528 140688 56556
rect 140682 56516 140688 56528
rect 140740 56516 140746 56568
rect 81526 55972 81532 56024
rect 81584 56012 81590 56024
rect 350626 56012 350632 56024
rect 81584 55984 350632 56012
rect 81584 55972 81590 55984
rect 350626 55972 350632 55984
rect 350684 55972 350690 56024
rect 354490 55972 354496 56024
rect 354548 56012 354554 56024
rect 419534 56012 419540 56024
rect 354548 55984 419540 56012
rect 354548 55972 354554 55984
rect 419534 55972 419540 55984
rect 419592 55972 419598 56024
rect 478874 55972 478880 56024
rect 478932 56012 478938 56024
rect 482002 56012 482008 56024
rect 478932 55984 482008 56012
rect 478932 55972 478938 55984
rect 482002 55972 482008 55984
rect 482060 55972 482066 56024
rect 220630 55904 220636 55956
rect 220688 55944 220694 55956
rect 505094 55944 505100 55956
rect 220688 55916 505100 55944
rect 220688 55904 220694 55916
rect 505094 55904 505100 55916
rect 505152 55904 505158 55956
rect 15102 55836 15108 55888
rect 15160 55876 15166 55888
rect 131758 55876 131764 55888
rect 15160 55848 131764 55876
rect 15160 55836 15166 55848
rect 131758 55836 131764 55848
rect 131816 55836 131822 55888
rect 136542 55836 136548 55888
rect 136600 55876 136606 55888
rect 503806 55876 503812 55888
rect 136600 55848 503812 55876
rect 136600 55836 136606 55848
rect 503806 55836 503812 55848
rect 503864 55836 503870 55888
rect 472894 53864 472900 53916
rect 472952 53904 472958 53916
rect 478874 53904 478880 53916
rect 472952 53876 478880 53904
rect 472952 53864 472958 53876
rect 478874 53864 478880 53876
rect 478932 53864 478938 53916
rect 464338 53796 464344 53848
rect 464396 53836 464402 53848
rect 467834 53836 467840 53848
rect 464396 53808 467840 53836
rect 464396 53796 464402 53808
rect 467834 53796 467840 53808
rect 467892 53796 467898 53848
rect 391750 53048 391756 53100
rect 391808 53088 391814 53100
rect 487154 53088 487160 53100
rect 391808 53060 487160 53088
rect 391808 53048 391814 53060
rect 487154 53048 487160 53060
rect 487212 53048 487218 53100
rect 467834 52436 467840 52488
rect 467892 52476 467898 52488
rect 472894 52476 472900 52488
rect 467892 52448 472900 52476
rect 467892 52436 467898 52448
rect 472894 52436 472900 52448
rect 472952 52436 472958 52488
rect 473998 52436 474004 52488
rect 474056 52476 474062 52488
rect 476758 52476 476764 52488
rect 474056 52448 476764 52476
rect 474056 52436 474062 52448
rect 476758 52436 476764 52448
rect 476816 52436 476822 52488
rect 80882 51688 80888 51740
rect 80940 51728 80946 51740
rect 382274 51728 382280 51740
rect 80940 51700 382280 51728
rect 80940 51688 80946 51700
rect 382274 51688 382280 51700
rect 382332 51688 382338 51740
rect 384942 51688 384948 51740
rect 385000 51728 385006 51740
rect 476114 51728 476120 51740
rect 385000 51700 476120 51728
rect 385000 51688 385006 51700
rect 476114 51688 476120 51700
rect 476172 51688 476178 51740
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 71038 51048 71044 51060
rect 3476 51020 71044 51048
rect 3476 51008 3482 51020
rect 71038 51008 71044 51020
rect 71096 51008 71102 51060
rect 151446 51008 151452 51060
rect 151504 51048 151510 51060
rect 151630 51048 151636 51060
rect 151504 51020 151636 51048
rect 151504 51008 151510 51020
rect 151630 51008 151636 51020
rect 151688 51008 151694 51060
rect 79870 50912 79876 50924
rect 79831 50884 79876 50912
rect 79870 50872 79876 50884
rect 79928 50872 79934 50924
rect 357250 50396 357256 50448
rect 357308 50436 357314 50448
rect 415394 50436 415400 50448
rect 357308 50408 415400 50436
rect 357308 50396 357314 50408
rect 415394 50396 415400 50408
rect 415452 50396 415458 50448
rect 78490 50328 78496 50380
rect 78548 50368 78554 50380
rect 234614 50368 234620 50380
rect 78548 50340 234620 50368
rect 78548 50328 78554 50340
rect 234614 50328 234620 50340
rect 234672 50328 234678 50380
rect 250990 50328 250996 50380
rect 251048 50368 251054 50380
rect 393314 50368 393320 50380
rect 251048 50340 393320 50368
rect 251048 50328 251054 50340
rect 393314 50328 393320 50340
rect 393372 50328 393378 50380
rect 461578 49648 461584 49700
rect 461636 49688 461642 49700
rect 462406 49688 462412 49700
rect 461636 49660 462412 49688
rect 461636 49648 461642 49660
rect 462406 49648 462412 49660
rect 462464 49648 462470 49700
rect 382182 49104 382188 49156
rect 382240 49144 382246 49156
rect 540974 49144 540980 49156
rect 382240 49116 540980 49144
rect 382240 49104 382246 49116
rect 540974 49104 540980 49116
rect 541032 49104 541038 49156
rect 81618 49036 81624 49088
rect 81676 49076 81682 49088
rect 404354 49076 404360 49088
rect 81676 49048 404360 49076
rect 81676 49036 81682 49048
rect 404354 49036 404360 49048
rect 404412 49036 404418 49088
rect 153102 48968 153108 49020
rect 153160 49008 153166 49020
rect 507026 49008 507032 49020
rect 153160 48980 507032 49008
rect 153160 48968 153166 48980
rect 507026 48968 507032 48980
rect 507084 48968 507090 49020
rect 89898 48328 89904 48340
rect 89859 48300 89904 48328
rect 89898 48288 89904 48300
rect 89956 48288 89962 48340
rect 144730 48328 144736 48340
rect 144691 48300 144736 48328
rect 144730 48288 144736 48300
rect 144788 48288 144794 48340
rect 176746 48328 176752 48340
rect 176707 48300 176752 48328
rect 176746 48288 176752 48300
rect 176804 48288 176810 48340
rect 198461 48331 198519 48337
rect 198461 48297 198473 48331
rect 198507 48328 198519 48331
rect 198550 48328 198556 48340
rect 198507 48300 198556 48328
rect 198507 48297 198519 48300
rect 198461 48291 198519 48297
rect 198550 48288 198556 48300
rect 198608 48288 198614 48340
rect 210970 48328 210976 48340
rect 210931 48300 210976 48328
rect 210970 48288 210976 48300
rect 211028 48288 211034 48340
rect 212442 48328 212448 48340
rect 212403 48300 212448 48328
rect 212442 48288 212448 48300
rect 212500 48288 212506 48340
rect 280338 48328 280344 48340
rect 280299 48300 280344 48328
rect 280338 48288 280344 48300
rect 280396 48288 280402 48340
rect 333882 48328 333888 48340
rect 333843 48300 333888 48328
rect 333882 48288 333888 48300
rect 333940 48288 333946 48340
rect 356609 48331 356667 48337
rect 356609 48297 356621 48331
rect 356655 48328 356667 48331
rect 356698 48328 356704 48340
rect 356655 48300 356704 48328
rect 356655 48297 356667 48300
rect 356609 48291 356667 48297
rect 356698 48288 356704 48300
rect 356756 48288 356762 48340
rect 411162 48328 411168 48340
rect 411123 48300 411168 48328
rect 411162 48288 411168 48300
rect 411220 48288 411226 48340
rect 151541 48263 151599 48269
rect 151541 48229 151553 48263
rect 151587 48260 151599 48263
rect 151630 48260 151636 48272
rect 151587 48232 151636 48260
rect 151587 48229 151599 48232
rect 151541 48223 151599 48229
rect 151630 48220 151636 48232
rect 151688 48220 151694 48272
rect 465810 47880 465816 47932
rect 465868 47920 465874 47932
rect 467834 47920 467840 47932
rect 465868 47892 467840 47920
rect 465868 47880 465874 47892
rect 467834 47880 467840 47892
rect 467892 47880 467898 47932
rect 90910 47540 90916 47592
rect 90968 47580 90974 47592
rect 200114 47580 200120 47592
rect 90968 47552 200120 47580
rect 90968 47540 90974 47552
rect 200114 47540 200120 47552
rect 200172 47540 200178 47592
rect 140685 46971 140743 46977
rect 140685 46937 140697 46971
rect 140731 46968 140743 46971
rect 140774 46968 140780 46980
rect 140731 46940 140780 46968
rect 140731 46937 140743 46940
rect 140685 46931 140743 46937
rect 140774 46928 140780 46940
rect 140832 46928 140838 46980
rect 210970 46968 210976 46980
rect 210931 46940 210976 46968
rect 210970 46928 210976 46940
rect 211028 46928 211034 46980
rect 512822 46900 512828 46912
rect 512783 46872 512828 46900
rect 512822 46860 512828 46872
rect 512880 46860 512886 46912
rect 83366 46248 83372 46300
rect 83424 46288 83430 46300
rect 237466 46288 237472 46300
rect 83424 46260 237472 46288
rect 83424 46248 83430 46260
rect 237466 46248 237472 46260
rect 237524 46248 237530 46300
rect 281442 46248 281448 46300
rect 281500 46288 281506 46300
rect 333974 46288 333980 46300
rect 281500 46260 333980 46288
rect 281500 46248 281506 46260
rect 333974 46248 333980 46260
rect 334032 46248 334038 46300
rect 335262 46248 335268 46300
rect 335320 46288 335326 46300
rect 429194 46288 429200 46300
rect 335320 46260 429200 46288
rect 335320 46248 335326 46260
rect 429194 46248 429200 46260
rect 429252 46248 429258 46300
rect 155862 46180 155868 46232
rect 155920 46220 155926 46232
rect 492674 46220 492680 46232
rect 155920 46192 492680 46220
rect 155920 46180 155926 46192
rect 492674 46180 492680 46192
rect 492732 46180 492738 46232
rect 140774 45540 140780 45552
rect 140735 45512 140780 45540
rect 140774 45500 140780 45512
rect 140832 45500 140838 45552
rect 103422 44888 103428 44940
rect 103480 44928 103486 44940
rect 425054 44928 425060 44940
rect 103480 44900 425060 44928
rect 103480 44888 103486 44900
rect 425054 44888 425060 44900
rect 425112 44888 425118 44940
rect 223482 44820 223488 44872
rect 223540 44860 223546 44872
rect 565814 44860 565820 44872
rect 223540 44832 565820 44860
rect 223540 44820 223546 44832
rect 565814 44820 565820 44832
rect 565872 44820 565878 44872
rect 461578 44180 461584 44192
rect 459572 44152 461584 44180
rect 456058 44004 456064 44056
rect 456116 44044 456122 44056
rect 459572 44044 459600 44152
rect 461578 44140 461584 44152
rect 461636 44140 461642 44192
rect 456116 44016 459600 44044
rect 456116 44004 456122 44016
rect 462682 43528 462688 43580
rect 462740 43568 462746 43580
rect 464338 43568 464344 43580
rect 462740 43540 464344 43568
rect 462740 43528 462746 43540
rect 464338 43528 464344 43540
rect 464396 43528 464402 43580
rect 110230 43460 110236 43512
rect 110288 43500 110294 43512
rect 506934 43500 506940 43512
rect 110288 43472 506940 43500
rect 110288 43460 110294 43472
rect 506934 43460 506940 43472
rect 506992 43460 506998 43512
rect 78030 43392 78036 43444
rect 78088 43432 78094 43444
rect 538214 43432 538220 43444
rect 78088 43404 538220 43432
rect 78088 43392 78094 43404
rect 538214 43392 538220 43404
rect 538272 43392 538278 43444
rect 463786 42780 463792 42832
rect 463844 42820 463850 42832
rect 465810 42820 465816 42832
rect 463844 42792 465816 42820
rect 463844 42780 463850 42792
rect 465810 42780 465816 42792
rect 465868 42780 465874 42832
rect 235902 42100 235908 42152
rect 235960 42140 235966 42152
rect 492674 42140 492680 42152
rect 235960 42112 492680 42140
rect 235960 42100 235966 42112
rect 492674 42100 492680 42112
rect 492732 42100 492738 42152
rect 79502 42032 79508 42084
rect 79560 42072 79566 42084
rect 358814 42072 358820 42084
rect 79560 42044 358820 42072
rect 79560 42032 79566 42044
rect 358814 42032 358820 42044
rect 358872 42032 358878 42084
rect 469306 42032 469312 42084
rect 469364 42072 469370 42084
rect 473998 42072 474004 42084
rect 469364 42044 474004 42072
rect 469364 42032 469370 42044
rect 473998 42032 474004 42044
rect 474056 42032 474062 42084
rect 198550 41460 198556 41472
rect 198476 41432 198556 41460
rect 198476 41404 198504 41432
rect 198550 41420 198556 41432
rect 198608 41420 198614 41472
rect 460198 41420 460204 41472
rect 460256 41460 460262 41472
rect 462682 41460 462688 41472
rect 460256 41432 462688 41460
rect 460256 41420 460262 41432
rect 462682 41420 462688 41432
rect 462740 41420 462746 41472
rect 89806 41352 89812 41404
rect 89864 41392 89870 41404
rect 89990 41392 89996 41404
rect 89864 41364 89996 41392
rect 89864 41352 89870 41364
rect 89990 41352 89996 41364
rect 90048 41352 90054 41404
rect 198458 41352 198464 41404
rect 198516 41352 198522 41404
rect 549898 41352 549904 41404
rect 549956 41392 549962 41404
rect 580166 41392 580172 41404
rect 549956 41364 580172 41392
rect 549956 41352 549962 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 76742 40740 76748 40792
rect 76800 40780 76806 40792
rect 367094 40780 367100 40792
rect 76800 40752 367100 40780
rect 76800 40740 76806 40752
rect 367094 40740 367100 40752
rect 367152 40740 367158 40792
rect 391842 40740 391848 40792
rect 391900 40780 391906 40792
rect 441614 40780 441620 40792
rect 391900 40752 441620 40780
rect 391900 40740 391906 40752
rect 441614 40740 441620 40752
rect 441672 40740 441678 40792
rect 104802 40672 104808 40724
rect 104860 40712 104866 40724
rect 494054 40712 494060 40724
rect 104860 40684 494060 40712
rect 104860 40672 104866 40684
rect 494054 40672 494060 40684
rect 494112 40672 494118 40724
rect 465718 40060 465724 40112
rect 465776 40100 465782 40112
rect 469306 40100 469312 40112
rect 465776 40072 469312 40100
rect 465776 40060 465782 40072
rect 469306 40060 469312 40072
rect 469364 40060 469370 40112
rect 461578 39856 461584 39908
rect 461636 39896 461642 39908
rect 463786 39896 463792 39908
rect 461636 39868 463792 39896
rect 461636 39856 461642 39868
rect 463786 39856 463792 39868
rect 463844 39856 463850 39908
rect 360838 39380 360844 39432
rect 360896 39420 360902 39432
rect 370498 39420 370504 39432
rect 360896 39392 370504 39420
rect 360896 39380 360902 39392
rect 370498 39380 370504 39392
rect 370556 39380 370562 39432
rect 307570 39312 307576 39364
rect 307628 39352 307634 39364
rect 520458 39352 520464 39364
rect 307628 39324 520464 39352
rect 307628 39312 307634 39324
rect 520458 39312 520464 39324
rect 520516 39312 520522 39364
rect 151538 38672 151544 38684
rect 151499 38644 151544 38672
rect 151538 38632 151544 38644
rect 151596 38632 151602 38684
rect 445570 38632 445576 38684
rect 445628 38672 445634 38684
rect 445662 38672 445668 38684
rect 445628 38644 445668 38672
rect 445628 38632 445634 38644
rect 445662 38632 445668 38644
rect 445720 38632 445726 38684
rect 144730 38604 144736 38616
rect 144691 38576 144736 38604
rect 144730 38564 144736 38576
rect 144788 38564 144794 38616
rect 176749 38607 176807 38613
rect 176749 38573 176761 38607
rect 176795 38604 176807 38607
rect 176838 38604 176844 38616
rect 176795 38576 176844 38604
rect 176795 38573 176807 38576
rect 176749 38567 176807 38573
rect 176838 38564 176844 38576
rect 176896 38564 176902 38616
rect 198458 38604 198464 38616
rect 198419 38576 198464 38604
rect 198458 38564 198464 38576
rect 198516 38564 198522 38616
rect 280341 38607 280399 38613
rect 280341 38573 280353 38607
rect 280387 38604 280399 38607
rect 280430 38604 280436 38616
rect 280387 38576 280436 38604
rect 280387 38573 280399 38576
rect 280341 38567 280399 38573
rect 280430 38564 280436 38576
rect 280488 38564 280494 38616
rect 161382 38020 161388 38072
rect 161440 38060 161446 38072
rect 356882 38060 356888 38072
rect 161440 38032 356888 38060
rect 161440 38020 161446 38032
rect 356882 38020 356888 38032
rect 356940 38020 356946 38072
rect 228818 37952 228824 38004
rect 228876 37992 228882 38004
rect 501506 37992 501512 38004
rect 228876 37964 501512 37992
rect 228876 37952 228882 37964
rect 501506 37952 501512 37964
rect 501564 37952 501570 38004
rect 79870 37884 79876 37936
rect 79928 37924 79934 37936
rect 436094 37924 436100 37936
rect 79928 37896 436100 37924
rect 79928 37884 79934 37896
rect 436094 37884 436100 37896
rect 436152 37884 436158 37936
rect 210970 37272 210976 37324
rect 211028 37312 211034 37324
rect 211062 37312 211068 37324
rect 211028 37284 211068 37312
rect 211028 37272 211034 37284
rect 211062 37272 211068 37284
rect 211120 37272 211126 37324
rect 512822 37312 512828 37324
rect 512783 37284 512828 37312
rect 512822 37272 512828 37284
rect 512880 37272 512886 37324
rect 140777 35955 140835 35961
rect 140777 35921 140789 35955
rect 140823 35952 140835 35955
rect 140866 35952 140872 35964
rect 140823 35924 140872 35952
rect 140823 35921 140835 35924
rect 140777 35915 140835 35921
rect 140866 35912 140872 35924
rect 140924 35912 140930 35964
rect 458266 34484 458272 34536
rect 458324 34524 458330 34536
rect 461578 34524 461584 34536
rect 458324 34496 461584 34524
rect 458324 34484 458330 34496
rect 461578 34484 461584 34496
rect 461636 34484 461642 34536
rect 462958 34484 462964 34536
rect 463016 34524 463022 34536
rect 465718 34524 465724 34536
rect 463016 34496 465724 34524
rect 463016 34484 463022 34496
rect 465718 34484 465724 34496
rect 465776 34484 465782 34536
rect 451182 33804 451188 33856
rect 451240 33844 451246 33856
rect 574738 33844 574744 33856
rect 451240 33816 574744 33844
rect 451240 33804 451246 33816
rect 574738 33804 574744 33816
rect 574796 33804 574802 33856
rect 248230 33736 248236 33788
rect 248288 33776 248294 33788
rect 495434 33776 495440 33788
rect 248288 33748 495440 33776
rect 248288 33736 248294 33748
rect 495434 33736 495440 33748
rect 495492 33736 495498 33788
rect 182082 32512 182088 32564
rect 182140 32552 182146 32564
rect 252554 32552 252560 32564
rect 182140 32524 252560 32552
rect 182140 32512 182146 32524
rect 252554 32512 252560 32524
rect 252612 32512 252618 32564
rect 219342 32444 219348 32496
rect 219400 32484 219406 32496
rect 294046 32484 294052 32496
rect 219400 32456 294052 32484
rect 219400 32444 219406 32456
rect 294046 32444 294052 32456
rect 294104 32444 294110 32496
rect 353294 32444 353300 32496
rect 353352 32484 353358 32496
rect 360838 32484 360844 32496
rect 353352 32456 360844 32484
rect 353352 32444 353358 32456
rect 360838 32444 360844 32456
rect 360896 32444 360902 32496
rect 78582 32376 78588 32428
rect 78640 32416 78646 32428
rect 223574 32416 223580 32428
rect 78640 32388 223580 32416
rect 78640 32376 78646 32388
rect 223574 32376 223580 32388
rect 223632 32376 223638 32428
rect 256602 32376 256608 32428
rect 256660 32416 256666 32428
rect 460934 32416 460940 32428
rect 256660 32388 460940 32416
rect 256660 32376 256666 32388
rect 460934 32376 460940 32388
rect 460992 32376 460998 32428
rect 89990 31804 89996 31816
rect 89951 31776 89996 31804
rect 89990 31764 89996 31776
rect 90048 31764 90054 31816
rect 176746 31736 176752 31748
rect 176707 31708 176752 31736
rect 176746 31696 176752 31708
rect 176804 31696 176810 31748
rect 280338 31736 280344 31748
rect 280299 31708 280344 31736
rect 280338 31696 280344 31708
rect 280396 31696 280402 31748
rect 198461 31671 198519 31677
rect 198461 31637 198473 31671
rect 198507 31668 198519 31671
rect 198550 31668 198556 31680
rect 198507 31640 198556 31668
rect 198507 31637 198519 31640
rect 198461 31631 198519 31637
rect 198550 31628 198556 31640
rect 198608 31628 198614 31680
rect 237190 31016 237196 31068
rect 237248 31056 237254 31068
rect 311894 31056 311900 31068
rect 237248 31028 311900 31056
rect 237248 31016 237254 31028
rect 311894 31016 311900 31028
rect 311952 31016 311958 31068
rect 409782 31016 409788 31068
rect 409840 31056 409846 31068
rect 469214 31056 469220 31068
rect 409840 31028 469220 31056
rect 409840 31016 409846 31028
rect 469214 31016 469220 31028
rect 469272 31016 469278 31068
rect 457438 30200 457444 30252
rect 457496 30240 457502 30252
rect 458266 30240 458272 30252
rect 457496 30212 458272 30240
rect 457496 30200 457502 30212
rect 458266 30200 458272 30212
rect 458324 30200 458330 30252
rect 9582 29724 9588 29776
rect 9640 29764 9646 29776
rect 207658 29764 207664 29776
rect 9640 29736 207664 29764
rect 9640 29724 9646 29736
rect 207658 29724 207664 29736
rect 207716 29724 207722 29776
rect 297818 29724 297824 29776
rect 297876 29764 297882 29776
rect 430574 29764 430580 29776
rect 297876 29736 430580 29764
rect 297876 29724 297882 29736
rect 430574 29724 430580 29736
rect 430632 29724 430638 29776
rect 184842 29656 184848 29708
rect 184900 29696 184906 29708
rect 484394 29696 484400 29708
rect 184900 29668 484400 29696
rect 184900 29656 184906 29668
rect 484394 29656 484400 29668
rect 484452 29656 484458 29708
rect 204070 29588 204076 29640
rect 204128 29628 204134 29640
rect 506842 29628 506848 29640
rect 204128 29600 506848 29628
rect 204128 29588 204134 29600
rect 506842 29588 506848 29600
rect 506900 29588 506906 29640
rect 553118 29180 553124 29232
rect 553176 29220 553182 29232
rect 560202 29220 560208 29232
rect 553176 29192 560208 29220
rect 553176 29180 553182 29192
rect 560202 29180 560208 29192
rect 560260 29180 560266 29232
rect 89898 29044 89904 29096
rect 89956 29084 89962 29096
rect 89993 29087 90051 29093
rect 89993 29084 90005 29087
rect 89956 29056 90005 29084
rect 89956 29044 89962 29056
rect 89993 29053 90005 29056
rect 90039 29053 90051 29087
rect 89993 29047 90051 29053
rect 144730 29016 144736 29028
rect 144691 28988 144736 29016
rect 144730 28976 144736 28988
rect 144788 28976 144794 29028
rect 411162 28908 411168 28960
rect 411220 28948 411226 28960
rect 411346 28948 411352 28960
rect 411220 28920 411352 28948
rect 411220 28908 411226 28920
rect 411346 28908 411352 28920
rect 411404 28908 411410 28960
rect 103422 28364 103428 28416
rect 103480 28404 103486 28416
rect 420914 28404 420920 28416
rect 103480 28376 420920 28404
rect 103480 28364 103486 28376
rect 420914 28364 420920 28376
rect 420972 28364 420978 28416
rect 423582 28364 423588 28416
rect 423640 28404 423646 28416
rect 440234 28404 440240 28416
rect 423640 28376 440240 28404
rect 423640 28364 423646 28376
rect 440234 28364 440240 28376
rect 440292 28364 440298 28416
rect 137922 28296 137928 28348
rect 137980 28336 137986 28348
rect 491294 28336 491300 28348
rect 137980 28308 491300 28336
rect 137980 28296 137986 28308
rect 491294 28296 491300 28308
rect 491352 28296 491358 28348
rect 144822 28228 144828 28280
rect 144880 28268 144886 28280
rect 581086 28268 581092 28280
rect 144880 28240 581092 28268
rect 144880 28228 144886 28240
rect 581086 28228 581092 28240
rect 581144 28228 581150 28280
rect 89806 27588 89812 27600
rect 89767 27560 89812 27588
rect 89806 27548 89812 27560
rect 89864 27548 89870 27600
rect 210970 27588 210976 27600
rect 210931 27560 210976 27588
rect 210970 27548 210976 27560
rect 211028 27548 211034 27600
rect 512457 27591 512515 27597
rect 512457 27557 512469 27591
rect 512503 27588 512515 27591
rect 512822 27588 512828 27600
rect 512503 27560 512828 27588
rect 512503 27557 512515 27560
rect 512457 27551 512515 27557
rect 512822 27548 512828 27560
rect 512880 27548 512886 27600
rect 351178 27208 351184 27260
rect 351236 27248 351242 27260
rect 353294 27248 353300 27260
rect 351236 27220 353300 27248
rect 351236 27208 351242 27220
rect 353294 27208 353300 27220
rect 353352 27208 353358 27260
rect 38562 26936 38568 26988
rect 38620 26976 38626 26988
rect 153194 26976 153200 26988
rect 38620 26948 153200 26976
rect 38620 26936 38626 26948
rect 153194 26936 153200 26948
rect 153252 26936 153258 26988
rect 266262 26936 266268 26988
rect 266320 26976 266326 26988
rect 401594 26976 401600 26988
rect 266320 26948 401600 26976
rect 266320 26936 266326 26948
rect 401594 26936 401600 26948
rect 401652 26936 401658 26988
rect 151446 26868 151452 26920
rect 151504 26908 151510 26920
rect 539594 26908 539600 26920
rect 151504 26880 539600 26908
rect 151504 26868 151510 26880
rect 539594 26868 539600 26880
rect 539652 26868 539658 26920
rect 97902 25712 97908 25764
rect 97960 25752 97966 25764
rect 251818 25752 251824 25764
rect 97960 25724 251824 25752
rect 97960 25712 97966 25724
rect 251818 25712 251824 25724
rect 251876 25712 251882 25764
rect 246942 25644 246948 25696
rect 247000 25684 247006 25696
rect 462314 25684 462320 25696
rect 247000 25656 462320 25684
rect 247000 25644 247006 25656
rect 462314 25644 462320 25656
rect 462372 25644 462378 25696
rect 100662 25576 100668 25628
rect 100720 25616 100726 25628
rect 408494 25616 408500 25628
rect 100720 25588 408500 25616
rect 100720 25576 100726 25588
rect 408494 25576 408500 25588
rect 408552 25576 408558 25628
rect 20622 25508 20628 25560
rect 20680 25548 20686 25560
rect 91094 25548 91100 25560
rect 20680 25520 91100 25548
rect 20680 25508 20686 25520
rect 91094 25508 91100 25520
rect 91152 25508 91158 25560
rect 110322 25508 110328 25560
rect 110380 25548 110386 25560
rect 550634 25548 550640 25560
rect 110380 25520 550640 25548
rect 110380 25508 110386 25520
rect 550634 25508 550640 25520
rect 550692 25508 550698 25560
rect 216490 24148 216496 24200
rect 216548 24188 216554 24200
rect 233326 24188 233332 24200
rect 216548 24160 233332 24188
rect 216548 24148 216554 24160
rect 233326 24148 233332 24160
rect 233384 24148 233390 24200
rect 75730 24080 75736 24132
rect 75788 24120 75794 24132
rect 281534 24120 281540 24132
rect 75788 24092 281540 24120
rect 75788 24080 75794 24092
rect 281534 24080 281540 24092
rect 281592 24080 281598 24132
rect 465718 23468 465724 23520
rect 465776 23508 465782 23520
rect 467098 23508 467104 23520
rect 465776 23480 467104 23508
rect 465776 23468 465782 23480
rect 467098 23468 467104 23480
rect 467156 23468 467162 23520
rect 26142 23128 26148 23180
rect 26200 23168 26206 23180
rect 28258 23168 28264 23180
rect 26200 23140 28264 23168
rect 26200 23128 26206 23140
rect 28258 23128 28264 23140
rect 28316 23128 28322 23180
rect 28902 22788 28908 22840
rect 28960 22828 28966 22840
rect 142798 22828 142804 22840
rect 28960 22800 142804 22828
rect 28960 22788 28966 22800
rect 142798 22788 142804 22800
rect 142856 22788 142862 22840
rect 269022 22788 269028 22840
rect 269080 22828 269086 22840
rect 400214 22828 400220 22840
rect 269080 22800 400220 22828
rect 269080 22788 269086 22800
rect 400214 22788 400220 22800
rect 400272 22788 400278 22840
rect 81802 22720 81808 22772
rect 81860 22760 81866 22772
rect 552014 22760 552020 22772
rect 81860 22732 552020 22760
rect 81860 22720 81866 22732
rect 552014 22720 552020 22732
rect 552072 22720 552078 22772
rect 140777 22695 140835 22701
rect 140777 22661 140789 22695
rect 140823 22692 140835 22695
rect 140866 22692 140872 22704
rect 140823 22664 140872 22692
rect 140823 22661 140835 22664
rect 140777 22655 140835 22661
rect 140866 22652 140872 22664
rect 140924 22652 140930 22704
rect 452562 22176 452568 22228
rect 452620 22216 452626 22228
rect 456058 22216 456064 22228
rect 452620 22188 456064 22216
rect 452620 22176 452626 22188
rect 456058 22176 456064 22188
rect 456116 22176 456122 22228
rect 455414 22108 455420 22160
rect 455472 22148 455478 22160
rect 457438 22148 457444 22160
rect 455472 22120 457444 22148
rect 455472 22108 455478 22120
rect 457438 22108 457444 22120
rect 457496 22108 457502 22160
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 514846 22080 514852 22092
rect 3200 22052 514852 22080
rect 3200 22040 3206 22052
rect 514846 22040 514852 22052
rect 514904 22040 514910 22092
rect 89809 21947 89867 21953
rect 89809 21913 89821 21947
rect 89855 21944 89867 21947
rect 89990 21944 89996 21956
rect 89855 21916 89996 21944
rect 89855 21913 89867 21916
rect 89809 21907 89867 21913
rect 89990 21904 89996 21916
rect 90048 21904 90054 21956
rect 297910 21428 297916 21480
rect 297968 21468 297974 21480
rect 576854 21468 576860 21480
rect 297968 21440 576860 21468
rect 297968 21428 297974 21440
rect 576854 21428 576860 21440
rect 576912 21428 576918 21480
rect 95142 21360 95148 21412
rect 95200 21400 95206 21412
rect 473354 21400 473360 21412
rect 95200 21372 473360 21400
rect 95200 21360 95206 21372
rect 473354 21360 473360 21372
rect 473412 21360 473418 21412
rect 478690 21360 478696 21412
rect 478748 21400 478754 21412
rect 484394 21400 484400 21412
rect 478748 21372 484400 21400
rect 478748 21360 478754 21372
rect 484394 21360 484400 21372
rect 484452 21360 484458 21412
rect 282822 20068 282828 20120
rect 282880 20108 282886 20120
rect 531314 20108 531320 20120
rect 282880 20080 531320 20108
rect 282880 20068 282886 20080
rect 531314 20068 531320 20080
rect 531372 20068 531378 20120
rect 79594 20000 79600 20052
rect 79652 20040 79658 20052
rect 338206 20040 338212 20052
rect 79652 20012 338212 20040
rect 79652 20000 79658 20012
rect 338206 20000 338212 20012
rect 338264 20000 338270 20052
rect 449158 20000 449164 20052
rect 449216 20040 449222 20052
rect 452562 20040 452568 20052
rect 449216 20012 452568 20040
rect 449216 20000 449222 20012
rect 452562 20000 452568 20012
rect 452620 20000 452626 20052
rect 21910 19932 21916 19984
rect 21968 19972 21974 19984
rect 117958 19972 117964 19984
rect 21968 19944 117964 19972
rect 21968 19932 21974 19944
rect 117958 19932 117964 19944
rect 118016 19932 118022 19984
rect 122742 19932 122748 19984
rect 122800 19972 122806 19984
rect 169754 19972 169760 19984
rect 122800 19944 169760 19972
rect 122800 19932 122806 19944
rect 169754 19932 169760 19944
rect 169812 19932 169818 19984
rect 173710 19932 173716 19984
rect 173768 19972 173774 19984
rect 456794 19972 456800 19984
rect 173768 19944 456800 19972
rect 173768 19932 173774 19944
rect 456794 19932 456800 19944
rect 456852 19932 456858 19984
rect 445570 19320 445576 19372
rect 445628 19360 445634 19372
rect 445662 19360 445668 19372
rect 445628 19332 445668 19360
rect 445628 19320 445634 19332
rect 445662 19320 445668 19332
rect 445720 19320 445726 19372
rect 144730 19292 144736 19304
rect 144691 19264 144736 19292
rect 144730 19252 144736 19264
rect 144788 19252 144794 19304
rect 176838 19292 176844 19304
rect 176799 19264 176844 19292
rect 176838 19252 176844 19264
rect 176896 19252 176902 19304
rect 210973 19295 211031 19301
rect 210973 19261 210985 19295
rect 211019 19292 211031 19295
rect 211154 19292 211160 19304
rect 211019 19264 211160 19292
rect 211019 19261 211031 19264
rect 210973 19255 211031 19261
rect 211154 19252 211160 19264
rect 211212 19252 211218 19304
rect 212442 19292 212448 19304
rect 212403 19264 212448 19292
rect 212442 19252 212448 19264
rect 212500 19252 212506 19304
rect 333882 19292 333888 19304
rect 333843 19264 333888 19292
rect 333882 19252 333888 19264
rect 333940 19252 333946 19304
rect 333974 19252 333980 19304
rect 334032 19292 334038 19304
rect 334802 19292 334808 19304
rect 334032 19264 334808 19292
rect 334032 19252 334038 19264
rect 334802 19252 334808 19264
rect 334860 19252 334866 19304
rect 338114 19252 338120 19304
rect 338172 19292 338178 19304
rect 389174 19292 389180 19304
rect 338172 19264 338217 19292
rect 389135 19264 389180 19292
rect 338172 19252 338178 19264
rect 389174 19252 389180 19264
rect 389232 19252 389238 19304
rect 391750 19292 391756 19304
rect 391711 19264 391756 19292
rect 391750 19252 391756 19264
rect 391808 19252 391814 19304
rect 411162 19292 411168 19304
rect 411123 19264 411168 19292
rect 411162 19252 411168 19264
rect 411220 19252 411226 19304
rect 414014 19252 414020 19304
rect 414072 19292 414078 19304
rect 414474 19292 414480 19304
rect 414072 19264 414480 19292
rect 414072 19252 414078 19264
rect 414474 19252 414480 19264
rect 414532 19252 414538 19304
rect 117222 18708 117228 18760
rect 117280 18748 117286 18760
rect 136634 18748 136640 18760
rect 117280 18720 136640 18748
rect 117280 18708 117286 18720
rect 136634 18708 136640 18720
rect 136692 18708 136698 18760
rect 364242 18708 364248 18760
rect 364300 18748 364306 18760
rect 546586 18748 546592 18760
rect 364300 18720 546592 18748
rect 364300 18708 364306 18720
rect 546586 18708 546592 18720
rect 546644 18708 546650 18760
rect 80790 18640 80796 18692
rect 80848 18680 80854 18692
rect 502334 18680 502340 18692
rect 80848 18652 502340 18680
rect 80848 18640 80854 18652
rect 502334 18640 502340 18652
rect 502392 18640 502398 18692
rect 37182 18572 37188 18624
rect 37240 18612 37246 18624
rect 64138 18612 64144 18624
rect 37240 18584 64144 18612
rect 37240 18572 37246 18584
rect 64138 18572 64144 18584
rect 64196 18572 64202 18624
rect 85482 18572 85488 18624
rect 85540 18612 85546 18624
rect 509418 18612 509424 18624
rect 85540 18584 509424 18612
rect 85540 18572 85546 18584
rect 509418 18572 509424 18584
rect 509476 18572 509482 18624
rect 547138 17960 547144 18012
rect 547196 18000 547202 18012
rect 549254 18000 549260 18012
rect 547196 17972 549260 18000
rect 547196 17960 547202 17972
rect 549254 17960 549260 17972
rect 549312 17960 549318 18012
rect 563698 17892 563704 17944
rect 563756 17932 563762 17944
rect 579798 17932 579804 17944
rect 563756 17904 579804 17932
rect 563756 17892 563762 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 231762 17348 231768 17400
rect 231820 17388 231826 17400
rect 365714 17388 365720 17400
rect 231820 17360 365720 17388
rect 231820 17348 231826 17360
rect 365714 17348 365720 17360
rect 365772 17348 365778 17400
rect 450538 17348 450544 17400
rect 450596 17388 450602 17400
rect 455322 17388 455328 17400
rect 450596 17360 455328 17388
rect 450596 17348 450602 17360
rect 455322 17348 455328 17360
rect 455380 17348 455386 17400
rect 125502 17280 125508 17332
rect 125560 17320 125566 17332
rect 452654 17320 452660 17332
rect 125560 17292 452660 17320
rect 125560 17280 125566 17292
rect 452654 17280 452660 17292
rect 452712 17280 452718 17332
rect 91002 17212 91008 17264
rect 91060 17252 91066 17264
rect 518986 17252 518992 17264
rect 91060 17224 518992 17252
rect 91060 17212 91066 17224
rect 518986 17212 518992 17224
rect 519044 17212 519050 17264
rect 202782 16056 202788 16108
rect 202840 16096 202846 16108
rect 368474 16096 368480 16108
rect 202840 16068 368480 16096
rect 202840 16056 202846 16068
rect 368474 16056 368480 16068
rect 368532 16056 368538 16108
rect 384942 16056 384948 16108
rect 385000 16096 385006 16108
rect 459554 16096 459560 16108
rect 385000 16068 459560 16096
rect 385000 16056 385006 16068
rect 459554 16056 459560 16068
rect 459612 16056 459618 16108
rect 115842 15988 115848 16040
rect 115900 16028 115906 16040
rect 186314 16028 186320 16040
rect 115900 16000 186320 16028
rect 115900 15988 115906 16000
rect 186314 15988 186320 16000
rect 186372 15988 186378 16040
rect 193122 15988 193128 16040
rect 193180 16028 193186 16040
rect 397454 16028 397460 16040
rect 193180 16000 397460 16028
rect 193180 15988 193186 16000
rect 397454 15988 397460 16000
rect 397512 15988 397518 16040
rect 59262 15920 59268 15972
rect 59320 15960 59326 15972
rect 233234 15960 233240 15972
rect 59320 15932 233240 15960
rect 59320 15920 59326 15932
rect 233234 15920 233240 15932
rect 233292 15920 233298 15972
rect 286962 15920 286968 15972
rect 287020 15960 287026 15972
rect 502794 15960 502800 15972
rect 287020 15932 502800 15960
rect 287020 15920 287026 15932
rect 502794 15920 502800 15932
rect 502852 15920 502858 15972
rect 39942 15852 39948 15904
rect 40000 15892 40006 15904
rect 327718 15892 327724 15904
rect 40000 15864 327724 15892
rect 40000 15852 40006 15864
rect 327718 15852 327724 15864
rect 327776 15852 327782 15904
rect 412542 15852 412548 15904
rect 412600 15892 412606 15904
rect 427814 15892 427820 15904
rect 412600 15864 427820 15892
rect 412600 15852 412606 15864
rect 427814 15852 427820 15864
rect 427872 15852 427878 15904
rect 448422 15852 448428 15904
rect 448480 15892 448486 15904
rect 525794 15892 525800 15904
rect 448480 15864 525800 15892
rect 448480 15852 448486 15864
rect 525794 15852 525800 15864
rect 525852 15852 525858 15904
rect 56502 15172 56508 15224
rect 56560 15212 56566 15224
rect 57238 15212 57244 15224
rect 56560 15184 57244 15212
rect 56560 15172 56566 15184
rect 57238 15172 57244 15184
rect 57296 15172 57302 15224
rect 288342 14968 288348 15020
rect 288400 15008 288406 15020
rect 310514 15008 310520 15020
rect 288400 14980 310520 15008
rect 288400 14968 288406 14980
rect 310514 14968 310520 14980
rect 310572 14968 310578 15020
rect 92382 14900 92388 14952
rect 92440 14940 92446 14952
rect 186958 14940 186964 14952
rect 92440 14912 186964 14940
rect 92440 14900 92446 14912
rect 186958 14900 186964 14912
rect 187016 14900 187022 14952
rect 204162 14900 204168 14952
rect 204220 14940 204226 14952
rect 351914 14940 351920 14952
rect 204220 14912 351920 14940
rect 204220 14900 204226 14912
rect 351914 14900 351920 14912
rect 351972 14900 351978 14952
rect 63126 14832 63132 14884
rect 63184 14872 63190 14884
rect 371234 14872 371240 14884
rect 63184 14844 371240 14872
rect 63184 14832 63190 14844
rect 371234 14832 371240 14844
rect 371292 14832 371298 14884
rect 375282 14832 375288 14884
rect 375340 14872 375346 14884
rect 528646 14872 528652 14884
rect 375340 14844 528652 14872
rect 375340 14832 375346 14844
rect 528646 14832 528652 14844
rect 528704 14832 528710 14884
rect 72694 14764 72700 14816
rect 72752 14804 72758 14816
rect 412634 14804 412640 14816
rect 72752 14776 412640 14804
rect 72752 14764 72758 14776
rect 412634 14764 412640 14776
rect 412692 14764 412698 14816
rect 158622 14696 158628 14748
rect 158680 14736 158686 14748
rect 503714 14736 503720 14748
rect 158680 14708 503720 14736
rect 158680 14696 158686 14708
rect 503714 14696 503720 14708
rect 503772 14696 503778 14748
rect 64598 14628 64604 14680
rect 64656 14668 64662 14680
rect 416774 14668 416780 14680
rect 64656 14640 416780 14668
rect 64656 14628 64662 14640
rect 416774 14628 416780 14640
rect 416832 14628 416838 14680
rect 73890 14560 73896 14612
rect 73948 14600 73954 14612
rect 427814 14600 427820 14612
rect 73948 14572 427820 14600
rect 73948 14560 73954 14572
rect 427814 14560 427820 14572
rect 427872 14560 427878 14612
rect 57790 14492 57796 14544
rect 57848 14532 57854 14544
rect 459554 14532 459560 14544
rect 57848 14504 459560 14532
rect 57848 14492 57854 14504
rect 459554 14492 459560 14504
rect 459612 14492 459618 14544
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 37918 14464 37924 14476
rect 11020 14436 37924 14464
rect 11020 14424 11026 14436
rect 37918 14424 37924 14436
rect 37976 14424 37982 14476
rect 68738 14424 68744 14476
rect 68796 14464 68802 14476
rect 560294 14464 560300 14476
rect 68796 14436 560300 14464
rect 68796 14424 68802 14436
rect 560294 14424 560300 14436
rect 560352 14424 560358 14476
rect 345014 13812 345020 13864
rect 345072 13852 345078 13864
rect 351178 13852 351184 13864
rect 345072 13824 351184 13852
rect 345072 13812 345078 13824
rect 351178 13812 351184 13824
rect 351236 13812 351242 13864
rect 72878 13064 72884 13116
rect 72936 13104 72942 13116
rect 124858 13104 124864 13116
rect 72936 13076 124864 13104
rect 72936 13064 72942 13076
rect 124858 13064 124864 13076
rect 124916 13064 124922 13116
rect 126882 13064 126888 13116
rect 126940 13104 126946 13116
rect 293954 13104 293960 13116
rect 126940 13076 293960 13104
rect 126940 13064 126946 13076
rect 293954 13064 293960 13076
rect 294012 13064 294018 13116
rect 426342 13064 426348 13116
rect 426400 13104 426406 13116
rect 500954 13104 500960 13116
rect 426400 13076 500960 13104
rect 426400 13064 426406 13076
rect 500954 13064 500960 13076
rect 501012 13064 501018 13116
rect 488169 12495 488227 12501
rect 488169 12461 488181 12495
rect 488215 12492 488227 12495
rect 488442 12492 488448 12504
rect 488215 12464 488448 12492
rect 488215 12461 488227 12464
rect 488169 12455 488227 12461
rect 488442 12452 488448 12464
rect 488500 12452 488506 12504
rect 65702 12384 65708 12436
rect 65760 12424 65766 12436
rect 142062 12424 142068 12436
rect 65760 12396 142068 12424
rect 65760 12384 65766 12396
rect 142062 12384 142068 12396
rect 142120 12384 142126 12436
rect 169754 12384 169760 12436
rect 169812 12424 169818 12436
rect 170582 12424 170588 12436
rect 169812 12396 170588 12424
rect 169812 12384 169818 12396
rect 170582 12384 170588 12396
rect 170640 12384 170646 12436
rect 204254 12384 204260 12436
rect 204312 12424 204318 12436
rect 205082 12424 205088 12436
rect 204312 12396 205088 12424
rect 204312 12384 204318 12396
rect 205082 12384 205088 12396
rect 205140 12384 205146 12436
rect 212534 12384 212540 12436
rect 212592 12424 212598 12436
rect 213454 12424 213460 12436
rect 212592 12396 213460 12424
rect 212592 12384 212598 12396
rect 213454 12384 213460 12396
rect 213512 12384 213518 12436
rect 213914 12384 213920 12436
rect 213972 12424 213978 12436
rect 214650 12424 214656 12436
rect 213972 12396 214656 12424
rect 213972 12384 213978 12396
rect 214650 12384 214656 12396
rect 214708 12384 214714 12436
rect 280246 12384 280252 12436
rect 280304 12424 280310 12436
rect 281166 12424 281172 12436
rect 280304 12396 281172 12424
rect 280304 12384 280310 12396
rect 281166 12384 281172 12396
rect 281224 12384 281230 12436
rect 281534 12384 281540 12436
rect 281592 12424 281598 12436
rect 282454 12424 282460 12436
rect 281592 12396 282460 12424
rect 281592 12384 281598 12396
rect 282454 12384 282460 12396
rect 282512 12384 282518 12436
rect 335354 12384 335360 12436
rect 335412 12424 335418 12436
rect 335906 12424 335912 12436
rect 335412 12396 335912 12424
rect 335412 12384 335418 12396
rect 335906 12384 335912 12396
rect 335964 12384 335970 12436
rect 350626 12384 350632 12436
rect 350684 12424 350690 12436
rect 351362 12424 351368 12436
rect 350684 12396 351368 12424
rect 350684 12384 350690 12396
rect 351362 12384 351368 12396
rect 351420 12384 351426 12436
rect 351914 12384 351920 12436
rect 351972 12424 351978 12436
rect 352558 12424 352564 12436
rect 351972 12396 352564 12424
rect 351972 12384 351978 12396
rect 352558 12384 352564 12396
rect 352616 12384 352622 12436
rect 404354 12384 404360 12436
rect 404412 12424 404418 12436
rect 404906 12424 404912 12436
rect 404412 12396 404912 12424
rect 404412 12384 404418 12396
rect 404906 12384 404912 12396
rect 404964 12384 404970 12436
rect 412634 12384 412640 12436
rect 412692 12424 412698 12436
rect 413278 12424 413284 12436
rect 412692 12396 413284 12424
rect 412692 12384 412698 12396
rect 413278 12384 413284 12396
rect 413336 12384 413342 12436
rect 448514 12384 448520 12436
rect 448572 12424 448578 12436
rect 448974 12424 448980 12436
rect 448572 12396 448980 12424
rect 448572 12384 448578 12396
rect 448974 12384 448980 12396
rect 449032 12384 449038 12436
rect 454034 12384 454040 12436
rect 454092 12424 454098 12436
rect 454862 12424 454868 12436
rect 454092 12396 454868 12424
rect 454092 12384 454098 12396
rect 454862 12384 454868 12396
rect 454920 12384 454926 12436
rect 473354 12384 473360 12436
rect 473412 12424 473418 12436
rect 473906 12424 473912 12436
rect 473412 12396 473912 12424
rect 473412 12384 473418 12396
rect 473906 12384 473912 12396
rect 473964 12384 473970 12436
rect 486878 12384 486884 12436
rect 486936 12424 486942 12436
rect 487062 12424 487068 12436
rect 486936 12396 487068 12424
rect 486936 12384 486942 12396
rect 487062 12384 487068 12396
rect 487120 12384 487126 12436
rect 502334 12384 502340 12436
rect 502392 12424 502398 12436
rect 502518 12424 502524 12436
rect 502392 12396 502524 12424
rect 502392 12384 502398 12396
rect 502518 12384 502524 12396
rect 502576 12384 502582 12436
rect 81250 12316 81256 12368
rect 81308 12356 81314 12368
rect 229094 12356 229100 12368
rect 81308 12328 229100 12356
rect 81308 12316 81314 12328
rect 229094 12316 229100 12328
rect 229152 12316 229158 12368
rect 61930 12248 61936 12300
rect 61988 12288 61994 12300
rect 260834 12288 260840 12300
rect 61988 12260 260840 12288
rect 61988 12248 61994 12260
rect 260834 12248 260840 12260
rect 260892 12248 260898 12300
rect 63310 12180 63316 12232
rect 63368 12220 63374 12232
rect 269114 12220 269120 12232
rect 63368 12192 269120 12220
rect 63368 12180 63374 12192
rect 269114 12180 269120 12192
rect 269172 12180 269178 12232
rect 68462 12112 68468 12164
rect 68520 12152 68526 12164
rect 276474 12152 276480 12164
rect 68520 12124 276480 12152
rect 68520 12112 68526 12124
rect 276474 12112 276480 12124
rect 276532 12112 276538 12164
rect 61562 12044 61568 12096
rect 61620 12084 61626 12096
rect 372614 12084 372620 12096
rect 61620 12056 372620 12084
rect 61620 12044 61626 12056
rect 372614 12044 372620 12056
rect 372672 12044 372678 12096
rect 61654 11976 61660 12028
rect 61712 12016 61718 12028
rect 472710 12016 472716 12028
rect 61712 11988 472716 12016
rect 61712 11976 61718 11988
rect 472710 11976 472716 11988
rect 472768 11976 472774 12028
rect 46750 11908 46756 11960
rect 46808 11948 46814 11960
rect 465074 11948 465080 11960
rect 46808 11920 465080 11948
rect 46808 11908 46814 11920
rect 465074 11908 465080 11920
rect 465132 11908 465138 11960
rect 50982 11840 50988 11892
rect 51040 11880 51046 11892
rect 494698 11880 494704 11892
rect 51040 11852 494704 11880
rect 51040 11840 51046 11852
rect 494698 11840 494704 11852
rect 494756 11840 494762 11892
rect 511350 11840 511356 11892
rect 511408 11880 511414 11892
rect 571334 11880 571340 11892
rect 511408 11852 571340 11880
rect 511408 11840 511414 11852
rect 571334 11840 571340 11852
rect 571392 11840 571398 11892
rect 64506 11772 64512 11824
rect 64564 11812 64570 11824
rect 516318 11812 516324 11824
rect 64564 11784 516324 11812
rect 64564 11772 64570 11784
rect 516318 11772 516324 11784
rect 516376 11772 516382 11824
rect 65886 11704 65892 11756
rect 65944 11744 65950 11756
rect 529934 11744 529940 11756
rect 65944 11716 529940 11744
rect 65944 11704 65950 11716
rect 529934 11704 529940 11716
rect 529992 11704 529998 11756
rect 457438 10956 457444 11008
rect 457496 10996 457502 11008
rect 462958 10996 462964 11008
rect 457496 10968 462964 10996
rect 457496 10956 457502 10968
rect 462958 10956 462964 10968
rect 463016 10956 463022 11008
rect 77110 10412 77116 10464
rect 77168 10452 77174 10464
rect 253934 10452 253940 10464
rect 77168 10424 253940 10452
rect 77168 10412 77174 10424
rect 253934 10412 253940 10424
rect 253992 10412 253998 10464
rect 34422 10344 34428 10396
rect 34480 10384 34486 10396
rect 350534 10384 350540 10396
rect 34480 10356 350540 10384
rect 34480 10344 34486 10356
rect 350534 10344 350540 10356
rect 350592 10344 350598 10396
rect 17862 10276 17868 10328
rect 17920 10316 17926 10328
rect 437474 10316 437480 10328
rect 17920 10288 437480 10316
rect 17920 10276 17926 10288
rect 437474 10276 437480 10288
rect 437532 10276 437538 10328
rect 411162 9772 411168 9784
rect 411123 9744 411168 9772
rect 411162 9732 411168 9744
rect 411220 9732 411226 9784
rect 140774 9704 140780 9716
rect 140735 9676 140780 9704
rect 140774 9664 140780 9676
rect 140832 9664 140838 9716
rect 144730 9704 144736 9716
rect 144691 9676 144736 9704
rect 144730 9664 144736 9676
rect 144788 9664 144794 9716
rect 176841 9707 176899 9713
rect 176841 9673 176853 9707
rect 176887 9704 176899 9707
rect 176930 9704 176936 9716
rect 176887 9676 176936 9704
rect 176887 9673 176899 9676
rect 176841 9667 176899 9673
rect 176930 9664 176936 9676
rect 176988 9664 176994 9716
rect 212442 9704 212448 9716
rect 212403 9676 212448 9704
rect 212442 9664 212448 9676
rect 212500 9664 212506 9716
rect 333882 9704 333888 9716
rect 333843 9676 333888 9704
rect 333882 9664 333888 9676
rect 333940 9664 333946 9716
rect 338117 9707 338175 9713
rect 338117 9673 338129 9707
rect 338163 9704 338175 9707
rect 338298 9704 338304 9716
rect 338163 9676 338304 9704
rect 338163 9673 338175 9676
rect 338117 9667 338175 9673
rect 338298 9664 338304 9676
rect 338356 9664 338362 9716
rect 389177 9707 389235 9713
rect 389177 9673 389189 9707
rect 389223 9704 389235 9707
rect 389450 9704 389456 9716
rect 389223 9676 389456 9704
rect 389223 9673 389235 9676
rect 389177 9667 389235 9673
rect 389450 9664 389456 9676
rect 389508 9664 389514 9716
rect 391753 9707 391811 9713
rect 391753 9673 391765 9707
rect 391799 9704 391811 9707
rect 391842 9704 391848 9716
rect 391799 9676 391848 9704
rect 391799 9673 391811 9676
rect 391753 9667 391811 9673
rect 391842 9664 391848 9676
rect 391900 9664 391906 9716
rect 488166 9704 488172 9716
rect 488127 9676 488172 9704
rect 488166 9664 488172 9676
rect 488224 9664 488230 9716
rect 512454 9704 512460 9716
rect 512415 9676 512460 9704
rect 512454 9664 512460 9676
rect 512512 9664 512518 9716
rect 61470 9596 61476 9648
rect 61528 9636 61534 9648
rect 121822 9636 121828 9648
rect 61528 9608 121828 9636
rect 61528 9596 61534 9608
rect 121822 9596 121828 9608
rect 121880 9596 121886 9648
rect 410889 9639 410947 9645
rect 410889 9605 410901 9639
rect 410935 9636 410947 9639
rect 411162 9636 411168 9648
rect 410935 9608 411168 9636
rect 410935 9605 410947 9608
rect 410889 9599 410947 9605
rect 411162 9596 411168 9608
rect 411220 9596 411226 9648
rect 502429 9639 502487 9645
rect 502429 9605 502441 9639
rect 502475 9636 502487 9639
rect 502518 9636 502524 9648
rect 502475 9608 502524 9636
rect 502475 9605 502487 9608
rect 502429 9599 502487 9605
rect 502518 9596 502524 9608
rect 502576 9596 502582 9648
rect 64782 9528 64788 9580
rect 64840 9568 64846 9580
rect 190822 9568 190828 9580
rect 64840 9540 190828 9568
rect 64840 9528 64846 9540
rect 190822 9528 190828 9540
rect 190880 9528 190886 9580
rect 445662 9568 445668 9580
rect 445623 9540 445668 9568
rect 445662 9528 445668 9540
rect 445720 9528 445726 9580
rect 59078 9460 59084 9512
rect 59136 9500 59142 9512
rect 206278 9500 206284 9512
rect 59136 9472 206284 9500
rect 59136 9460 59142 9472
rect 206278 9460 206284 9472
rect 206336 9460 206342 9512
rect 63402 9392 63408 9444
rect 63460 9432 63466 9444
rect 279970 9432 279976 9444
rect 63460 9404 279976 9432
rect 63460 9392 63466 9404
rect 279970 9392 279976 9404
rect 280028 9392 280034 9444
rect 113542 9324 113548 9376
rect 113600 9364 113606 9376
rect 336734 9364 336740 9376
rect 113600 9336 336740 9364
rect 113600 9324 113606 9336
rect 336734 9324 336740 9336
rect 336792 9324 336798 9376
rect 60458 9256 60464 9308
rect 60516 9296 60522 9308
rect 290734 9296 290740 9308
rect 60516 9268 290740 9296
rect 60516 9256 60522 9268
rect 290734 9256 290740 9268
rect 290792 9256 290798 9308
rect 65610 9188 65616 9240
rect 65668 9228 65674 9240
rect 244366 9228 244372 9240
rect 65668 9200 244372 9228
rect 65668 9188 65674 9200
rect 244366 9188 244372 9200
rect 244424 9188 244430 9240
rect 273162 9188 273168 9240
rect 273220 9228 273226 9240
rect 510798 9228 510804 9240
rect 273220 9200 510804 9228
rect 273220 9188 273226 9200
rect 510798 9188 510804 9200
rect 510856 9188 510862 9240
rect 68554 9120 68560 9172
rect 68612 9160 68618 9172
rect 308582 9160 308588 9172
rect 68612 9132 308588 9160
rect 68612 9120 68618 9132
rect 308582 9120 308588 9132
rect 308640 9120 308646 9172
rect 30190 9052 30196 9104
rect 30248 9092 30254 9104
rect 286318 9092 286324 9104
rect 30248 9064 286324 9092
rect 30248 9052 30254 9064
rect 286318 9052 286324 9064
rect 286376 9052 286382 9104
rect 444190 9052 444196 9104
rect 444248 9092 444254 9104
rect 518894 9092 518900 9104
rect 444248 9064 518900 9092
rect 444248 9052 444254 9064
rect 518894 9052 518900 9064
rect 518952 9052 518958 9104
rect 70026 8984 70032 9036
rect 70084 9024 70090 9036
rect 340690 9024 340696 9036
rect 70084 8996 340696 9024
rect 70084 8984 70090 8996
rect 340690 8984 340696 8996
rect 340748 8984 340754 9036
rect 376386 8984 376392 9036
rect 376444 9024 376450 9036
rect 512086 9024 512092 9036
rect 376444 8996 512092 9024
rect 376444 8984 376450 8996
rect 512086 8984 512092 8996
rect 512144 8984 512150 9036
rect 71222 8916 71228 8968
rect 71280 8956 71286 8968
rect 358538 8956 358544 8968
rect 71280 8928 358544 8956
rect 71280 8916 71286 8928
rect 358538 8916 358544 8928
rect 358596 8916 358602 8968
rect 382366 8916 382372 8968
rect 382424 8956 382430 8968
rect 521654 8956 521660 8968
rect 382424 8928 521660 8956
rect 382424 8916 382430 8928
rect 521654 8916 521660 8928
rect 521712 8916 521718 8968
rect 540238 8916 540244 8968
rect 540296 8956 540302 8968
rect 573818 8956 573824 8968
rect 540296 8928 573824 8956
rect 540296 8916 540302 8928
rect 573818 8916 573824 8928
rect 573876 8916 573882 8968
rect 462314 8848 462320 8900
rect 462372 8888 462378 8900
rect 465718 8888 465724 8900
rect 462372 8860 465724 8888
rect 462372 8848 462378 8860
rect 465718 8848 465724 8860
rect 465776 8848 465782 8900
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 513742 8276 513748 8288
rect 3476 8248 513748 8276
rect 3476 8236 3482 8248
rect 513742 8236 513748 8248
rect 513800 8236 513806 8288
rect 54018 7624 54024 7676
rect 54076 7664 54082 7676
rect 299474 7664 299480 7676
rect 54076 7636 299480 7664
rect 54076 7624 54082 7636
rect 299474 7624 299480 7636
rect 299532 7624 299538 7676
rect 331214 7624 331220 7676
rect 331272 7664 331278 7676
rect 332410 7664 332416 7676
rect 331272 7636 332416 7664
rect 331272 7624 331278 7636
rect 332410 7624 332416 7636
rect 332468 7624 332474 7676
rect 408494 7624 408500 7676
rect 408552 7664 408558 7676
rect 409690 7664 409696 7676
rect 408552 7636 409696 7664
rect 408552 7624 408558 7636
rect 409690 7624 409696 7636
rect 409748 7624 409754 7676
rect 416774 7624 416780 7676
rect 416832 7664 416838 7676
rect 417970 7664 417976 7676
rect 416832 7636 417976 7664
rect 416832 7624 416838 7636
rect 417970 7624 417976 7636
rect 418028 7624 418034 7676
rect 447410 7624 447416 7676
rect 447468 7664 447474 7676
rect 449158 7664 449164 7676
rect 447468 7636 449164 7664
rect 447468 7624 447474 7636
rect 449158 7624 449164 7636
rect 449216 7624 449222 7676
rect 117130 7556 117136 7608
rect 117188 7596 117194 7608
rect 149698 7596 149704 7608
rect 117188 7568 149704 7596
rect 117188 7556 117194 7568
rect 149698 7556 149704 7568
rect 149756 7556 149762 7608
rect 178954 7556 178960 7608
rect 179012 7596 179018 7608
rect 442994 7596 443000 7608
rect 179012 7568 443000 7596
rect 179012 7556 179018 7568
rect 442994 7556 443000 7568
rect 443052 7556 443058 7608
rect 451274 7556 451280 7608
rect 451332 7596 451338 7608
rect 452470 7596 452476 7608
rect 451332 7568 452476 7596
rect 451332 7556 451338 7568
rect 452470 7556 452476 7568
rect 452528 7556 452534 7608
rect 494054 7556 494060 7608
rect 494112 7596 494118 7608
rect 495342 7596 495348 7608
rect 494112 7568 495348 7596
rect 494112 7556 494118 7568
rect 495342 7556 495348 7568
rect 495400 7556 495406 7608
rect 552750 7556 552756 7608
rect 552808 7596 552814 7608
rect 564342 7596 564348 7608
rect 552808 7568 564348 7596
rect 552808 7556 552814 7568
rect 564342 7556 564348 7568
rect 564400 7556 564406 7608
rect 201494 7488 201500 7540
rect 201552 7528 201558 7540
rect 202690 7528 202696 7540
rect 201552 7500 202696 7528
rect 201552 7488 201558 7500
rect 202690 7488 202696 7500
rect 202748 7488 202754 7540
rect 71130 6808 71136 6860
rect 71188 6848 71194 6860
rect 153930 6848 153936 6860
rect 71188 6820 153936 6848
rect 71188 6808 71194 6820
rect 153930 6808 153936 6820
rect 153988 6808 153994 6860
rect 60550 6740 60556 6792
rect 60608 6780 60614 6792
rect 159910 6780 159916 6792
rect 60608 6752 159916 6780
rect 60608 6740 60614 6752
rect 159910 6740 159916 6752
rect 159968 6740 159974 6792
rect 72418 6672 72424 6724
rect 72476 6712 72482 6724
rect 183738 6712 183744 6724
rect 72476 6684 183744 6712
rect 72476 6672 72482 6684
rect 183738 6672 183744 6684
rect 183796 6672 183802 6724
rect 445665 6715 445723 6721
rect 445665 6681 445677 6715
rect 445711 6712 445723 6715
rect 475102 6712 475108 6724
rect 445711 6684 475108 6712
rect 445711 6681 445723 6684
rect 445665 6675 445723 6681
rect 475102 6672 475108 6684
rect 475160 6672 475166 6724
rect 481082 6672 481088 6724
rect 481140 6712 481146 6724
rect 515214 6712 515220 6724
rect 481140 6684 515220 6712
rect 481140 6672 481146 6684
rect 515214 6672 515220 6684
rect 515272 6672 515278 6724
rect 68922 6604 68928 6656
rect 68980 6644 68986 6656
rect 125410 6644 125416 6656
rect 68980 6616 125416 6644
rect 68980 6604 68986 6616
rect 125410 6604 125416 6616
rect 125468 6604 125474 6656
rect 138474 6604 138480 6656
rect 138532 6644 138538 6656
rect 256694 6644 256700 6656
rect 138532 6616 256700 6644
rect 138532 6604 138538 6616
rect 256694 6604 256700 6616
rect 256752 6604 256758 6656
rect 406102 6604 406108 6656
rect 406160 6644 406166 6656
rect 434714 6644 434720 6656
rect 406160 6616 434720 6644
rect 406160 6604 406166 6616
rect 434714 6604 434720 6616
rect 434772 6604 434778 6656
rect 459646 6604 459652 6656
rect 459704 6644 459710 6656
rect 510614 6644 510620 6656
rect 459704 6616 510620 6644
rect 459704 6604 459710 6616
rect 510614 6604 510620 6616
rect 510672 6604 510678 6656
rect 70670 6536 70676 6588
rect 70728 6576 70734 6588
rect 225598 6576 225604 6588
rect 70728 6548 225604 6576
rect 70728 6536 70734 6548
rect 225598 6536 225604 6548
rect 225656 6536 225662 6588
rect 229002 6536 229008 6588
rect 229060 6576 229066 6588
rect 416866 6576 416872 6588
rect 229060 6548 416872 6576
rect 229060 6536 229066 6548
rect 416866 6536 416872 6548
rect 416924 6536 416930 6588
rect 447778 6536 447784 6588
rect 447836 6576 447842 6588
rect 514754 6576 514760 6588
rect 447836 6548 514760 6576
rect 447836 6536 447842 6548
rect 514754 6536 514760 6548
rect 514812 6536 514818 6588
rect 67358 6468 67364 6520
rect 67416 6508 67422 6520
rect 258626 6508 258632 6520
rect 67416 6480 258632 6508
rect 67416 6468 67422 6480
rect 258626 6468 258632 6480
rect 258684 6468 258690 6520
rect 263502 6468 263508 6520
rect 263560 6508 263566 6520
rect 313366 6508 313372 6520
rect 263560 6480 313372 6508
rect 263560 6468 263566 6480
rect 313366 6468 313372 6480
rect 313424 6468 313430 6520
rect 423950 6468 423956 6520
rect 424008 6508 424014 6520
rect 513558 6508 513564 6520
rect 424008 6480 513564 6508
rect 424008 6468 424014 6480
rect 513558 6468 513564 6480
rect 513616 6468 513622 6520
rect 67542 6400 67548 6452
rect 67600 6440 67606 6452
rect 318058 6440 318064 6452
rect 67600 6412 318064 6440
rect 67600 6400 67606 6412
rect 318058 6400 318064 6412
rect 318116 6400 318122 6452
rect 422754 6400 422760 6452
rect 422812 6440 422818 6452
rect 516226 6440 516232 6452
rect 422812 6412 516232 6440
rect 422812 6400 422818 6412
rect 516226 6400 516232 6412
rect 516284 6400 516290 6452
rect 531958 6400 531964 6452
rect 532016 6440 532022 6452
rect 572622 6440 572628 6452
rect 532016 6412 572628 6440
rect 532016 6400 532022 6412
rect 572622 6400 572628 6412
rect 572680 6400 572686 6452
rect 73982 6332 73988 6384
rect 74040 6372 74046 6384
rect 554866 6372 554872 6384
rect 74040 6344 554872 6372
rect 74040 6332 74046 6344
rect 554866 6332 554872 6344
rect 554924 6332 554930 6384
rect 66070 6264 66076 6316
rect 66128 6304 66134 6316
rect 558362 6304 558368 6316
rect 66128 6276 558368 6304
rect 66128 6264 66134 6276
rect 558362 6264 558368 6276
rect 558420 6264 558426 6316
rect 65978 6196 65984 6248
rect 66036 6236 66042 6248
rect 561950 6236 561956 6248
rect 66036 6208 561956 6236
rect 66036 6196 66042 6208
rect 561950 6196 561956 6208
rect 562008 6196 562014 6248
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 19978 6168 19984 6180
rect 11296 6140 19984 6168
rect 11296 6128 11302 6140
rect 19978 6128 19984 6140
rect 20036 6128 20042 6180
rect 38470 6128 38476 6180
rect 38528 6168 38534 6180
rect 46198 6168 46204 6180
rect 38528 6140 46204 6168
rect 38528 6128 38534 6140
rect 46198 6128 46204 6140
rect 46256 6128 46262 6180
rect 66898 6128 66904 6180
rect 66956 6168 66962 6180
rect 569034 6168 569040 6180
rect 66956 6140 569040 6168
rect 66956 6128 66962 6140
rect 569034 6128 569040 6140
rect 569092 6128 569098 6180
rect 432322 5992 432328 6044
rect 432380 6032 432386 6044
rect 433242 6032 433248 6044
rect 432380 6004 433248 6032
rect 432380 5992 432386 6004
rect 433242 5992 433248 6004
rect 433300 5992 433306 6044
rect 201586 5924 201592 5976
rect 201644 5964 201650 5976
rect 211062 5964 211068 5976
rect 201644 5936 211068 5964
rect 201644 5924 201650 5936
rect 211062 5924 211068 5936
rect 211120 5924 211126 5976
rect 481818 5924 481824 5976
rect 481876 5964 481882 5976
rect 491202 5964 491208 5976
rect 481876 5936 491208 5964
rect 481876 5924 481882 5936
rect 491202 5924 491208 5936
rect 491260 5924 491266 5976
rect 259822 5856 259828 5908
rect 259880 5896 259886 5908
rect 260742 5896 260748 5908
rect 259880 5868 260748 5896
rect 259880 5856 259886 5868
rect 260742 5856 260748 5868
rect 260800 5856 260806 5908
rect 135254 5720 135260 5772
rect 135312 5760 135318 5772
rect 144822 5760 144828 5772
rect 135312 5732 144828 5760
rect 135312 5720 135318 5732
rect 144822 5720 144828 5732
rect 144880 5720 144886 5772
rect 438118 5720 438124 5772
rect 438176 5760 438182 5772
rect 442902 5760 442908 5772
rect 438176 5732 442908 5760
rect 438176 5720 438182 5732
rect 442902 5720 442908 5732
rect 442960 5720 442966 5772
rect 182174 5652 182180 5704
rect 182232 5692 182238 5704
rect 199930 5692 199936 5704
rect 182232 5664 199936 5692
rect 182232 5652 182238 5664
rect 199930 5652 199936 5664
rect 199988 5652 199994 5704
rect 46934 5516 46940 5568
rect 46992 5556 46998 5568
rect 50338 5556 50344 5568
rect 46992 5528 50344 5556
rect 46992 5516 46998 5528
rect 50338 5516 50344 5528
rect 50396 5516 50402 5568
rect 571978 5516 571984 5568
rect 572036 5556 572042 5568
rect 576210 5556 576216 5568
rect 572036 5528 576216 5556
rect 572036 5516 572042 5528
rect 576210 5516 576216 5528
rect 576268 5516 576274 5568
rect 331048 5188 333284 5216
rect 320082 5108 320088 5160
rect 320140 5148 320146 5160
rect 331048 5148 331076 5188
rect 320140 5120 331076 5148
rect 320140 5108 320146 5120
rect 333256 5080 333284 5188
rect 350258 5080 350264 5092
rect 333256 5052 350264 5080
rect 350258 5040 350264 5052
rect 350316 5040 350322 5092
rect 378686 5040 378692 5092
rect 378744 5080 378750 5092
rect 462222 5080 462228 5092
rect 378744 5052 462228 5080
rect 378744 5040 378750 5052
rect 462222 5040 462228 5052
rect 462280 5040 462286 5092
rect 327626 4972 327632 5024
rect 327684 5012 327690 5024
rect 457438 5012 457444 5024
rect 327684 4984 457444 5012
rect 327684 4972 327690 4984
rect 457438 4972 457444 4984
rect 457496 4972 457502 5024
rect 291930 4904 291936 4956
rect 291988 4944 291994 4956
rect 447410 4944 447416 4956
rect 291988 4916 447416 4944
rect 291988 4904 291994 4916
rect 447410 4904 447416 4916
rect 447468 4904 447474 4956
rect 456702 4904 456708 4956
rect 456760 4944 456766 4956
rect 467926 4944 467932 4956
rect 456760 4916 467932 4944
rect 456760 4904 456766 4916
rect 467926 4904 467932 4916
rect 467984 4904 467990 4956
rect 206922 4836 206928 4888
rect 206980 4876 206986 4888
rect 225322 4876 225328 4888
rect 206980 4848 225328 4876
rect 206980 4836 206986 4848
rect 225322 4836 225328 4848
rect 225380 4836 225386 4888
rect 287146 4836 287152 4888
rect 287204 4876 287210 4888
rect 450538 4876 450544 4888
rect 287204 4848 450544 4876
rect 287204 4836 287210 4848
rect 450538 4836 450544 4848
rect 450596 4836 450602 4888
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 14458 4808 14464 4820
rect 6512 4780 14464 4808
rect 6512 4768 6518 4780
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 40954 4768 40960 4820
rect 41012 4808 41018 4820
rect 55858 4808 55864 4820
rect 41012 4780 55864 4808
rect 41012 4768 41018 4780
rect 55858 4768 55864 4780
rect 55916 4768 55922 4820
rect 112346 4768 112352 4820
rect 112404 4808 112410 4820
rect 237374 4808 237380 4820
rect 112404 4780 237380 4808
rect 112404 4768 112410 4780
rect 237374 4768 237380 4780
rect 237432 4768 237438 4820
rect 272886 4768 272892 4820
rect 272944 4808 272950 4820
rect 460198 4808 460204 4820
rect 272944 4780 460204 4808
rect 272944 4768 272950 4780
rect 460198 4768 460204 4780
rect 460256 4768 460262 4820
rect 527818 4768 527824 4820
rect 527876 4808 527882 4820
rect 548886 4808 548892 4820
rect 527876 4780 548892 4808
rect 527876 4768 527882 4780
rect 548886 4768 548892 4780
rect 548944 4768 548950 4820
rect 554038 4768 554044 4820
rect 554096 4808 554102 4820
rect 578602 4808 578608 4820
rect 554096 4780 578608 4808
rect 554096 4768 554102 4780
rect 578602 4768 578608 4780
rect 578660 4768 578666 4820
rect 502426 4632 502432 4684
rect 502484 4672 502490 4684
rect 503622 4672 503628 4684
rect 502484 4644 503628 4672
rect 502484 4632 502490 4644
rect 503622 4632 503628 4644
rect 503680 4632 503686 4684
rect 12434 4360 12440 4412
rect 12492 4400 12498 4412
rect 17218 4400 17224 4412
rect 12492 4372 17224 4400
rect 12492 4360 12498 4372
rect 17218 4360 17224 4372
rect 17276 4360 17282 4412
rect 133690 4156 133696 4208
rect 133748 4196 133754 4208
rect 133748 4168 133920 4196
rect 133748 4156 133754 4168
rect 64414 4088 64420 4140
rect 64472 4128 64478 4140
rect 133782 4128 133788 4140
rect 64472 4100 133788 4128
rect 64472 4088 64478 4100
rect 133782 4088 133788 4100
rect 133840 4088 133846 4140
rect 133892 4128 133920 4168
rect 133892 4100 508636 4128
rect 566 4020 572 4072
rect 624 4060 630 4072
rect 9030 4060 9036 4072
rect 624 4032 9036 4060
rect 624 4020 630 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 64322 4020 64328 4072
rect 64380 4060 64386 4072
rect 80238 4060 80244 4072
rect 64380 4032 80244 4060
rect 64380 4020 64386 4032
rect 80238 4020 80244 4032
rect 80296 4020 80302 4072
rect 84838 4020 84844 4072
rect 84896 4060 84902 4072
rect 93857 4063 93915 4069
rect 93857 4060 93869 4063
rect 84896 4032 93869 4060
rect 84896 4020 84902 4032
rect 93857 4029 93869 4032
rect 93903 4029 93915 4063
rect 93857 4023 93915 4029
rect 103425 4063 103483 4069
rect 103425 4029 103437 4063
rect 103471 4060 103483 4063
rect 113177 4063 113235 4069
rect 113177 4060 113189 4063
rect 103471 4032 113189 4060
rect 103471 4029 103483 4032
rect 103425 4023 103483 4029
rect 113177 4029 113189 4032
rect 113223 4029 113235 4063
rect 113177 4023 113235 4029
rect 122745 4063 122803 4069
rect 122745 4029 122757 4063
rect 122791 4060 122803 4063
rect 132497 4063 132555 4069
rect 132497 4060 132509 4063
rect 122791 4032 132509 4060
rect 122791 4029 122803 4032
rect 122745 4023 122803 4029
rect 132497 4029 132509 4032
rect 132543 4029 132555 4063
rect 132497 4023 132555 4029
rect 142154 4020 142160 4072
rect 142212 4060 142218 4072
rect 143258 4060 143264 4072
rect 142212 4032 143264 4060
rect 142212 4020 142218 4032
rect 143258 4020 143264 4032
rect 143316 4020 143322 4072
rect 145650 4020 145656 4072
rect 145708 4060 145714 4072
rect 146202 4060 146208 4072
rect 145708 4032 146208 4060
rect 145708 4020 145714 4032
rect 146202 4020 146208 4032
rect 146260 4020 146266 4072
rect 146294 4020 146300 4072
rect 146352 4060 146358 4072
rect 146846 4060 146852 4072
rect 146352 4032 146852 4060
rect 146352 4020 146358 4032
rect 146846 4020 146852 4032
rect 146904 4020 146910 4072
rect 146941 4063 146999 4069
rect 146941 4029 146953 4063
rect 146987 4060 146999 4063
rect 157337 4063 157395 4069
rect 157337 4060 157349 4063
rect 146987 4032 157349 4060
rect 146987 4029 146999 4032
rect 146941 4023 146999 4029
rect 157337 4029 157349 4032
rect 157383 4029 157395 4063
rect 157337 4023 157395 4029
rect 157518 4020 157524 4072
rect 157576 4060 157582 4072
rect 158622 4060 158628 4072
rect 157576 4032 158628 4060
rect 157576 4020 157582 4032
rect 158622 4020 158628 4032
rect 158680 4020 158686 4072
rect 166994 4020 167000 4072
rect 167052 4060 167058 4072
rect 168190 4060 168196 4072
rect 167052 4032 168196 4060
rect 167052 4020 167058 4032
rect 168190 4020 168196 4032
rect 168248 4020 168254 4072
rect 176930 4020 176936 4072
rect 176988 4060 176994 4072
rect 177758 4060 177764 4072
rect 176988 4032 177764 4060
rect 176988 4020 176994 4032
rect 177758 4020 177764 4032
rect 177816 4020 177822 4072
rect 179414 4020 179420 4072
rect 179472 4060 179478 4072
rect 180150 4060 180156 4072
rect 179472 4032 180156 4060
rect 179472 4020 179478 4032
rect 180150 4020 180156 4032
rect 180208 4020 180214 4072
rect 197998 4020 198004 4072
rect 198056 4060 198062 4072
rect 198642 4060 198648 4072
rect 198056 4032 198648 4060
rect 198056 4020 198062 4032
rect 198642 4020 198648 4032
rect 198700 4020 198706 4072
rect 199194 4020 199200 4072
rect 199252 4060 199258 4072
rect 200022 4060 200028 4072
rect 199252 4032 200028 4060
rect 199252 4020 199258 4032
rect 200022 4020 200028 4032
rect 200080 4020 200086 4072
rect 201494 4020 201500 4072
rect 201552 4060 201558 4072
rect 202782 4060 202788 4072
rect 201552 4032 202788 4060
rect 201552 4020 201558 4032
rect 202782 4020 202788 4032
rect 202840 4020 202846 4072
rect 207014 4020 207020 4072
rect 207072 4060 207078 4072
rect 207474 4060 207480 4072
rect 207072 4032 207480 4060
rect 207072 4020 207078 4032
rect 207474 4020 207480 4032
rect 207532 4020 207538 4072
rect 208670 4020 208676 4072
rect 208728 4060 208734 4072
rect 209682 4060 209688 4072
rect 208728 4032 209688 4060
rect 208728 4020 208734 4032
rect 209682 4020 209688 4032
rect 209740 4020 209746 4072
rect 209866 4020 209872 4072
rect 209924 4060 209930 4072
rect 210878 4060 210884 4072
rect 209924 4032 210884 4060
rect 209924 4020 209930 4032
rect 210878 4020 210884 4032
rect 210936 4020 210942 4072
rect 217042 4020 217048 4072
rect 217100 4060 217106 4072
rect 217962 4060 217968 4072
rect 217100 4032 217968 4060
rect 217100 4020 217106 4032
rect 217962 4020 217968 4032
rect 218020 4020 218026 4072
rect 218054 4020 218060 4072
rect 218112 4060 218118 4072
rect 219342 4060 219348 4072
rect 218112 4032 219348 4060
rect 218112 4020 218118 4032
rect 219342 4020 219348 4032
rect 219400 4020 219406 4072
rect 274082 4020 274088 4072
rect 274140 4060 274146 4072
rect 274542 4060 274548 4072
rect 274140 4032 274548 4060
rect 274140 4020 274146 4032
rect 274542 4020 274548 4032
rect 274600 4020 274606 4072
rect 275278 4020 275284 4072
rect 275336 4060 275342 4072
rect 275922 4060 275928 4072
rect 275336 4032 275928 4060
rect 275336 4020 275342 4032
rect 275922 4020 275928 4032
rect 275980 4020 275986 4072
rect 278866 4020 278872 4072
rect 278924 4060 278930 4072
rect 280062 4060 280068 4072
rect 278924 4032 280068 4060
rect 278924 4020 278930 4032
rect 280062 4020 280068 4032
rect 280120 4020 280126 4072
rect 331214 4020 331220 4072
rect 331272 4060 331278 4072
rect 332502 4060 332508 4072
rect 331272 4032 332508 4060
rect 331272 4020 331278 4032
rect 332502 4020 332508 4032
rect 332560 4020 332566 4072
rect 337102 4020 337108 4072
rect 337160 4060 337166 4072
rect 338022 4060 338028 4072
rect 337160 4032 338028 4060
rect 337160 4020 337166 4032
rect 338022 4020 338028 4032
rect 338080 4020 338086 4072
rect 356146 4020 356152 4072
rect 356204 4060 356210 4072
rect 357342 4060 357348 4072
rect 356204 4032 357348 4060
rect 356204 4020 356210 4032
rect 357342 4020 357348 4032
rect 357400 4020 357406 4072
rect 397822 4020 397828 4072
rect 397880 4060 397886 4072
rect 398742 4060 398748 4072
rect 397880 4032 398748 4060
rect 397880 4020 397886 4032
rect 398742 4020 398748 4032
rect 398800 4020 398806 4072
rect 399018 4020 399024 4072
rect 399076 4060 399082 4072
rect 400122 4060 400128 4072
rect 399076 4032 400128 4060
rect 399076 4020 399082 4032
rect 400122 4020 400128 4032
rect 400180 4020 400186 4072
rect 408494 4020 408500 4072
rect 408552 4060 408558 4072
rect 409782 4060 409788 4072
rect 408552 4032 409788 4060
rect 408552 4020 408558 4032
rect 409782 4020 409788 4032
rect 409840 4020 409846 4072
rect 412082 4020 412088 4072
rect 412140 4060 412146 4072
rect 412542 4060 412548 4072
rect 412140 4032 412548 4060
rect 412140 4020 412146 4032
rect 412542 4020 412548 4032
rect 412600 4020 412606 4072
rect 456058 4020 456064 4072
rect 456116 4060 456122 4072
rect 456610 4060 456616 4072
rect 456116 4032 456616 4060
rect 456116 4020 456122 4032
rect 456610 4020 456616 4032
rect 456668 4020 456674 4072
rect 466822 4020 466828 4072
rect 466880 4060 466886 4072
rect 467742 4060 467748 4072
rect 466880 4032 467748 4060
rect 466880 4020 466886 4032
rect 467742 4020 467748 4032
rect 467800 4020 467806 4072
rect 485774 4020 485780 4072
rect 485832 4060 485838 4072
rect 486970 4060 486976 4072
rect 485832 4032 486976 4060
rect 485832 4020 485838 4032
rect 486970 4020 486976 4032
rect 487028 4020 487034 4072
rect 498930 4020 498936 4072
rect 498988 4060 498994 4072
rect 499482 4060 499488 4072
rect 498988 4032 499488 4060
rect 498988 4020 498994 4032
rect 499482 4020 499488 4032
rect 499540 4020 499546 4072
rect 503717 4063 503775 4069
rect 503717 4029 503729 4063
rect 503763 4060 503775 4063
rect 508501 4063 508559 4069
rect 508501 4060 508513 4063
rect 503763 4032 508513 4060
rect 503763 4029 503775 4032
rect 503717 4023 503775 4029
rect 508501 4029 508513 4032
rect 508547 4029 508559 4063
rect 508608 4060 508636 4100
rect 511442 4088 511448 4140
rect 511500 4128 511506 4140
rect 513190 4128 513196 4140
rect 511500 4100 513196 4128
rect 511500 4088 511506 4100
rect 513190 4088 513196 4100
rect 513248 4088 513254 4140
rect 512178 4060 512184 4072
rect 508608 4032 512184 4060
rect 508501 4023 508559 4029
rect 512178 4020 512184 4032
rect 512236 4020 512242 4072
rect 69934 3952 69940 4004
rect 69992 3992 69998 4004
rect 150434 3992 150440 4004
rect 69992 3964 150440 3992
rect 69992 3952 69998 3964
rect 150434 3952 150440 3964
rect 150492 3952 150498 4004
rect 470318 3952 470324 4004
rect 470376 3992 470382 4004
rect 494146 3992 494152 4004
rect 470376 3964 494152 3992
rect 470376 3952 470382 3964
rect 494146 3952 494152 3964
rect 494204 3952 494210 4004
rect 497734 3952 497740 4004
rect 497792 3992 497798 4004
rect 517698 3992 517704 4004
rect 497792 3964 517704 3992
rect 497792 3952 497798 3964
rect 517698 3952 517704 3964
rect 517756 3952 517762 4004
rect 68646 3884 68652 3936
rect 68704 3924 68710 3936
rect 162302 3924 162308 3936
rect 68704 3896 162308 3924
rect 68704 3884 68710 3896
rect 162302 3884 162308 3896
rect 162360 3884 162366 3936
rect 477494 3884 477500 3936
rect 477552 3924 477558 3936
rect 496449 3927 496507 3933
rect 496449 3924 496461 3927
rect 477552 3896 496461 3924
rect 477552 3884 477558 3896
rect 496449 3893 496461 3896
rect 496495 3893 496507 3927
rect 496449 3887 496507 3893
rect 500126 3884 500132 3936
rect 500184 3924 500190 3936
rect 500862 3924 500868 3936
rect 500184 3896 500868 3924
rect 500184 3884 500190 3896
rect 500862 3884 500868 3896
rect 500920 3884 500926 3936
rect 508501 3927 508559 3933
rect 508501 3893 508513 3927
rect 508547 3924 508559 3927
rect 513466 3924 513472 3936
rect 508547 3896 513472 3924
rect 508547 3893 508559 3896
rect 508501 3887 508559 3893
rect 513466 3884 513472 3896
rect 513524 3884 513530 3936
rect 64690 3816 64696 3868
rect 64748 3856 64754 3868
rect 165890 3856 165896 3868
rect 64748 3828 165896 3856
rect 64748 3816 64754 3828
rect 165890 3816 165896 3828
rect 165948 3816 165954 3868
rect 257430 3856 257436 3868
rect 251376 3828 257436 3856
rect 60366 3748 60372 3800
rect 60424 3788 60430 3800
rect 167086 3788 167092 3800
rect 60424 3760 167092 3788
rect 60424 3748 60430 3760
rect 167086 3748 167092 3760
rect 167144 3748 167150 3800
rect 66990 3680 66996 3732
rect 67048 3720 67054 3732
rect 73065 3723 73123 3729
rect 73065 3720 73077 3723
rect 67048 3692 73077 3720
rect 67048 3680 67054 3692
rect 73065 3689 73077 3692
rect 73111 3689 73123 3723
rect 73065 3683 73123 3689
rect 74442 3680 74448 3732
rect 74500 3720 74506 3732
rect 251376 3720 251404 3828
rect 257430 3816 257436 3828
rect 257488 3816 257494 3868
rect 375282 3816 375288 3868
rect 375340 3856 375346 3868
rect 406378 3856 406384 3868
rect 375340 3828 406384 3856
rect 375340 3816 375346 3828
rect 406378 3816 406384 3828
rect 406436 3816 406442 3868
rect 431126 3816 431132 3868
rect 431184 3856 431190 3868
rect 439498 3856 439504 3868
rect 431184 3828 439504 3856
rect 431184 3816 431190 3828
rect 439498 3816 439504 3828
rect 439556 3816 439562 3868
rect 442994 3816 443000 3868
rect 443052 3856 443058 3868
rect 502978 3856 502984 3868
rect 443052 3828 502984 3856
rect 443052 3816 443058 3828
rect 502978 3816 502984 3828
rect 503036 3816 503042 3868
rect 300302 3748 300308 3800
rect 300360 3788 300366 3800
rect 378686 3788 378692 3800
rect 300360 3760 378692 3788
rect 300360 3748 300366 3760
rect 378686 3748 378692 3760
rect 378744 3748 378750 3800
rect 401318 3748 401324 3800
rect 401376 3788 401382 3800
rect 512362 3788 512368 3800
rect 401376 3760 512368 3788
rect 401376 3748 401382 3760
rect 512362 3748 512368 3760
rect 512420 3748 512426 3800
rect 74500 3692 251404 3720
rect 74500 3680 74506 3692
rect 270494 3680 270500 3732
rect 270552 3720 270558 3732
rect 513374 3720 513380 3732
rect 270552 3692 513380 3720
rect 270552 3680 270558 3692
rect 513374 3680 513380 3692
rect 513432 3680 513438 3732
rect 63218 3612 63224 3664
rect 63276 3652 63282 3664
rect 222930 3652 222936 3664
rect 63276 3624 222936 3652
rect 63276 3612 63282 3624
rect 222930 3612 222936 3624
rect 222988 3612 222994 3664
rect 227714 3612 227720 3664
rect 227772 3652 227778 3664
rect 228910 3652 228916 3664
rect 227772 3624 228916 3652
rect 227772 3612 227778 3624
rect 228910 3612 228916 3624
rect 228968 3612 228974 3664
rect 235994 3612 236000 3664
rect 236052 3652 236058 3664
rect 237190 3652 237196 3664
rect 236052 3624 237196 3652
rect 236052 3612 236058 3624
rect 237190 3612 237196 3624
rect 237248 3612 237254 3664
rect 252646 3612 252652 3664
rect 252704 3652 252710 3664
rect 253842 3652 253848 3664
rect 252704 3624 253848 3652
rect 252704 3612 252710 3624
rect 253842 3612 253848 3624
rect 253900 3612 253906 3664
rect 253937 3655 253995 3661
rect 253937 3621 253949 3655
rect 253983 3652 253995 3655
rect 520366 3652 520372 3664
rect 253983 3624 520372 3652
rect 253983 3621 253995 3624
rect 253937 3615 253995 3621
rect 520366 3612 520372 3624
rect 520424 3612 520430 3664
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 15838 3584 15844 3596
rect 7708 3556 15844 3584
rect 7708 3544 7714 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21910 3584 21916 3596
rect 20772 3556 21916 3584
rect 20772 3544 20778 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 30282 3584 30288 3596
rect 29144 3556 30288 3584
rect 29144 3544 29150 3556
rect 30282 3544 30288 3556
rect 30340 3544 30346 3596
rect 43346 3544 43352 3596
rect 43404 3584 43410 3596
rect 315298 3584 315304 3596
rect 43404 3556 315304 3584
rect 43404 3544 43410 3556
rect 315298 3544 315304 3556
rect 315356 3544 315362 3596
rect 321646 3544 321652 3596
rect 321704 3584 321710 3596
rect 322842 3584 322848 3596
rect 321704 3556 322848 3584
rect 321704 3544 321710 3556
rect 322842 3544 322848 3556
rect 322900 3544 322906 3596
rect 322934 3544 322940 3596
rect 322992 3584 322998 3596
rect 517606 3584 517612 3596
rect 322992 3556 517612 3584
rect 322992 3544 322998 3556
rect 517606 3544 517612 3556
rect 517664 3544 517670 3596
rect 520274 3544 520280 3596
rect 520332 3584 520338 3596
rect 521470 3584 521476 3596
rect 520332 3556 521476 3584
rect 520332 3544 520338 3556
rect 521470 3544 521476 3556
rect 521528 3544 521534 3596
rect 574738 3544 574744 3596
rect 574796 3544 574802 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17862 3516 17868 3528
rect 17276 3488 17868 3516
rect 17276 3476 17282 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19242 3516 19248 3528
rect 18380 3488 19248 3516
rect 18380 3476 18386 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20622 3516 20628 3528
rect 19576 3488 20628 3516
rect 19576 3476 19582 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 26142 3516 26148 3528
rect 25556 3488 26148 3516
rect 25556 3476 25562 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27522 3516 27528 3528
rect 26752 3488 27528 3516
rect 26752 3476 26758 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 28902 3516 28908 3528
rect 27948 3488 28908 3516
rect 27948 3476 27954 3488
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 33870 3476 33876 3528
rect 33928 3516 33934 3528
rect 34422 3516 34428 3528
rect 33928 3488 34428 3516
rect 33928 3476 33934 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34974 3476 34980 3528
rect 35032 3516 35038 3528
rect 35802 3516 35808 3528
rect 35032 3488 35808 3516
rect 35032 3476 35038 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 37182 3516 37188 3528
rect 36228 3488 37188 3516
rect 36228 3476 36234 3488
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 37366 3476 37372 3528
rect 37424 3516 37430 3528
rect 38562 3516 38568 3528
rect 37424 3488 38568 3516
rect 37424 3476 37430 3488
rect 38562 3476 38568 3488
rect 38620 3476 38626 3528
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 42702 3516 42708 3528
rect 42208 3488 42708 3516
rect 42208 3476 42214 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 44542 3476 44548 3528
rect 44600 3516 44606 3528
rect 45462 3516 45468 3528
rect 44600 3488 45468 3516
rect 44600 3476 44606 3488
rect 45462 3476 45468 3488
rect 45520 3476 45526 3528
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46750 3516 46756 3528
rect 45796 3488 46756 3516
rect 45796 3476 45802 3488
rect 46750 3476 46756 3488
rect 46808 3476 46814 3528
rect 51626 3476 51632 3528
rect 51684 3516 51690 3528
rect 52362 3516 52368 3528
rect 51684 3488 52368 3516
rect 51684 3476 51690 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 52822 3476 52828 3528
rect 52880 3516 52886 3528
rect 53742 3516 53748 3528
rect 52880 3488 53748 3516
rect 52880 3476 52886 3488
rect 53742 3476 53748 3488
rect 53800 3476 53806 3528
rect 59998 3476 60004 3528
rect 60056 3516 60062 3528
rect 60642 3516 60648 3528
rect 60056 3488 60648 3516
rect 60056 3476 60062 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 61194 3476 61200 3528
rect 61252 3516 61258 3528
rect 62022 3516 62028 3528
rect 61252 3488 62028 3516
rect 61252 3476 61258 3488
rect 62022 3476 62028 3488
rect 62080 3476 62086 3528
rect 62390 3476 62396 3528
rect 62448 3516 62454 3528
rect 63034 3516 63040 3528
rect 62448 3488 63040 3516
rect 62448 3476 62454 3488
rect 63034 3476 63040 3488
rect 63092 3476 63098 3528
rect 63586 3476 63592 3528
rect 63644 3516 63650 3528
rect 64230 3516 64236 3528
rect 63644 3488 64236 3516
rect 63644 3476 63650 3488
rect 64230 3476 64236 3488
rect 64288 3476 64294 3528
rect 68278 3476 68284 3528
rect 68336 3516 68342 3528
rect 68830 3516 68836 3528
rect 68336 3488 68836 3516
rect 68336 3476 68342 3488
rect 68830 3476 68836 3488
rect 68888 3476 68894 3528
rect 71866 3476 71872 3528
rect 71924 3516 71930 3528
rect 72878 3516 72884 3528
rect 71924 3488 72884 3516
rect 71924 3476 71930 3488
rect 72878 3476 72884 3488
rect 72936 3476 72942 3528
rect 515582 3516 515588 3528
rect 72988 3488 515588 3516
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 13078 3448 13084 3460
rect 2924 3420 13084 3448
rect 2924 3408 2930 3420
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 58802 3408 58808 3460
rect 58860 3448 58866 3460
rect 59262 3448 59268 3460
rect 58860 3420 59268 3448
rect 58860 3408 58866 3420
rect 59262 3408 59268 3420
rect 59320 3408 59326 3460
rect 72786 3408 72792 3460
rect 72844 3448 72850 3460
rect 72988 3448 73016 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 518158 3476 518164 3528
rect 518216 3516 518222 3528
rect 542906 3516 542912 3528
rect 518216 3488 542912 3516
rect 518216 3476 518222 3488
rect 542906 3476 542912 3488
rect 542964 3476 542970 3528
rect 554774 3476 554780 3528
rect 554832 3516 554838 3528
rect 555970 3516 555976 3528
rect 554832 3488 555976 3516
rect 554832 3476 554838 3488
rect 555970 3476 555976 3488
rect 556028 3476 556034 3528
rect 574756 3516 574784 3544
rect 580994 3516 581000 3528
rect 574756 3488 581000 3516
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 72844 3420 73016 3448
rect 73065 3451 73123 3457
rect 72844 3408 72850 3420
rect 73065 3417 73077 3451
rect 73111 3448 73123 3451
rect 522666 3448 522672 3460
rect 73111 3420 522672 3448
rect 73111 3417 73123 3420
rect 73065 3411 73123 3417
rect 522666 3408 522672 3420
rect 522724 3408 522730 3460
rect 528554 3408 528560 3460
rect 528612 3448 528618 3460
rect 529842 3448 529848 3460
rect 528612 3420 529848 3448
rect 528612 3408 528618 3420
rect 529842 3408 529848 3420
rect 529900 3408 529906 3460
rect 573358 3408 573364 3460
rect 573416 3448 573422 3460
rect 579798 3448 579804 3460
rect 573416 3420 579804 3448
rect 573416 3408 573422 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 76650 3340 76656 3392
rect 76708 3380 76714 3392
rect 77202 3380 77208 3392
rect 76708 3352 77208 3380
rect 76708 3340 76714 3352
rect 77202 3340 77208 3352
rect 77260 3340 77266 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 78306 3380 78312 3392
rect 77904 3352 78312 3380
rect 77904 3340 77910 3352
rect 78306 3340 78312 3352
rect 78364 3340 78370 3392
rect 81894 3340 81900 3392
rect 81952 3380 81958 3392
rect 82630 3380 82636 3392
rect 81952 3352 82636 3380
rect 81952 3340 81958 3352
rect 82630 3340 82636 3352
rect 82688 3340 82694 3392
rect 87322 3340 87328 3392
rect 87380 3380 87386 3392
rect 88242 3380 88248 3392
rect 87380 3352 88248 3380
rect 87380 3340 87386 3352
rect 88242 3340 88248 3352
rect 88300 3340 88306 3392
rect 89714 3340 89720 3392
rect 89772 3380 89778 3392
rect 90910 3380 90916 3392
rect 89772 3352 90916 3380
rect 89772 3340 89778 3352
rect 90910 3340 90916 3352
rect 90968 3340 90974 3392
rect 93302 3340 93308 3392
rect 93360 3380 93366 3392
rect 93762 3380 93768 3392
rect 93360 3352 93768 3380
rect 93360 3340 93366 3352
rect 93762 3340 93768 3352
rect 93820 3340 93826 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 94498 3380 94504 3392
rect 94004 3352 94504 3380
rect 94004 3340 94010 3352
rect 94498 3340 94504 3352
rect 94556 3340 94562 3392
rect 95694 3340 95700 3392
rect 95752 3380 95758 3392
rect 96522 3380 96528 3392
rect 95752 3352 96528 3380
rect 95752 3340 95758 3352
rect 96522 3340 96528 3352
rect 96580 3340 96586 3392
rect 96890 3340 96896 3392
rect 96948 3380 96954 3392
rect 97902 3380 97908 3392
rect 96948 3352 97908 3380
rect 96948 3340 96954 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 98086 3340 98092 3392
rect 98144 3380 98150 3392
rect 99374 3380 99380 3392
rect 98144 3352 99380 3380
rect 98144 3340 98150 3352
rect 99374 3340 99380 3352
rect 99432 3340 99438 3392
rect 101582 3340 101588 3392
rect 101640 3380 101646 3392
rect 102042 3380 102048 3392
rect 101640 3352 102048 3380
rect 101640 3340 101646 3352
rect 102042 3340 102048 3352
rect 102100 3340 102106 3392
rect 102778 3340 102784 3392
rect 102836 3380 102842 3392
rect 103422 3380 103428 3392
rect 102836 3352 103428 3380
rect 102836 3340 102842 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 105170 3340 105176 3392
rect 105228 3380 105234 3392
rect 106182 3380 106188 3392
rect 105228 3352 106188 3380
rect 105228 3340 105234 3352
rect 106182 3340 106188 3352
rect 106240 3340 106246 3392
rect 106366 3340 106372 3392
rect 106424 3380 106430 3392
rect 107654 3380 107660 3392
rect 106424 3352 107660 3380
rect 106424 3340 106430 3352
rect 107654 3340 107660 3352
rect 107712 3340 107718 3392
rect 114738 3340 114744 3392
rect 114796 3380 114802 3392
rect 115750 3380 115756 3392
rect 114796 3352 115756 3380
rect 114796 3340 114802 3352
rect 115750 3340 115756 3352
rect 115808 3340 115814 3392
rect 117314 3340 117320 3392
rect 117372 3380 117378 3392
rect 118234 3380 118240 3392
rect 117372 3352 118240 3380
rect 117372 3340 117378 3352
rect 118234 3340 118240 3352
rect 118292 3340 118298 3392
rect 119430 3340 119436 3392
rect 119488 3380 119494 3392
rect 119982 3380 119988 3392
rect 119488 3352 119988 3380
rect 119488 3340 119494 3352
rect 119982 3340 119988 3352
rect 120040 3340 120046 3392
rect 124214 3340 124220 3392
rect 124272 3380 124278 3392
rect 125502 3380 125508 3392
rect 124272 3352 125508 3380
rect 124272 3340 124278 3352
rect 125502 3340 125508 3352
rect 125560 3340 125566 3392
rect 127802 3340 127808 3392
rect 127860 3380 127866 3392
rect 128262 3380 128268 3392
rect 127860 3352 128268 3380
rect 127860 3340 127866 3352
rect 128262 3340 128268 3352
rect 128320 3340 128326 3392
rect 129734 3340 129740 3392
rect 129792 3380 129798 3392
rect 130194 3380 130200 3392
rect 129792 3352 130200 3380
rect 129792 3340 129798 3352
rect 130194 3340 130200 3352
rect 130252 3340 130258 3392
rect 136082 3340 136088 3392
rect 136140 3380 136146 3392
rect 136542 3380 136548 3392
rect 136140 3352 136548 3380
rect 136140 3340 136146 3352
rect 136542 3340 136548 3352
rect 136600 3340 136606 3392
rect 148042 3340 148048 3392
rect 148100 3380 148106 3392
rect 148962 3380 148968 3392
rect 148100 3352 148968 3380
rect 148100 3340 148106 3352
rect 148962 3340 148968 3352
rect 149020 3340 149026 3392
rect 157337 3383 157395 3389
rect 157337 3349 157349 3383
rect 157383 3380 157395 3383
rect 158714 3380 158720 3392
rect 157383 3352 158720 3380
rect 157383 3349 157395 3352
rect 157337 3343 157395 3349
rect 158714 3340 158720 3352
rect 158772 3340 158778 3392
rect 187786 3340 187792 3392
rect 187844 3380 187850 3392
rect 188430 3380 188436 3392
rect 187844 3352 188436 3380
rect 187844 3340 187850 3352
rect 188430 3340 188436 3352
rect 188488 3340 188494 3392
rect 189626 3340 189632 3392
rect 189684 3380 189690 3392
rect 190362 3380 190368 3392
rect 189684 3352 190368 3380
rect 189684 3340 189690 3352
rect 190362 3340 190368 3352
rect 190420 3340 190426 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 193122 3380 193128 3392
rect 192076 3352 193128 3380
rect 192076 3340 192082 3352
rect 193122 3340 193128 3352
rect 193180 3340 193186 3392
rect 226518 3340 226524 3392
rect 226576 3380 226582 3392
rect 227622 3380 227628 3392
rect 226576 3352 227628 3380
rect 226576 3340 226582 3352
rect 227622 3340 227628 3352
rect 227680 3340 227686 3392
rect 232498 3340 232504 3392
rect 232556 3380 232562 3392
rect 233142 3380 233148 3392
rect 232556 3352 233148 3380
rect 232556 3340 232562 3352
rect 233142 3340 233148 3352
rect 233200 3340 233206 3392
rect 239582 3340 239588 3392
rect 239640 3380 239646 3392
rect 240042 3380 240048 3392
rect 239640 3352 240048 3380
rect 239640 3340 239646 3352
rect 240042 3340 240048 3352
rect 240100 3340 240106 3392
rect 240778 3340 240784 3392
rect 240836 3380 240842 3392
rect 241422 3380 241428 3392
rect 240836 3352 241428 3380
rect 240836 3340 240842 3352
rect 241422 3340 241428 3352
rect 241480 3340 241486 3392
rect 249150 3340 249156 3392
rect 249208 3380 249214 3392
rect 249702 3380 249708 3392
rect 249208 3352 249708 3380
rect 249208 3340 249214 3352
rect 249702 3340 249708 3352
rect 249760 3340 249766 3392
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 251082 3380 251088 3392
rect 250404 3352 251088 3380
rect 250404 3340 250410 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 251450 3340 251456 3392
rect 251508 3380 251514 3392
rect 253937 3383 253995 3389
rect 253937 3380 253949 3383
rect 251508 3352 253949 3380
rect 251508 3340 251514 3352
rect 253937 3349 253949 3352
rect 253983 3349 253995 3383
rect 253937 3343 253995 3349
rect 262214 3340 262220 3392
rect 262272 3380 262278 3392
rect 263410 3380 263416 3392
rect 262272 3352 263416 3380
rect 262272 3340 262278 3352
rect 263410 3340 263416 3352
rect 263468 3340 263474 3392
rect 283650 3340 283656 3392
rect 283708 3380 283714 3392
rect 284202 3380 284208 3392
rect 283708 3352 284208 3380
rect 283708 3340 283714 3352
rect 284202 3340 284208 3352
rect 284260 3340 284266 3392
rect 285950 3340 285956 3392
rect 286008 3380 286014 3392
rect 286962 3380 286968 3392
rect 286008 3352 286968 3380
rect 286008 3340 286014 3352
rect 286962 3340 286968 3352
rect 287020 3340 287026 3392
rect 287054 3340 287060 3392
rect 287112 3380 287118 3392
rect 288342 3380 288348 3392
rect 287112 3352 288348 3380
rect 287112 3340 287118 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 293126 3340 293132 3392
rect 293184 3380 293190 3392
rect 293862 3380 293868 3392
rect 293184 3352 293868 3380
rect 293184 3340 293190 3352
rect 293862 3340 293868 3352
rect 293920 3340 293926 3392
rect 296714 3340 296720 3392
rect 296772 3380 296778 3392
rect 298002 3380 298008 3392
rect 296772 3352 298008 3380
rect 296772 3340 296778 3352
rect 298002 3340 298008 3352
rect 298060 3340 298066 3392
rect 301406 3340 301412 3392
rect 301464 3380 301470 3392
rect 302142 3380 302148 3392
rect 301464 3352 302148 3380
rect 301464 3340 301470 3352
rect 302142 3340 302148 3352
rect 302200 3340 302206 3392
rect 303798 3340 303804 3392
rect 303856 3380 303862 3392
rect 304902 3380 304908 3392
rect 303856 3352 304908 3380
rect 303856 3340 303862 3352
rect 304902 3340 304908 3352
rect 304960 3340 304966 3392
rect 304994 3340 305000 3392
rect 305052 3380 305058 3392
rect 306190 3380 306196 3392
rect 305052 3352 306196 3380
rect 305052 3340 305058 3352
rect 306190 3340 306196 3352
rect 306248 3340 306254 3392
rect 326430 3340 326436 3392
rect 326488 3380 326494 3392
rect 326982 3380 326988 3392
rect 326488 3352 326988 3380
rect 326488 3340 326494 3352
rect 326982 3340 326988 3352
rect 327040 3340 327046 3392
rect 330018 3340 330024 3392
rect 330076 3380 330082 3392
rect 331122 3380 331128 3392
rect 330076 3352 331128 3380
rect 330076 3340 330082 3352
rect 331122 3340 331128 3352
rect 331180 3340 331186 3392
rect 344278 3340 344284 3392
rect 344336 3380 344342 3392
rect 344922 3380 344928 3392
rect 344336 3352 344928 3380
rect 344336 3340 344342 3352
rect 344922 3340 344928 3352
rect 344980 3340 344986 3392
rect 361574 3340 361580 3392
rect 361632 3380 361638 3392
rect 362126 3380 362132 3392
rect 361632 3352 362132 3380
rect 361632 3340 361638 3352
rect 362126 3340 362132 3352
rect 362184 3340 362190 3392
rect 363322 3340 363328 3392
rect 363380 3380 363386 3392
rect 364150 3380 364156 3392
rect 363380 3352 364156 3380
rect 363380 3340 363386 3352
rect 364150 3340 364156 3352
rect 364208 3340 364214 3392
rect 364518 3340 364524 3392
rect 364576 3380 364582 3392
rect 365622 3380 365628 3392
rect 364576 3352 365628 3380
rect 364576 3340 364582 3352
rect 365622 3340 365628 3352
rect 365680 3340 365686 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 366910 3380 366916 3392
rect 365772 3352 366916 3380
rect 365772 3340 365778 3352
rect 366910 3340 366916 3352
rect 366968 3340 366974 3392
rect 370406 3340 370412 3392
rect 370464 3380 370470 3392
rect 371142 3380 371148 3392
rect 370464 3352 371148 3380
rect 370464 3340 370470 3352
rect 371142 3340 371148 3352
rect 371200 3340 371206 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375190 3380 375196 3392
rect 374052 3352 375196 3380
rect 374052 3340 374058 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 379974 3340 379980 3392
rect 380032 3380 380038 3392
rect 380802 3380 380808 3392
rect 380032 3352 380808 3380
rect 380032 3340 380038 3352
rect 380802 3340 380808 3352
rect 380860 3340 380866 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 385862 3340 385868 3392
rect 385920 3380 385926 3392
rect 386322 3380 386328 3392
rect 385920 3352 386328 3380
rect 385920 3340 385926 3352
rect 386322 3340 386328 3352
rect 386380 3340 386386 3392
rect 388254 3340 388260 3392
rect 388312 3380 388318 3392
rect 389082 3380 389088 3392
rect 388312 3352 389088 3380
rect 388312 3340 388318 3352
rect 389082 3340 389088 3352
rect 389140 3340 389146 3392
rect 421558 3340 421564 3392
rect 421616 3380 421622 3392
rect 422202 3380 422208 3392
rect 421616 3352 422208 3380
rect 421616 3340 421622 3352
rect 422202 3340 422208 3352
rect 422260 3340 422266 3392
rect 425054 3340 425060 3392
rect 425112 3380 425118 3392
rect 426342 3380 426348 3392
rect 425112 3352 426348 3380
rect 425112 3340 425118 3352
rect 426342 3340 426348 3352
rect 426400 3340 426406 3392
rect 433334 3340 433340 3392
rect 433392 3380 433398 3392
rect 434622 3380 434628 3392
rect 433392 3352 434628 3380
rect 433392 3340 433398 3352
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 439406 3340 439412 3392
rect 439464 3380 439470 3392
rect 440142 3380 440148 3392
rect 439464 3352 440148 3380
rect 439464 3340 439470 3352
rect 440142 3340 440148 3352
rect 440200 3340 440206 3392
rect 459554 3340 459560 3392
rect 459612 3380 459618 3392
rect 460842 3380 460848 3392
rect 459612 3352 460848 3380
rect 459612 3340 459618 3352
rect 460842 3340 460848 3352
rect 460900 3340 460906 3392
rect 483474 3340 483480 3392
rect 483532 3380 483538 3392
rect 484302 3380 484308 3392
rect 483532 3352 484308 3380
rect 483532 3340 483538 3352
rect 484302 3340 484308 3352
rect 484360 3340 484366 3392
rect 496449 3383 496507 3389
rect 496449 3349 496461 3383
rect 496495 3380 496507 3383
rect 507854 3380 507860 3392
rect 496495 3352 507860 3380
rect 496495 3349 496507 3352
rect 496449 3343 496507 3349
rect 507854 3340 507860 3352
rect 507912 3340 507918 3392
rect 113177 3315 113235 3321
rect 113177 3281 113189 3315
rect 113223 3312 113235 3315
rect 122745 3315 122803 3321
rect 122745 3312 122757 3315
rect 113223 3284 122757 3312
rect 113223 3281 113235 3284
rect 113177 3275 113235 3281
rect 122745 3281 122757 3284
rect 122791 3281 122803 3315
rect 122745 3275 122803 3281
rect 132497 3315 132555 3321
rect 132497 3281 132509 3315
rect 132543 3312 132555 3315
rect 146941 3315 146999 3321
rect 146941 3312 146953 3315
rect 132543 3284 146953 3312
rect 132543 3281 132555 3284
rect 132497 3275 132555 3281
rect 146941 3281 146953 3284
rect 146987 3281 146999 3315
rect 146941 3275 146999 3281
rect 155126 3272 155132 3324
rect 155184 3312 155190 3324
rect 155862 3312 155868 3324
rect 155184 3284 155868 3312
rect 155184 3272 155190 3284
rect 155862 3272 155868 3284
rect 155920 3272 155926 3324
rect 175366 3272 175372 3324
rect 175424 3312 175430 3324
rect 176562 3312 176568 3324
rect 175424 3284 176568 3312
rect 175424 3272 175430 3284
rect 176562 3272 176568 3284
rect 176620 3272 176626 3324
rect 182542 3272 182548 3324
rect 182600 3312 182606 3324
rect 183462 3312 183468 3324
rect 182600 3284 183468 3312
rect 182600 3272 182606 3284
rect 183462 3272 183468 3284
rect 183520 3272 183526 3324
rect 241974 3272 241980 3324
rect 242032 3312 242038 3324
rect 242802 3312 242808 3324
rect 242032 3284 242808 3312
rect 242032 3272 242038 3284
rect 242802 3272 242808 3284
rect 242860 3272 242866 3324
rect 339494 3272 339500 3324
rect 339552 3312 339558 3324
rect 340782 3312 340788 3324
rect 339552 3284 340788 3312
rect 339552 3272 339558 3284
rect 340782 3272 340788 3284
rect 340840 3272 340846 3324
rect 494146 3272 494152 3324
rect 494204 3312 494210 3324
rect 503717 3315 503775 3321
rect 503717 3312 503729 3315
rect 494204 3284 503729 3312
rect 494204 3272 494210 3284
rect 503717 3281 503729 3284
rect 503763 3281 503775 3315
rect 503717 3275 503775 3281
rect 542998 3272 543004 3324
rect 543056 3312 543062 3324
rect 546494 3312 546500 3324
rect 543056 3284 546500 3312
rect 543056 3272 543062 3284
rect 546494 3272 546500 3284
rect 546552 3272 546558 3324
rect 89990 3204 89996 3256
rect 90048 3244 90054 3256
rect 90910 3244 90916 3256
rect 90048 3216 90916 3244
rect 90048 3204 90054 3216
rect 90910 3204 90916 3216
rect 90968 3204 90974 3256
rect 93857 3247 93915 3253
rect 93857 3213 93869 3247
rect 93903 3244 93915 3247
rect 103425 3247 103483 3253
rect 103425 3244 103437 3247
rect 93903 3216 103437 3244
rect 93903 3213 93915 3216
rect 93857 3207 93915 3213
rect 103425 3213 103437 3216
rect 103471 3213 103483 3247
rect 103425 3207 103483 3213
rect 218146 3204 218152 3256
rect 218204 3244 218210 3256
rect 219250 3244 219256 3256
rect 218204 3216 219256 3244
rect 218204 3204 218210 3216
rect 219250 3204 219256 3216
rect 219308 3204 219314 3256
rect 277670 3204 277676 3256
rect 277728 3244 277734 3256
rect 278682 3244 278688 3256
rect 277728 3216 278688 3244
rect 277728 3204 277734 3216
rect 278682 3204 278688 3216
rect 278740 3204 278746 3256
rect 304994 3204 305000 3256
rect 305052 3244 305058 3256
rect 306282 3244 306288 3256
rect 305052 3216 306288 3244
rect 305052 3204 305058 3216
rect 306282 3204 306288 3216
rect 306340 3204 306346 3256
rect 365714 3204 365720 3256
rect 365772 3244 365778 3256
rect 367002 3244 367008 3256
rect 365772 3216 367008 3244
rect 365772 3204 365778 3216
rect 367002 3204 367008 3216
rect 367060 3204 367066 3256
rect 200390 3136 200396 3188
rect 200448 3176 200454 3188
rect 201402 3176 201408 3188
rect 200448 3148 201408 3176
rect 200448 3136 200454 3148
rect 201402 3136 201408 3148
rect 201460 3136 201466 3188
rect 215846 3136 215852 3188
rect 215904 3176 215910 3188
rect 216582 3176 216588 3188
rect 215904 3148 216588 3176
rect 215904 3136 215910 3148
rect 216582 3136 216588 3148
rect 216640 3136 216646 3188
rect 328822 3136 328828 3188
rect 328880 3176 328886 3188
rect 329742 3176 329748 3188
rect 328880 3148 329748 3176
rect 328880 3136 328886 3148
rect 329742 3136 329748 3148
rect 329800 3136 329806 3188
rect 353754 3136 353760 3188
rect 353812 3176 353818 3188
rect 354582 3176 354588 3188
rect 353812 3148 354588 3176
rect 353812 3136 353818 3148
rect 354582 3136 354588 3148
rect 354640 3136 354646 3188
rect 354950 3136 354956 3188
rect 355008 3176 355014 3188
rect 355962 3176 355968 3188
rect 355008 3148 355968 3176
rect 355008 3136 355014 3148
rect 355962 3136 355968 3148
rect 356020 3136 356026 3188
rect 172974 3068 172980 3120
rect 173032 3108 173038 3120
rect 173802 3108 173808 3120
rect 173032 3080 173808 3108
rect 173032 3068 173038 3080
rect 173802 3068 173808 3080
rect 173860 3068 173866 3120
rect 415670 3068 415676 3120
rect 415728 3108 415734 3120
rect 416682 3108 416688 3120
rect 415728 3080 416688 3108
rect 415728 3068 415734 3080
rect 416682 3068 416688 3080
rect 416740 3068 416746 3120
rect 84930 3000 84936 3052
rect 84988 3040 84994 3052
rect 85482 3040 85488 3052
rect 84988 3012 85488 3040
rect 84988 3000 84994 3012
rect 85482 3000 85488 3012
rect 85540 3000 85546 3052
rect 163498 3000 163504 3052
rect 163556 3040 163562 3052
rect 164142 3040 164148 3052
rect 163556 3012 164148 3040
rect 163556 3000 163562 3012
rect 164142 3000 164148 3012
rect 164200 3000 164206 3052
rect 164694 3000 164700 3052
rect 164752 3040 164758 3052
rect 165522 3040 165528 3052
rect 164752 3012 165528 3040
rect 164752 3000 164758 3012
rect 165522 3000 165528 3012
rect 165580 3000 165586 3052
rect 319254 3000 319260 3052
rect 319312 3040 319318 3052
rect 319990 3040 319996 3052
rect 319312 3012 319996 3040
rect 319312 3000 319318 3012
rect 319990 3000 319996 3012
rect 320048 3000 320054 3052
rect 347866 3000 347872 3052
rect 347924 3040 347930 3052
rect 349062 3040 349068 3052
rect 347924 3012 349068 3040
rect 347924 3000 347930 3012
rect 349062 3000 349068 3012
rect 349120 3000 349126 3052
rect 504358 3000 504364 3052
rect 504416 3040 504422 3052
rect 507210 3040 507216 3052
rect 504416 3012 507216 3040
rect 504416 3000 504422 3012
rect 507210 3000 507216 3012
rect 507268 3000 507274 3052
rect 181346 2932 181352 2984
rect 181404 2972 181410 2984
rect 182082 2972 182088 2984
rect 181404 2944 182088 2972
rect 181404 2932 181410 2944
rect 182082 2932 182088 2944
rect 182140 2932 182146 2984
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 8938 2904 8944 2916
rect 4120 2876 8944 2904
rect 4120 2864 4126 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 50522 2864 50528 2916
rect 50580 2904 50586 2916
rect 50982 2904 50988 2916
rect 50580 2876 50988 2904
rect 50580 2864 50586 2876
rect 50982 2864 50988 2876
rect 51040 2864 51046 2916
rect 69474 2864 69480 2916
rect 69532 2904 69538 2916
rect 70118 2904 70124 2916
rect 69532 2876 70124 2904
rect 69532 2864 69538 2876
rect 70118 2864 70124 2876
rect 70176 2864 70182 2916
rect 139670 2864 139676 2916
rect 139728 2904 139734 2916
rect 140682 2904 140688 2916
rect 139728 2876 140688 2904
rect 139728 2864 139734 2876
rect 140682 2864 140688 2876
rect 140740 2864 140746 2916
rect 144730 2836 144736 2848
rect 144472 2808 144736 2836
rect 144472 2780 144500 2808
rect 144730 2796 144736 2808
rect 144788 2796 144794 2848
rect 161106 2796 161112 2848
rect 161164 2836 161170 2848
rect 161382 2836 161388 2848
rect 161164 2808 161388 2836
rect 161164 2796 161170 2808
rect 161382 2796 161388 2808
rect 161440 2796 161446 2848
rect 203889 2839 203947 2845
rect 203889 2805 203901 2839
rect 203935 2836 203947 2839
rect 204070 2836 204076 2848
rect 203935 2808 204076 2836
rect 203935 2805 203947 2808
rect 203889 2799 203947 2805
rect 204070 2796 204076 2808
rect 204128 2796 204134 2848
rect 212442 2836 212448 2848
rect 212276 2808 212448 2836
rect 212276 2780 212304 2808
rect 212442 2796 212448 2808
rect 212500 2796 212506 2848
rect 333882 2836 333888 2848
rect 333624 2808 333888 2836
rect 333624 2780 333652 2808
rect 333882 2796 333888 2808
rect 333940 2796 333946 2848
rect 393041 2839 393099 2845
rect 393041 2805 393053 2839
rect 393087 2836 393099 2839
rect 393222 2836 393228 2848
rect 393087 2808 393228 2836
rect 393087 2805 393099 2808
rect 393041 2799 393099 2805
rect 393222 2796 393228 2808
rect 393280 2796 393286 2848
rect 453666 2796 453672 2848
rect 453724 2836 453730 2848
rect 453942 2836 453948 2848
rect 453724 2808 453948 2836
rect 453724 2796 453730 2808
rect 453942 2796 453948 2808
rect 454000 2796 454006 2848
rect 144454 2728 144460 2780
rect 144512 2728 144518 2780
rect 212258 2728 212264 2780
rect 212316 2728 212322 2780
rect 333606 2728 333612 2780
rect 333664 2728 333670 2780
rect 511994 2728 512000 2780
rect 512052 2768 512058 2780
rect 512546 2768 512552 2780
rect 512052 2740 512552 2768
rect 512052 2728 512058 2740
rect 512546 2728 512552 2740
rect 512604 2728 512610 2780
rect 536834 2320 536840 2372
rect 536892 2360 536898 2372
rect 538122 2360 538128 2372
rect 536892 2332 538128 2360
rect 536892 2320 536898 2332
rect 538122 2320 538128 2332
rect 538180 2320 538186 2372
rect 445754 2184 445760 2236
rect 445812 2224 445818 2236
rect 446582 2224 446588 2236
rect 445812 2196 446588 2224
rect 445812 2184 445818 2196
rect 446582 2184 446588 2196
rect 446640 2184 446646 2236
rect 99466 552 99472 604
rect 99524 592 99530 604
rect 100478 592 100484 604
rect 99524 564 100484 592
rect 99524 552 99530 564
rect 100478 552 100484 564
rect 100536 552 100542 604
rect 120074 552 120080 604
rect 120132 592 120138 604
rect 120626 592 120632 604
rect 120132 564 120632 592
rect 120132 552 120138 564
rect 120626 552 120632 564
rect 120684 552 120690 604
rect 128354 552 128360 604
rect 128412 592 128418 604
rect 128998 592 129004 604
rect 128412 564 129004 592
rect 128412 552 128418 564
rect 128998 552 129004 564
rect 129056 552 129062 604
rect 171134 552 171140 604
rect 171192 592 171198 604
rect 171778 592 171784 604
rect 171192 564 171784 592
rect 171192 552 171198 564
rect 171778 552 171784 564
rect 171836 552 171842 604
rect 186314 552 186320 604
rect 186372 592 186378 604
rect 187234 592 187240 604
rect 186372 564 187240 592
rect 186372 552 186378 564
rect 187234 552 187240 564
rect 187292 552 187298 604
rect 195974 552 195980 604
rect 196032 592 196038 604
rect 196802 592 196808 604
rect 196032 564 196808 592
rect 196032 552 196038 564
rect 196802 552 196808 564
rect 196860 552 196866 604
rect 203886 592 203892 604
rect 203847 564 203892 592
rect 203886 552 203892 564
rect 203944 552 203950 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 223574 552 223580 604
rect 223632 592 223638 604
rect 224126 592 224132 604
rect 223632 564 224132 592
rect 223632 552 223638 564
rect 224126 552 224132 564
rect 224184 552 224190 604
rect 247954 552 247960 604
rect 248012 592 248018 604
rect 248322 592 248328 604
rect 248012 564 248328 592
rect 248012 552 248018 564
rect 248322 552 248328 564
rect 248380 552 248386 604
rect 358814 552 358820 604
rect 358872 592 358878 604
rect 359734 592 359740 604
rect 358872 564 359740 592
rect 358872 552 358878 564
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 393038 592 393044 604
rect 392999 564 393044 592
rect 393038 552 393044 564
rect 393096 552 393102 604
rect 393314 552 393320 604
rect 393372 592 393378 604
rect 394234 592 394240 604
rect 393372 564 394240 592
rect 393372 552 393378 564
rect 394234 552 394240 564
rect 394292 552 394298 604
rect 396074 552 396080 604
rect 396132 592 396138 604
rect 396626 592 396632 604
rect 396132 564 396632 592
rect 396132 552 396138 564
rect 396626 552 396632 564
rect 396684 552 396690 604
rect 401594 552 401600 604
rect 401652 592 401658 604
rect 402514 592 402520 604
rect 401652 564 402520 592
rect 401652 552 401658 564
rect 402514 552 402520 564
rect 402572 552 402578 604
rect 410886 592 410892 604
rect 410847 564 410892 592
rect 410886 552 410892 564
rect 410944 552 410950 604
rect 492674 552 492680 604
rect 492732 592 492738 604
rect 492950 592 492956 604
rect 492732 564 492956 592
rect 492732 552 492738 564
rect 492950 552 492956 564
rect 493008 552 493014 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 500954 552 500960 604
rect 501012 592 501018 604
rect 501230 592 501236 604
rect 501012 564 501236 592
rect 501012 552 501018 564
rect 501230 552 501236 564
rect 501288 552 501294 604
rect 502426 592 502432 604
rect 502387 564 502432 592
rect 502426 552 502432 564
rect 502484 552 502490 604
rect 505094 552 505100 604
rect 505152 592 505158 604
rect 506014 592 506020 604
rect 505152 564 506020 592
rect 505152 552 505158 564
rect 506014 552 506020 564
rect 506072 552 506078 604
rect 508130 552 508136 604
rect 508188 592 508194 604
rect 508406 592 508412 604
rect 508188 564 508412 592
rect 508188 552 508194 564
rect 508406 552 508412 564
rect 508464 552 508470 604
rect 513650 552 513656 604
rect 513708 592 513714 604
rect 514386 592 514392 604
rect 513708 564 514392 592
rect 513708 552 513714 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 576854 552 576860 604
rect 576912 592 576918 604
rect 577406 592 577412 604
rect 576912 564 577412 592
rect 576912 552 576918 564
rect 577406 552 577412 564
rect 577464 552 577470 604
rect 581086 552 581092 604
rect 581144 592 581150 604
rect 582190 592 582196 604
rect 581144 564 582196 592
rect 581144 552 581150 564
rect 582190 552 582196 564
rect 582248 552 582254 604
<< via1 >>
rect 137836 700680 137888 700732
rect 138664 700680 138716 700732
rect 70308 700612 70360 700664
rect 154120 700612 154172 700664
rect 81348 700544 81400 700596
rect 218980 700544 219032 700596
rect 75828 700476 75880 700528
rect 235172 700476 235224 700528
rect 283840 700476 283892 700528
rect 298744 700476 298796 700528
rect 332508 700476 332560 700528
rect 520464 700476 520516 700528
rect 77208 700408 77260 700460
rect 348792 700408 348844 700460
rect 364984 700408 365036 700460
rect 509976 700408 510028 700460
rect 67456 700340 67508 700392
rect 413652 700340 413704 700392
rect 68744 700272 68796 700324
rect 462320 700272 462372 700324
rect 529204 700272 529256 700324
rect 543464 700272 543516 700324
rect 543556 700272 543608 700324
rect 559656 700272 559708 700324
rect 8116 700204 8168 700256
rect 14464 700204 14516 700256
rect 397460 699932 397512 699984
rect 398748 699932 398800 699984
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 40500 699660 40552 699712
rect 43444 699660 43496 699712
rect 88340 699660 88392 699712
rect 89168 699660 89220 699712
rect 104900 699660 104952 699712
rect 105452 699660 105504 699712
rect 543004 699660 543056 699712
rect 543556 699660 543608 699712
rect 259368 698912 259420 698964
rect 300124 698912 300176 698964
rect 202788 697552 202840 697604
rect 502340 697552 502392 697604
rect 169944 695444 169996 695496
rect 170312 695444 170364 695496
rect 72700 694084 72752 694136
rect 429200 692792 429252 692844
rect 429936 692792 429988 692844
rect 477500 692792 477552 692844
rect 478604 692792 478656 692844
rect 169944 687896 169996 687948
rect 170128 687896 170180 687948
rect 522304 685856 522356 685908
rect 580172 685856 580224 685908
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 169760 683068 169812 683120
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 173900 673956 173952 674008
rect 178316 673956 178368 674008
rect 154580 673752 154632 673804
rect 162216 673752 162268 673804
rect 477500 673480 477552 673532
rect 477684 673480 477736 673532
rect 429200 673412 429252 673464
rect 429476 673412 429528 673464
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 3424 667904 3476 667956
rect 502432 667904 502484 667956
rect 170220 666544 170272 666596
rect 72884 659608 72936 659660
rect 73068 659608 73120 659660
rect 73068 656820 73120 656872
rect 477500 654100 477552 654152
rect 477684 654100 477736 654152
rect 3056 652740 3108 652792
rect 17224 652740 17276 652792
rect 177948 650020 178000 650072
rect 580172 650020 580224 650072
rect 72976 647275 73028 647284
rect 72976 647241 72985 647275
rect 72985 647241 73019 647275
rect 73019 647241 73028 647275
rect 72976 647232 73028 647241
rect 169944 647232 169996 647284
rect 170036 647232 170088 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 72976 640364 73028 640416
rect 169944 640364 169996 640416
rect 170036 640364 170088 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 72792 640228 72844 640280
rect 515404 638936 515456 638988
rect 580172 638936 580224 638988
rect 72792 637551 72844 637560
rect 72792 637517 72801 637551
rect 72801 637517 72835 637551
rect 72835 637517 72844 637551
rect 72792 637508 72844 637517
rect 477500 634788 477552 634840
rect 477684 634788 477736 634840
rect 169852 630640 169904 630692
rect 170036 630640 170088 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 398748 628532 398800 628584
rect 501604 628532 501656 628584
rect 73068 627920 73120 627972
rect 81716 626560 81768 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 55864 623772 55916 623824
rect 72976 618264 73028 618316
rect 73068 618264 73120 618316
rect 72976 618171 73028 618180
rect 72976 618137 72985 618171
rect 72985 618137 73019 618171
rect 73019 618137 73028 618171
rect 72976 618128 73028 618137
rect 79876 617516 79928 617568
rect 477684 617516 477736 617568
rect 43444 616088 43496 616140
rect 398840 616088 398892 616140
rect 138664 614728 138716 614780
rect 382280 614728 382332 614780
rect 169760 611328 169812 611380
rect 170036 611328 170088 611380
rect 429200 611328 429252 611380
rect 429476 611328 429528 611380
rect 128360 610580 128412 610632
rect 543004 610580 543056 610632
rect 3424 609968 3476 610020
rect 48964 609968 49016 610020
rect 73068 608676 73120 608728
rect 380440 608676 380492 608728
rect 521844 608676 521896 608728
rect 57888 608608 57940 608660
rect 313648 608608 313700 608660
rect 375472 608608 375524 608660
rect 520372 608608 520424 608660
rect 501788 608540 501840 608592
rect 501972 608540 502024 608592
rect 81624 607860 81676 607912
rect 169760 607860 169812 607912
rect 298744 607860 298796 607912
rect 338304 607860 338356 607912
rect 67548 607316 67600 607368
rect 155592 607316 155644 607368
rect 372896 607316 372948 607368
rect 521660 607316 521712 607368
rect 64788 607248 64840 607300
rect 180248 607248 180300 607300
rect 353208 607248 353260 607300
rect 504824 607248 504876 607300
rect 81256 607180 81308 607232
rect 204904 607180 204956 607232
rect 340880 607180 340932 607232
rect 505744 607180 505796 607232
rect 69756 606568 69808 606620
rect 461952 606568 462004 606620
rect 66168 606500 66220 606552
rect 190184 606500 190236 606552
rect 61844 606432 61896 606484
rect 224776 606432 224828 606484
rect 328552 606432 328604 606484
rect 429200 606432 429252 606484
rect 61752 606364 61804 606416
rect 244464 606364 244516 606416
rect 81164 606296 81216 606348
rect 318616 606296 318668 606348
rect 471704 606296 471756 606348
rect 514944 606296 514996 606348
rect 74264 606228 74316 606280
rect 323584 606228 323636 606280
rect 390192 606228 390244 606280
rect 520556 606228 520608 606280
rect 71596 606160 71648 606212
rect 199936 606160 199988 606212
rect 209872 606160 209924 606212
rect 554044 606160 554096 606212
rect 82084 606092 82136 606144
rect 165344 606092 165396 606144
rect 508504 606092 508556 606144
rect 167920 606024 167972 606076
rect 456984 606024 457036 606076
rect 517796 606024 517848 606076
rect 168288 605956 168340 606008
rect 573364 605956 573416 606008
rect 86408 605888 86460 605940
rect 523040 605888 523092 605940
rect 39396 605820 39448 605872
rect 503904 605820 503956 605872
rect 72424 605276 72476 605328
rect 246856 605276 246908 605328
rect 72976 605208 73028 605260
rect 192576 605208 192628 605260
rect 82268 605140 82320 605192
rect 360568 605140 360620 605192
rect 83280 605072 83332 605124
rect 145656 605072 145708 605124
rect 79324 605004 79376 605056
rect 160376 605004 160428 605056
rect 444656 605004 444708 605056
rect 521752 605004 521804 605056
rect 67272 604936 67324 604988
rect 222200 604936 222252 604988
rect 419816 604936 419868 604988
rect 513564 604936 513616 604988
rect 57244 604868 57296 604920
rect 276664 604868 276716 604920
rect 412456 604868 412508 604920
rect 513380 604868 513432 604920
rect 21364 604800 21416 604852
rect 256792 604800 256844 604852
rect 387800 604800 387852 604852
rect 516416 604800 516468 604852
rect 79968 604732 80020 604784
rect 325976 604732 326028 604784
rect 333336 604732 333388 604784
rect 502984 604732 503036 604784
rect 68928 604664 68980 604716
rect 101128 604664 101180 604716
rect 358176 604664 358228 604716
rect 503812 604664 503864 604716
rect 242072 604596 242124 604648
rect 554780 604596 554832 604648
rect 68284 604528 68336 604580
rect 153016 604528 153068 604580
rect 172888 604528 172940 604580
rect 514116 604528 514168 604580
rect 140688 604460 140740 604512
rect 503720 604460 503772 604512
rect 289820 604052 289872 604104
rect 299388 604052 299440 604104
rect 328460 604052 328512 604104
rect 338028 604052 338080 604104
rect 347780 604052 347832 604104
rect 357348 604052 357400 604104
rect 345848 603916 345900 603968
rect 492680 603916 492732 603968
rect 64604 603848 64656 603900
rect 98736 603848 98788 603900
rect 363144 603848 363196 603900
rect 481732 603848 481784 603900
rect 483020 603848 483072 603900
rect 492772 603848 492824 603900
rect 81440 603780 81492 603832
rect 410064 603780 410116 603832
rect 452016 603780 452068 603832
rect 502064 603780 502116 603832
rect 71044 603712 71096 603764
rect 96160 603712 96212 603764
rect 190092 603712 190144 603764
rect 417424 603712 417476 603764
rect 444472 603712 444524 603764
rect 449164 603712 449216 603764
rect 454408 603712 454460 603764
rect 513472 603712 513524 603764
rect 516876 603712 516928 603764
rect 525708 603712 525760 603764
rect 79416 603644 79468 603696
rect 108488 603644 108540 603696
rect 148048 603644 148100 603696
rect 309232 603644 309284 603696
rect 318708 603644 318760 603696
rect 469312 603644 469364 603696
rect 479248 603644 479300 603696
rect 502248 603644 502300 603696
rect 533988 603644 534040 603696
rect 540888 603644 540940 603696
rect 71688 603576 71740 603628
rect 125784 603576 125836 603628
rect 422392 603576 422444 603628
rect 56508 603508 56560 603560
rect 111064 603508 111116 603560
rect 321008 603508 321060 603560
rect 381452 603508 381504 603560
rect 432328 603508 432380 603560
rect 515496 603508 515548 603560
rect 97908 603440 97960 603492
rect 197544 603440 197596 603492
rect 351828 603440 351880 603492
rect 466920 603440 466972 603492
rect 484216 603440 484268 603492
rect 517612 603440 517664 603492
rect 67180 603372 67232 603424
rect 202512 603372 202564 603424
rect 481640 603372 481692 603424
rect 531964 603372 532016 603424
rect 64144 603304 64196 603356
rect 150624 603304 150676 603356
rect 175280 603304 175332 603356
rect 318800 603304 318852 603356
rect 493968 603304 494020 603356
rect 516324 603304 516376 603356
rect 83188 603236 83240 603288
rect 261760 603236 261812 603288
rect 343272 603236 343324 603288
rect 512092 603236 512144 603288
rect 28264 603168 28316 603220
rect 303712 603168 303764 603220
rect 311256 603168 311308 603220
rect 552664 603168 552716 603220
rect 60556 603100 60608 603152
rect 88800 603100 88852 603152
rect 301320 603100 301372 603152
rect 346400 603100 346452 603152
rect 395160 603100 395212 603152
rect 407488 603100 407540 603152
rect 507216 603100 507268 603152
rect 88340 603032 88392 603084
rect 351828 603032 351880 603084
rect 492680 602760 492732 602812
rect 498200 602760 498252 602812
rect 31668 602624 31720 602676
rect 239496 602624 239548 602676
rect 70216 602556 70268 602608
rect 232136 602556 232188 602608
rect 8944 602488 8996 602540
rect 133328 602488 133380 602540
rect 59268 602420 59320 602472
rect 68836 602420 68888 602472
rect 88248 602420 88300 602472
rect 481732 602420 481784 602472
rect 517704 602420 517756 602472
rect 71504 602352 71556 602404
rect 104808 602352 104860 602404
rect 381452 602352 381504 602404
rect 580264 602352 580316 602404
rect 104900 602284 104952 602336
rect 464344 602284 464396 602336
rect 82176 602216 82228 602268
rect 143080 602216 143132 602268
rect 474280 602216 474332 602268
rect 507860 602216 507912 602268
rect 74448 602148 74500 602200
rect 135720 602148 135772 602200
rect 377864 602148 377916 602200
rect 524420 602148 524472 602200
rect 9036 602080 9088 602132
rect 121000 602080 121052 602132
rect 370504 602080 370556 602132
rect 569960 602080 570012 602132
rect 83464 602012 83516 602064
rect 226892 602012 226944 602064
rect 269488 602012 269540 602064
rect 481824 602012 481876 602064
rect 27528 601944 27580 601996
rect 263876 601944 263928 601996
rect 309048 601944 309100 601996
rect 543004 601944 543056 601996
rect 237288 601876 237340 601928
rect 514760 601876 514812 601928
rect 229928 601808 229980 601860
rect 510620 601808 510672 601860
rect 72516 601740 72568 601792
rect 115940 601740 115992 601792
rect 459560 601740 459612 601792
rect 118608 601672 118660 601724
rect 507124 601672 507176 601724
rect 92388 601604 92440 601656
rect 504824 601332 504876 601384
rect 507308 601332 507360 601384
rect 91100 601307 91152 601316
rect 91100 601273 91109 601307
rect 91109 601273 91143 601307
rect 91143 601273 91152 601307
rect 91100 601264 91152 601273
rect 97908 601307 97960 601316
rect 97908 601273 97917 601307
rect 97917 601273 97951 601307
rect 97951 601273 97960 601307
rect 97908 601264 97960 601273
rect 105820 601307 105872 601316
rect 105820 601273 105829 601307
rect 105829 601273 105863 601307
rect 105863 601273 105872 601307
rect 105820 601264 105872 601273
rect 113180 601307 113232 601316
rect 113180 601273 113189 601307
rect 113189 601273 113223 601307
rect 113223 601273 113232 601307
rect 113180 601264 113232 601273
rect 123116 601307 123168 601316
rect 123116 601273 123125 601307
rect 123125 601273 123159 601307
rect 123159 601273 123168 601307
rect 123116 601264 123168 601273
rect 131028 601307 131080 601316
rect 131028 601273 131037 601307
rect 131037 601273 131071 601307
rect 131071 601273 131080 601307
rect 131028 601264 131080 601273
rect 183008 601307 183060 601316
rect 183008 601273 183017 601307
rect 183017 601273 183051 601307
rect 183051 601273 183060 601307
rect 183008 601264 183060 601273
rect 187332 601307 187384 601316
rect 187332 601273 187341 601307
rect 187341 601273 187375 601307
rect 187375 601273 187384 601307
rect 187332 601264 187384 601273
rect 215024 601307 215076 601316
rect 215024 601273 215033 601307
rect 215033 601273 215067 601307
rect 215067 601273 215076 601307
rect 215024 601264 215076 601273
rect 217600 601307 217652 601316
rect 217600 601273 217609 601307
rect 217609 601273 217643 601307
rect 217643 601273 217652 601307
rect 217600 601264 217652 601273
rect 234252 601264 234304 601316
rect 254216 601264 254268 601316
rect 271420 601307 271472 601316
rect 271420 601273 271429 601307
rect 271429 601273 271463 601307
rect 271463 601273 271472 601307
rect 271420 601264 271472 601273
rect 274456 601307 274508 601316
rect 274456 601273 274465 601307
rect 274465 601273 274499 601307
rect 274499 601273 274508 601307
rect 274456 601264 274508 601273
rect 283748 601307 283800 601316
rect 283748 601273 283757 601307
rect 283757 601273 283791 601307
rect 283791 601273 283800 601307
rect 283748 601264 283800 601273
rect 291200 601264 291252 601316
rect 347964 601307 348016 601316
rect 347964 601273 347973 601307
rect 347973 601273 348007 601307
rect 348007 601273 348016 601307
rect 347964 601264 348016 601273
rect 355876 601264 355928 601316
rect 365720 601307 365772 601316
rect 365720 601273 365729 601307
rect 365729 601273 365763 601307
rect 365763 601273 365772 601307
rect 365720 601264 365772 601273
rect 425152 601307 425204 601316
rect 425152 601273 425161 601307
rect 425161 601273 425195 601307
rect 425195 601273 425204 601307
rect 425152 601264 425204 601273
rect 437296 601307 437348 601316
rect 437296 601273 437305 601307
rect 437305 601273 437339 601307
rect 437339 601273 437348 601307
rect 437296 601264 437348 601273
rect 498200 601264 498252 601316
rect 503996 601264 504048 601316
rect 83464 601060 83516 601112
rect 83648 601060 83700 601112
rect 75552 600992 75604 601044
rect 81072 600924 81124 600976
rect 74356 600856 74408 600908
rect 71136 600788 71188 600840
rect 72884 600720 72936 600772
rect 543740 600924 543792 600976
rect 509332 600788 509384 600840
rect 511356 600720 511408 600772
rect 76564 600652 76616 600704
rect 516232 600652 516284 600704
rect 69664 600584 69716 600636
rect 556160 600584 556212 600636
rect 62028 600516 62080 600568
rect 518164 600516 518216 600568
rect 83648 600448 83700 600500
rect 532700 600448 532752 600500
rect 61936 600380 61988 600432
rect 518900 600380 518952 600432
rect 15844 600312 15896 600364
rect 509884 600312 509936 600364
rect 501512 600244 501564 600296
rect 83464 599972 83516 600024
rect 75644 599768 75696 599820
rect 501696 599632 501748 599684
rect 514024 599632 514076 599684
rect 580356 599564 580408 599616
rect 2688 599224 2740 599276
rect 64696 598952 64748 599004
rect 78680 598952 78732 599004
rect 503996 598272 504048 598324
rect 523132 598272 523184 598324
rect 502064 598204 502116 598256
rect 534080 598204 534132 598256
rect 30288 596776 30340 596828
rect 81440 596776 81492 596828
rect 502248 596776 502300 596828
rect 512828 596776 512880 596828
rect 504364 596207 504416 596216
rect 504364 596173 504373 596207
rect 504373 596173 504407 596207
rect 504407 596173 504416 596207
rect 504364 596164 504416 596173
rect 2872 594804 2924 594856
rect 32404 594804 32456 594856
rect 20076 594056 20128 594108
rect 78680 594056 78732 594108
rect 42708 592628 42760 592680
rect 82912 592628 82964 592680
rect 60464 592016 60516 592068
rect 78680 592016 78732 592068
rect 511264 592016 511316 592068
rect 579896 592016 579948 592068
rect 507308 587120 507360 587172
rect 523224 587120 523276 587172
rect 503904 586508 503956 586560
rect 540244 586508 540296 586560
rect 72792 586440 72844 586492
rect 73068 586440 73120 586492
rect 503904 582360 503956 582412
rect 574100 582360 574152 582412
rect 560944 579640 560996 579692
rect 580172 579640 580224 579692
rect 504364 578212 504416 578264
rect 504456 578212 504508 578264
rect 75736 577124 75788 577176
rect 78956 577124 79008 577176
rect 72792 576852 72844 576904
rect 73068 576852 73120 576904
rect 501696 574064 501748 574116
rect 501972 574064 502024 574116
rect 76932 572704 76984 572756
rect 78772 572704 78824 572756
rect 504364 572772 504416 572824
rect 504272 572636 504324 572688
rect 503904 571344 503956 571396
rect 538864 571344 538916 571396
rect 50344 569916 50396 569968
rect 78680 569916 78732 569968
rect 3424 567196 3476 567248
rect 25504 567196 25556 567248
rect 503904 567196 503956 567248
rect 517980 567196 518032 567248
rect 46848 565836 46900 565888
rect 78680 565836 78732 565888
rect 503904 564408 503956 564460
rect 514852 564408 514904 564460
rect 504364 562912 504416 562964
rect 504548 562912 504600 562964
rect 67364 561688 67416 561740
rect 78680 561688 78732 561740
rect 503904 560260 503956 560312
rect 520648 560260 520700 560312
rect 77024 558900 77076 558952
rect 79600 558900 79652 558952
rect 512828 558900 512880 558952
rect 513012 558900 513064 558952
rect 569316 556180 569368 556232
rect 580172 556180 580224 556232
rect 501512 556112 501564 556164
rect 501512 555976 501564 556028
rect 501696 554820 501748 554872
rect 63408 554752 63460 554804
rect 78680 554752 78732 554804
rect 501604 554752 501656 554804
rect 503904 554684 503956 554736
rect 529204 554684 529256 554736
rect 3148 552032 3200 552084
rect 39304 552032 39356 552084
rect 503904 549244 503956 549296
rect 518992 549244 519044 549296
rect 72792 547816 72844 547868
rect 73068 547816 73120 547868
rect 504456 547136 504508 547188
rect 536840 547136 536892 547188
rect 503904 545164 503956 545216
rect 515036 545164 515088 545216
rect 512644 545096 512696 545148
rect 579896 545096 579948 545148
rect 503904 541628 503956 541680
rect 565084 541628 565136 541680
rect 3424 538228 3476 538280
rect 43444 538228 43496 538280
rect 72792 538228 72844 538280
rect 73068 538228 73120 538280
rect 503904 538228 503956 538280
rect 521936 538228 521988 538280
rect 501604 536800 501656 536852
rect 501696 536664 501748 536716
rect 504456 534148 504508 534200
rect 507216 534012 507268 534064
rect 580172 534012 580224 534064
rect 504364 531335 504416 531344
rect 504364 531301 504373 531335
rect 504373 531301 504407 531335
rect 504407 531301 504416 531335
rect 504364 531292 504416 531301
rect 512828 531292 512880 531344
rect 513012 531292 513064 531344
rect 504456 531267 504508 531276
rect 504456 531233 504465 531267
rect 504465 531233 504499 531267
rect 504499 531233 504508 531267
rect 504456 531224 504508 531233
rect 512828 529864 512880 529916
rect 513012 529864 513064 529916
rect 76840 525784 76892 525836
rect 78680 525784 78732 525836
rect 503904 524424 503956 524476
rect 506480 524424 506532 524476
rect 504456 524331 504508 524340
rect 504456 524297 504465 524331
rect 504465 524297 504499 524331
rect 504499 524297 504508 524331
rect 504456 524288 504508 524297
rect 503904 520276 503956 520328
rect 520740 520276 520792 520328
rect 501696 520208 501748 520260
rect 75460 518916 75512 518968
rect 78864 518916 78916 518968
rect 504364 514811 504416 514820
rect 504364 514777 504373 514811
rect 504373 514777 504407 514811
rect 504407 514777 504416 514811
rect 504364 514768 504416 514777
rect 504364 512023 504416 512032
rect 504364 511989 504373 512023
rect 504373 511989 504407 512023
rect 504407 511989 504416 512023
rect 504364 511980 504416 511989
rect 512828 511980 512880 512032
rect 513012 511980 513064 512032
rect 63316 510620 63368 510672
rect 78680 510620 78732 510672
rect 501604 510663 501656 510672
rect 501604 510629 501613 510663
rect 501613 510629 501647 510663
rect 501647 510629 501656 510663
rect 501604 510620 501656 510629
rect 512828 510552 512880 510604
rect 513012 510552 513064 510604
rect 565084 510552 565136 510604
rect 580172 510552 580224 510604
rect 3148 509260 3200 509312
rect 9128 509260 9180 509312
rect 64512 507832 64564 507884
rect 78680 507832 78732 507884
rect 82912 507875 82964 507884
rect 82912 507841 82921 507875
rect 82921 507841 82955 507875
rect 82955 507841 82964 507875
rect 82912 507832 82964 507841
rect 501604 507807 501656 507816
rect 501604 507773 501613 507807
rect 501613 507773 501647 507807
rect 501647 507773 501656 507807
rect 501604 507764 501656 507773
rect 504364 505112 504416 505164
rect 504456 504976 504508 505028
rect 66076 503684 66128 503736
rect 78680 503684 78732 503736
rect 82912 501712 82964 501764
rect 82912 501619 82964 501628
rect 82912 501585 82921 501619
rect 82921 501585 82955 501619
rect 82955 501585 82964 501619
rect 82912 501576 82964 501585
rect 77116 500012 77168 500064
rect 79048 500012 79100 500064
rect 508504 499468 508556 499520
rect 580172 499468 580224 499520
rect 501696 498176 501748 498228
rect 503904 498176 503956 498228
rect 507952 498176 508004 498228
rect 504180 497496 504232 497548
rect 504364 497496 504416 497548
rect 61660 496816 61712 496868
rect 78680 496816 78732 496868
rect 3424 496748 3476 496800
rect 503904 494028 503956 494080
rect 513656 494028 513708 494080
rect 512828 491283 512880 491292
rect 512828 491249 512837 491283
rect 512837 491249 512871 491283
rect 512871 491249 512880 491283
rect 512828 491240 512880 491249
rect 72792 489812 72844 489864
rect 73068 489812 73120 489864
rect 503904 487160 503956 487212
rect 571984 487160 572036 487212
rect 65984 485800 66036 485852
rect 78680 485800 78732 485852
rect 504364 485800 504416 485852
rect 567844 485800 567896 485852
rect 580172 485800 580224 485852
rect 504456 485664 504508 485716
rect 503904 483012 503956 483064
rect 522028 483012 522080 483064
rect 504456 482944 504508 482996
rect 504640 482944 504692 482996
rect 512828 481695 512880 481704
rect 512828 481661 512837 481695
rect 512837 481661 512871 481695
rect 512871 481661 512880 481695
rect 512828 481652 512880 481661
rect 3792 481584 3844 481636
rect 39396 481584 39448 481636
rect 72792 480224 72844 480276
rect 73068 480224 73120 480276
rect 501604 480224 501656 480276
rect 501696 480224 501748 480276
rect 61568 478864 61620 478916
rect 78680 478864 78732 478916
rect 503904 476076 503956 476128
rect 516508 476076 516560 476128
rect 83004 474920 83056 474972
rect 503904 473356 503956 473408
rect 523316 473356 523368 473408
rect 48964 471928 49016 471980
rect 78680 471928 78732 471980
rect 512828 471971 512880 471980
rect 512828 471937 512837 471971
rect 512837 471937 512871 471971
rect 512871 471937 512880 471971
rect 512828 471928 512880 471937
rect 83004 469208 83056 469260
rect 503904 469208 503956 469260
rect 510804 469208 510856 469260
rect 501604 467780 501656 467832
rect 501696 467780 501748 467832
rect 504364 466420 504416 466472
rect 504456 466352 504508 466404
rect 504180 463632 504232 463684
rect 504456 463632 504508 463684
rect 512828 462383 512880 462392
rect 512828 462349 512837 462383
rect 512837 462349 512871 462383
rect 512871 462349 512880 462383
rect 512828 462340 512880 462349
rect 565084 462340 565136 462392
rect 580172 462340 580224 462392
rect 503904 461524 503956 461576
rect 508044 461524 508096 461576
rect 68652 459552 68704 459604
rect 78680 459552 78732 459604
rect 75368 456764 75420 456816
rect 78680 456764 78732 456816
rect 509884 452548 509936 452600
rect 580172 452548 580224 452600
rect 512828 452523 512880 452532
rect 512828 452489 512837 452523
rect 512837 452489 512871 452523
rect 512871 452489 512880 452523
rect 512828 452480 512880 452489
rect 72792 451188 72844 451240
rect 73068 451188 73120 451240
rect 501604 449896 501656 449948
rect 501696 449896 501748 449948
rect 74080 448536 74132 448588
rect 78680 448536 78732 448588
rect 82912 448579 82964 448588
rect 82912 448545 82921 448579
rect 82921 448545 82955 448579
rect 82955 448545 82964 448579
rect 82912 448536 82964 448545
rect 501604 448468 501656 448520
rect 501696 448468 501748 448520
rect 503904 447108 503956 447160
rect 506572 447108 506624 447160
rect 60372 445748 60424 445800
rect 78680 445748 78732 445800
rect 82912 444320 82964 444372
rect 504456 444320 504508 444372
rect 503904 442960 503956 443012
rect 509608 442960 509660 443012
rect 512828 443003 512880 443012
rect 512828 442969 512837 443003
rect 512837 442969 512871 443003
rect 512871 442969 512880 443003
rect 512828 442960 512880 442969
rect 82912 441940 82964 441992
rect 72792 441668 72844 441720
rect 73068 441668 73120 441720
rect 82912 441711 82964 441720
rect 82912 441677 82921 441711
rect 82921 441677 82955 441711
rect 82955 441677 82964 441711
rect 82912 441668 82964 441677
rect 64420 441600 64472 441652
rect 78680 441600 78732 441652
rect 503904 440240 503956 440292
rect 509516 440240 509568 440292
rect 82820 440172 82872 440224
rect 82912 440172 82964 440224
rect 514116 440172 514168 440224
rect 579620 440172 579672 440224
rect 503904 436092 503956 436144
rect 519084 436092 519136 436144
rect 504364 434775 504416 434784
rect 504364 434741 504373 434775
rect 504373 434741 504407 434775
rect 504407 434741 504416 434775
rect 504364 434732 504416 434741
rect 512828 433279 512880 433288
rect 512828 433245 512837 433279
rect 512837 433245 512871 433279
rect 512871 433245 512880 433279
rect 512828 433236 512880 433245
rect 503904 432488 503956 432540
rect 506756 432488 506808 432540
rect 72792 431876 72844 431928
rect 73068 431876 73120 431928
rect 59084 430584 59136 430636
rect 78680 430584 78732 430636
rect 82820 430516 82872 430568
rect 83004 430516 83056 430568
rect 503904 429156 503956 429208
rect 522120 429156 522172 429208
rect 19984 427796 20036 427848
rect 78680 427796 78732 427848
rect 504364 427796 504416 427848
rect 504456 427728 504508 427780
rect 503904 425076 503956 425128
rect 509424 425076 509476 425128
rect 3240 425008 3292 425060
rect 69756 425008 69808 425060
rect 504456 425008 504508 425060
rect 501972 423648 502024 423700
rect 502064 423648 502116 423700
rect 512828 423691 512880 423700
rect 512828 423657 512837 423691
rect 512837 423657 512871 423691
rect 512871 423657 512880 423691
rect 512828 423648 512880 423657
rect 72792 422288 72844 422340
rect 73068 422288 73120 422340
rect 503904 420928 503956 420980
rect 506664 420928 506716 420980
rect 46204 419500 46256 419552
rect 78680 419500 78732 419552
rect 3424 417392 3476 417444
rect 69756 417392 69808 417444
rect 76748 416780 76800 416832
rect 78680 416780 78732 416832
rect 504364 415463 504416 415472
rect 504364 415429 504373 415463
rect 504373 415429 504407 415463
rect 504407 415429 504416 415463
rect 504364 415420 504416 415429
rect 512828 413967 512880 413976
rect 512828 413933 512837 413967
rect 512837 413933 512871 413967
rect 512871 413933 512880 413967
rect 512828 413924 512880 413933
rect 65892 412632 65944 412684
rect 78680 412632 78732 412684
rect 72792 412564 72844 412616
rect 73068 412564 73120 412616
rect 501604 411272 501656 411324
rect 501788 411272 501840 411324
rect 504364 408484 504416 408536
rect 504456 408348 504508 408400
rect 503904 407124 503956 407176
rect 508228 407124 508280 407176
rect 63224 405696 63276 405748
rect 78680 405696 78732 405748
rect 512828 404379 512880 404388
rect 512828 404345 512837 404379
rect 512837 404345 512871 404379
rect 512871 404345 512880 404379
rect 512828 404336 512880 404345
rect 516784 404336 516836 404388
rect 580172 404336 580224 404388
rect 72792 402976 72844 403028
rect 73068 402976 73120 403028
rect 503904 402976 503956 403028
rect 513748 402976 513800 403028
rect 64328 401616 64380 401668
rect 78680 401616 78732 401668
rect 504456 400868 504508 400920
rect 504640 400868 504692 400920
rect 503904 398828 503956 398880
rect 520832 398828 520884 398880
rect 33784 397468 33836 397520
rect 78680 397468 78732 397520
rect 3332 394680 3384 394732
rect 69848 394680 69900 394732
rect 512828 394655 512880 394664
rect 512828 394621 512837 394655
rect 512837 394621 512871 394655
rect 512871 394621 512880 394655
rect 512828 394612 512880 394621
rect 72792 393252 72844 393304
rect 73068 393252 73120 393304
rect 504364 393252 504416 393304
rect 504456 393252 504508 393304
rect 507124 393252 507176 393304
rect 580172 393252 580224 393304
rect 501696 391892 501748 391944
rect 501788 391892 501840 391944
rect 503904 389172 503956 389224
rect 573456 389172 573508 389224
rect 63132 386384 63184 386436
rect 78680 386384 78732 386436
rect 82912 386248 82964 386300
rect 512828 385135 512880 385144
rect 512828 385101 512837 385135
rect 512837 385101 512871 385135
rect 512871 385101 512880 385135
rect 512828 385092 512880 385101
rect 503904 385024 503956 385076
rect 549904 385024 549956 385076
rect 72792 383732 72844 383784
rect 73068 383732 73120 383784
rect 65800 383664 65852 383716
rect 78680 383664 78732 383716
rect 502984 382916 503036 382968
rect 523408 382916 523460 382968
rect 503904 380876 503956 380928
rect 519176 380876 519228 380928
rect 3424 379516 3476 379568
rect 13176 379516 13228 379568
rect 503904 378156 503956 378208
rect 506940 378156 506992 378208
rect 501696 376660 501748 376712
rect 501788 376660 501840 376712
rect 503904 375300 503956 375352
rect 522304 375300 522356 375352
rect 512828 375275 512880 375284
rect 512828 375241 512837 375275
rect 512837 375241 512871 375275
rect 512871 375241 512880 375275
rect 512828 375232 512880 375241
rect 82820 374799 82872 374808
rect 82820 374765 82829 374799
rect 82829 374765 82863 374799
rect 82863 374765 82872 374799
rect 82820 374756 82872 374765
rect 72792 373940 72844 373992
rect 73068 373940 73120 373992
rect 49608 368500 49660 368552
rect 78680 368500 78732 368552
rect 514116 368500 514168 368552
rect 580172 368500 580224 368552
rect 503996 367072 504048 367124
rect 506848 367072 506900 367124
rect 504456 367004 504508 367056
rect 504364 366936 504416 366988
rect 512828 365755 512880 365764
rect 512828 365721 512837 365755
rect 512837 365721 512871 365755
rect 512871 365721 512880 365755
rect 512828 365712 512880 365721
rect 72792 364352 72844 364404
rect 73068 364352 73120 364404
rect 503996 362924 504048 362976
rect 516600 362924 516652 362976
rect 37924 361564 37976 361616
rect 78680 361564 78732 361616
rect 501696 358776 501748 358828
rect 501788 358776 501840 358828
rect 512828 357552 512880 357604
rect 75276 357416 75328 357468
rect 78680 357416 78732 357468
rect 512828 357416 512880 357468
rect 569224 357416 569276 357468
rect 580172 357416 580224 357468
rect 501604 357348 501656 357400
rect 501696 357348 501748 357400
rect 512828 356031 512880 356040
rect 512828 355997 512837 356031
rect 512837 355997 512871 356031
rect 512871 355997 512880 356031
rect 512828 355988 512880 355997
rect 505744 355308 505796 355360
rect 519636 355308 519688 355360
rect 13176 351840 13228 351892
rect 78680 351840 78732 351892
rect 15936 346400 15988 346452
rect 78680 346400 78732 346452
rect 512828 346443 512880 346452
rect 512828 346409 512837 346443
rect 512837 346409 512871 346443
rect 512871 346409 512880 346443
rect 512828 346400 512880 346409
rect 504088 345040 504140 345092
rect 513840 345040 513892 345092
rect 82912 342499 82964 342508
rect 82912 342465 82921 342499
rect 82921 342465 82955 342499
rect 82955 342465 82964 342499
rect 82912 342456 82964 342465
rect 504088 340892 504140 340944
rect 527824 340892 527876 340944
rect 501604 339396 501656 339448
rect 501696 339396 501748 339448
rect 504088 338104 504140 338156
rect 519268 338104 519320 338156
rect 82912 336855 82964 336864
rect 82912 336821 82921 336855
rect 82921 336821 82955 336855
rect 82955 336821 82964 336855
rect 82912 336812 82964 336821
rect 3424 336744 3476 336796
rect 72608 336744 72660 336796
rect 512828 336719 512880 336728
rect 512828 336685 512837 336719
rect 512837 336685 512871 336719
rect 512871 336685 512880 336719
rect 512828 336676 512880 336685
rect 57796 335316 57848 335368
rect 78680 335316 78732 335368
rect 504088 335248 504140 335300
rect 569316 335248 569368 335300
rect 63040 332596 63092 332648
rect 78680 332596 78732 332648
rect 17224 329740 17276 329792
rect 78680 329740 78732 329792
rect 512828 327131 512880 327140
rect 512828 327097 512837 327131
rect 512837 327097 512871 327131
rect 512871 327097 512880 327131
rect 512828 327088 512880 327097
rect 76656 324300 76708 324352
rect 78680 324300 78732 324352
rect 3240 324232 3292 324284
rect 76564 324232 76616 324284
rect 504088 322940 504140 322992
rect 512184 322940 512236 322992
rect 9128 322872 9180 322924
rect 78680 322872 78732 322924
rect 514024 322872 514076 322924
rect 580172 322872 580224 322924
rect 82820 318792 82872 318844
rect 82912 318792 82964 318844
rect 504088 318792 504140 318844
rect 515128 318792 515180 318844
rect 9128 317432 9180 317484
rect 78680 317432 78732 317484
rect 512828 317364 512880 317416
rect 512920 317364 512972 317416
rect 504088 316004 504140 316056
rect 558184 316004 558236 316056
rect 72792 315936 72844 315988
rect 73068 315936 73120 315988
rect 504364 314644 504416 314696
rect 504456 314644 504508 314696
rect 515496 311788 515548 311840
rect 580172 311788 580224 311840
rect 71320 310496 71372 310548
rect 78680 310496 78732 310548
rect 3424 308932 3476 308984
rect 9128 308932 9180 308984
rect 72792 306348 72844 306400
rect 73068 306348 73120 306400
rect 504088 306280 504140 306332
rect 567844 306280 567896 306332
rect 76564 299480 76616 299532
rect 79232 299480 79284 299532
rect 82912 299523 82964 299532
rect 82912 299489 82921 299523
rect 82921 299489 82955 299523
rect 82955 299489 82964 299523
rect 82912 299480 82964 299489
rect 540244 299412 540296 299464
rect 579804 299412 579856 299464
rect 512828 298052 512880 298104
rect 512920 298052 512972 298104
rect 72792 296624 72844 296676
rect 73068 296624 73120 296676
rect 70124 295332 70176 295384
rect 78680 295332 78732 295384
rect 3424 295264 3476 295316
rect 21364 295264 21416 295316
rect 82912 294720 82964 294772
rect 82912 294627 82964 294636
rect 82912 294593 82921 294627
rect 82921 294593 82955 294627
rect 82955 294593 82964 294627
rect 82912 294584 82964 294593
rect 82912 294244 82964 294296
rect 504088 293972 504140 294024
rect 512276 293972 512328 294024
rect 68560 292544 68612 292596
rect 78680 292544 78732 292596
rect 504088 289824 504140 289876
rect 508320 289824 508372 289876
rect 72792 287036 72844 287088
rect 73068 287036 73120 287088
rect 504088 285676 504140 285728
rect 540244 285676 540296 285728
rect 504088 282888 504140 282940
rect 545120 282888 545172 282940
rect 72792 281528 72844 281580
rect 78680 281528 78732 281580
rect 66996 277380 67048 277432
rect 78680 277380 78732 277432
rect 72700 277312 72752 277364
rect 73068 277312 73120 277364
rect 554044 275952 554096 276004
rect 580172 275952 580224 276004
rect 504088 274660 504140 274712
rect 519360 274660 519412 274712
rect 82912 273819 82964 273828
rect 82912 273785 82921 273819
rect 82921 273785 82955 273819
rect 82955 273785 82964 273819
rect 82912 273776 82964 273785
rect 70032 273232 70084 273284
rect 78680 273232 78732 273284
rect 512828 269084 512880 269136
rect 513012 269084 513064 269136
rect 72700 267724 72752 267776
rect 73068 267724 73120 267776
rect 504088 267724 504140 267776
rect 515312 267724 515364 267776
rect 57704 266364 57756 266416
rect 78680 266364 78732 266416
rect 3424 264936 3476 264988
rect 68376 264936 68428 264988
rect 55864 263508 55916 263560
rect 78680 263508 78732 263560
rect 504088 260856 504140 260908
rect 507124 260856 507176 260908
rect 82912 259471 82964 259480
rect 82912 259437 82921 259471
rect 82921 259437 82955 259471
rect 82955 259437 82964 259471
rect 82912 259428 82964 259437
rect 82820 259360 82872 259412
rect 82912 259156 82964 259208
rect 72700 258748 72752 258800
rect 73068 258748 73120 258800
rect 504088 256708 504140 256760
rect 508136 256708 508188 256760
rect 66904 251268 66956 251320
rect 78680 251268 78732 251320
rect 3424 251200 3476 251252
rect 68468 251200 68520 251252
rect 567844 251200 567896 251252
rect 580172 251200 580224 251252
rect 512828 249840 512880 249892
rect 513012 249840 513064 249892
rect 504088 249772 504140 249824
rect 518072 249772 518124 249824
rect 67088 249704 67140 249756
rect 78680 249704 78732 249756
rect 72700 249092 72752 249144
rect 73068 249092 73120 249144
rect 504088 245624 504140 245676
rect 547144 245624 547196 245676
rect 78312 245556 78364 245608
rect 79508 245556 79560 245608
rect 504088 242904 504140 242956
rect 507032 242904 507084 242956
rect 73988 241476 74040 241528
rect 78680 241476 78732 241528
rect 72700 239436 72752 239488
rect 73068 239436 73120 239488
rect 69940 237396 69992 237448
rect 78680 237396 78732 237448
rect 3424 237328 3476 237380
rect 69664 237328 69716 237380
rect 504088 234608 504140 234660
rect 516692 234608 516744 234660
rect 55864 233248 55916 233300
rect 78680 233248 78732 233300
rect 504088 231820 504140 231872
rect 519544 231820 519596 231872
rect 519636 231412 519688 231464
rect 520924 231412 520976 231464
rect 512828 230460 512880 230512
rect 513012 230460 513064 230512
rect 72700 229712 72752 229764
rect 73068 229712 73120 229764
rect 61476 229100 61528 229152
rect 78680 229100 78732 229152
rect 531964 229032 532016 229084
rect 580172 229032 580224 229084
rect 504088 227740 504140 227792
rect 510896 227740 510948 227792
rect 504088 223592 504140 223644
rect 512460 223592 512512 223644
rect 3148 223524 3200 223576
rect 72516 223524 72568 223576
rect 68744 223456 68796 223508
rect 78680 223456 78732 223508
rect 504088 220872 504140 220924
rect 509700 220872 509752 220924
rect 82912 219512 82964 219564
rect 82912 219011 82964 219020
rect 82912 218977 82921 219011
rect 82921 218977 82955 219011
rect 82955 218977 82964 219011
rect 82912 218968 82964 218977
rect 540244 217948 540296 218000
rect 580172 217948 580224 218000
rect 83004 217404 83056 217456
rect 72700 216928 72752 216980
rect 73068 216928 73120 216980
rect 504088 212508 504140 212560
rect 540244 212508 540296 212560
rect 72516 211148 72568 211200
rect 78680 211148 78732 211200
rect 82912 210672 82964 210724
rect 72700 210400 72752 210452
rect 73068 210400 73120 210452
rect 79508 210400 79560 210452
rect 79692 210400 79744 210452
rect 82912 209924 82964 209976
rect 82912 209788 82964 209840
rect 504088 209788 504140 209840
rect 512552 209788 512604 209840
rect 73896 208360 73948 208412
rect 78680 208360 78732 208412
rect 3424 208292 3476 208344
rect 57244 208292 57296 208344
rect 82912 207723 82964 207732
rect 82912 207689 82921 207723
rect 82921 207689 82955 207723
rect 82955 207689 82964 207723
rect 82912 207680 82964 207689
rect 82912 207476 82964 207528
rect 511448 204280 511500 204332
rect 580172 204280 580224 204332
rect 512828 201424 512880 201476
rect 513012 201424 513064 201476
rect 72332 200744 72384 200796
rect 73068 200744 73120 200796
rect 79508 199520 79560 199572
rect 79692 199520 79744 199572
rect 82912 195279 82964 195288
rect 82912 195245 82921 195279
rect 82921 195245 82955 195279
rect 82955 195245 82964 195279
rect 82912 195236 82964 195245
rect 504180 194556 504232 194608
rect 513932 194556 513984 194608
rect 3148 194488 3200 194540
rect 71136 194488 71188 194540
rect 504364 193808 504416 193860
rect 515220 193808 515272 193860
rect 72700 193196 72752 193248
rect 78680 193196 78732 193248
rect 68744 190476 68796 190528
rect 78680 190476 78732 190528
rect 79508 190476 79560 190528
rect 79692 190476 79744 190528
rect 504180 187688 504232 187740
rect 554044 187688 554096 187740
rect 82912 182928 82964 182980
rect 82912 182724 82964 182776
rect 71228 182180 71280 182232
rect 78680 182180 78732 182232
rect 512828 182112 512880 182164
rect 513012 182112 513064 182164
rect 3240 180752 3292 180804
rect 20076 180752 20128 180804
rect 72332 180752 72384 180804
rect 73068 180752 73120 180804
rect 79508 180752 79560 180804
rect 79692 180752 79744 180804
rect 81072 179324 81124 179376
rect 81900 179324 81952 179376
rect 75184 178100 75236 178152
rect 82268 178100 82320 178152
rect 65708 178032 65760 178084
rect 78680 178032 78732 178084
rect 79968 176672 80020 176724
rect 80704 176672 80756 176724
rect 82912 173476 82964 173528
rect 82912 173340 82964 173392
rect 82912 172252 82964 172304
rect 509240 171776 509292 171828
rect 527180 171776 527232 171828
rect 72332 171164 72384 171216
rect 73068 171164 73120 171216
rect 65616 171096 65668 171148
rect 78680 171096 78732 171148
rect 79508 171096 79560 171148
rect 79692 171096 79744 171148
rect 511356 171028 511408 171080
rect 580172 171028 580224 171080
rect 503720 170756 503772 170808
rect 509240 170756 509292 170808
rect 79508 166268 79560 166320
rect 79692 166268 79744 166320
rect 503720 165588 503772 165640
rect 512368 165588 512420 165640
rect 3516 165520 3568 165572
rect 72424 165520 72476 165572
rect 68468 165452 68520 165504
rect 78680 165452 78732 165504
rect 512828 162843 512880 162852
rect 512828 162809 512837 162843
rect 512837 162809 512871 162843
rect 512871 162809 512880 162843
rect 512828 162800 512880 162809
rect 72424 161372 72476 161424
rect 73068 161372 73120 161424
rect 14464 158652 14516 158704
rect 78680 158652 78732 158704
rect 82820 158652 82872 158704
rect 573456 158652 573508 158704
rect 579804 158652 579856 158704
rect 82912 158380 82964 158432
rect 82912 158015 82964 158024
rect 82912 157981 82921 158015
rect 82921 157981 82955 158015
rect 82955 157981 82964 158015
rect 82912 157972 82964 157981
rect 82820 157836 82872 157888
rect 82728 157403 82780 157412
rect 82728 157369 82737 157403
rect 82737 157369 82771 157403
rect 82771 157369 82780 157403
rect 82728 157360 82780 157369
rect 69664 155184 69716 155236
rect 82176 155184 82228 155236
rect 68468 153212 68520 153264
rect 78680 153212 78732 153264
rect 512828 153255 512880 153264
rect 512828 153221 512837 153255
rect 512837 153221 512871 153255
rect 512871 153221 512880 153255
rect 512828 153212 512880 153221
rect 72424 151784 72476 151836
rect 73068 151784 73120 151836
rect 79508 151784 79560 151836
rect 79692 151784 79744 151836
rect 503720 151784 503772 151836
rect 552756 151784 552808 151836
rect 3148 151716 3200 151768
rect 68284 151716 68336 151768
rect 14464 149064 14516 149116
rect 78680 149064 78732 149116
rect 82912 148248 82964 148300
rect 17224 146276 17276 146328
rect 78680 146276 78732 146328
rect 82912 145188 82964 145240
rect 82912 144984 82964 145036
rect 82820 144848 82872 144900
rect 82912 144823 82964 144832
rect 82912 144789 82921 144823
rect 82921 144789 82955 144823
rect 82955 144789 82964 144823
rect 82912 144780 82964 144789
rect 82912 143692 82964 143744
rect 82912 143556 82964 143608
rect 504548 143556 504600 143608
rect 510988 143556 511040 143608
rect 512828 143531 512880 143540
rect 512828 143497 512837 143531
rect 512837 143497 512871 143531
rect 512871 143497 512880 143531
rect 512828 143488 512880 143497
rect 72424 142060 72476 142112
rect 73068 142060 73120 142112
rect 79692 142060 79744 142112
rect 79968 142060 80020 142112
rect 504548 140768 504600 140820
rect 508412 140768 508464 140820
rect 82820 140267 82872 140276
rect 82820 140233 82829 140267
rect 82829 140233 82863 140267
rect 82863 140233 82872 140267
rect 82820 140224 82872 140233
rect 71136 140020 71188 140072
rect 82912 140020 82964 140072
rect 82820 137207 82872 137216
rect 82820 137173 82829 137207
rect 82829 137173 82863 137207
rect 82863 137173 82872 137207
rect 82820 137164 82872 137173
rect 3516 135804 3568 135856
rect 9128 135804 9180 135856
rect 552664 135192 552716 135244
rect 580172 135192 580224 135244
rect 82636 134716 82688 134768
rect 82912 134716 82964 134768
rect 512828 133943 512880 133952
rect 512828 133909 512837 133943
rect 512837 133909 512871 133943
rect 512871 133909 512880 133943
rect 512828 133900 512880 133909
rect 503076 133016 503128 133068
rect 508504 133016 508556 133068
rect 82912 132608 82964 132660
rect 72424 132472 72476 132524
rect 73068 132472 73120 132524
rect 79692 132472 79744 132524
rect 79968 132472 80020 132524
rect 82544 132472 82596 132524
rect 57244 131112 57296 131164
rect 78680 131112 78732 131164
rect 72424 126964 72476 127016
rect 78680 126964 78732 127016
rect 73804 126216 73856 126268
rect 79324 126216 79376 126268
rect 504548 125604 504600 125656
rect 509792 125604 509844 125656
rect 82912 124176 82964 124228
rect 512828 124151 512880 124160
rect 512828 124117 512837 124151
rect 512837 124117 512871 124151
rect 512871 124117 512880 124151
rect 512828 124108 512880 124117
rect 538864 124108 538916 124160
rect 580172 124108 580224 124160
rect 82912 124083 82964 124092
rect 82912 124049 82921 124083
rect 82921 124049 82955 124083
rect 82955 124049 82964 124083
rect 82912 124040 82964 124049
rect 72332 122748 72384 122800
rect 73068 122748 73120 122800
rect 79692 122748 79744 122800
rect 79968 122748 80020 122800
rect 3424 121456 3476 121508
rect 11704 121456 11756 121508
rect 81072 120028 81124 120080
rect 81900 120028 81952 120080
rect 82912 118711 82964 118720
rect 82912 118677 82921 118711
rect 82921 118677 82955 118711
rect 82955 118677 82964 118711
rect 82912 118668 82964 118677
rect 82912 115243 82964 115252
rect 82912 115209 82921 115243
rect 82921 115209 82955 115243
rect 82955 115209 82964 115243
rect 82912 115200 82964 115209
rect 512828 114563 512880 114572
rect 512828 114529 512837 114563
rect 512837 114529 512871 114563
rect 512871 114529 512880 114563
rect 512828 114520 512880 114529
rect 72332 113160 72384 113212
rect 73068 113160 73120 113212
rect 79692 113160 79744 113212
rect 79968 113160 80020 113212
rect 82912 110984 82964 111036
rect 503260 110440 503312 110492
rect 509240 110440 509292 110492
rect 73068 110372 73120 110424
rect 78680 110372 78732 110424
rect 73068 109012 73120 109064
rect 73804 109012 73856 109064
rect 73804 107856 73856 107908
rect 74172 107856 74224 107908
rect 4068 107652 4120 107704
rect 74264 107652 74316 107704
rect 503352 107652 503404 107704
rect 531964 107652 532016 107704
rect 503904 107516 503956 107568
rect 504364 107516 504416 107568
rect 82636 106700 82688 106752
rect 82912 106700 82964 106752
rect 502984 105476 503036 105528
rect 504456 105476 504508 105528
rect 83004 104796 83056 104848
rect 512828 104796 512880 104848
rect 82912 104728 82964 104780
rect 504548 103504 504600 103556
rect 511356 103504 511408 103556
rect 9128 102688 9180 102740
rect 82728 102756 82780 102808
rect 81072 102688 81124 102740
rect 72976 102620 73028 102672
rect 74172 102552 74224 102604
rect 173992 102552 174044 102604
rect 201500 102688 201552 102740
rect 370504 102620 370556 102672
rect 509240 102824 509292 102876
rect 523408 102756 523460 102808
rect 416688 102663 416740 102672
rect 416688 102629 416697 102663
rect 416697 102629 416731 102663
rect 416731 102629 416740 102663
rect 416688 102620 416740 102629
rect 83096 102416 83148 102468
rect 83648 102416 83700 102468
rect 79876 102348 79928 102400
rect 84844 102348 84896 102400
rect 83372 102280 83424 102332
rect 125508 102484 125560 102536
rect 133696 102484 133748 102536
rect 149060 102416 149112 102468
rect 79692 102212 79744 102264
rect 79876 102212 79928 102264
rect 74264 102076 74316 102128
rect 510896 102076 510948 102128
rect 499488 101940 499540 101992
rect 513840 101940 513892 101992
rect 81992 101872 82044 101924
rect 106464 101872 106516 101924
rect 488448 101872 488500 101924
rect 508504 101872 508556 101924
rect 83648 101804 83700 101856
rect 107660 101804 107712 101856
rect 187792 101804 187844 101856
rect 480076 101804 480128 101856
rect 502524 101804 502576 101856
rect 67180 101736 67232 101788
rect 93952 101736 94004 101788
rect 487068 101736 487120 101788
rect 509792 101736 509844 101788
rect 56508 101668 56560 101720
rect 88524 101668 88576 101720
rect 484308 101668 484360 101720
rect 513932 101668 513984 101720
rect 71596 101600 71648 101652
rect 103612 101600 103664 101652
rect 453948 101600 454000 101652
rect 505652 101600 505704 101652
rect 75552 101532 75604 101584
rect 117320 101532 117372 101584
rect 439504 101532 439556 101584
rect 504364 101532 504416 101584
rect 80980 101464 81032 101516
rect 128360 101464 128412 101516
rect 198740 101464 198792 101516
rect 512460 101464 512512 101516
rect 85580 101396 85632 101448
rect 495256 101396 495308 101448
rect 500868 101396 500920 101448
rect 519176 101396 519228 101448
rect 82176 101260 82228 101312
rect 85580 101260 85632 101312
rect 88340 100852 88392 100904
rect 419448 100852 419500 100904
rect 39304 100784 39356 100836
rect 166448 100784 166500 100836
rect 245568 100784 245620 100836
rect 511448 100784 511500 100836
rect 72608 100716 72660 100768
rect 467840 100716 467892 100768
rect 513288 100716 513340 100768
rect 520924 100716 520976 100768
rect 11704 100648 11756 100700
rect 285128 100648 285180 100700
rect 292488 100648 292540 100700
rect 514116 100648 514168 100700
rect 68376 100580 68428 100632
rect 322112 100580 322164 100632
rect 327080 100580 327132 100632
rect 516784 100580 516836 100632
rect 82544 100512 82596 100564
rect 84936 100512 84988 100564
rect 329472 100512 329524 100564
rect 359096 100512 359148 100564
rect 360108 100512 360160 100564
rect 410984 100512 411036 100564
rect 560944 100512 560996 100564
rect 68836 100444 68888 100496
rect 186136 100444 186188 100496
rect 218336 100444 218388 100496
rect 219348 100444 219400 100496
rect 230664 100444 230716 100496
rect 231768 100444 231820 100496
rect 255320 100444 255372 100496
rect 256608 100444 256660 100496
rect 267832 100444 267884 100496
rect 269028 100444 269080 100496
rect 280160 100444 280212 100496
rect 281448 100444 281500 100496
rect 388904 100444 388956 100496
rect 511264 100444 511316 100496
rect 69756 100376 69808 100428
rect 176384 100376 176436 100428
rect 401232 100376 401284 100428
rect 520464 100376 520516 100428
rect 71504 100308 71556 100360
rect 164056 100308 164108 100360
rect 403624 100308 403676 100360
rect 515404 100308 515456 100360
rect 70308 100240 70360 100292
rect 131856 100240 131908 100292
rect 136824 100240 136876 100292
rect 137928 100240 137980 100292
rect 206008 100240 206060 100292
rect 206928 100240 206980 100292
rect 207664 100240 207716 100292
rect 277584 100240 277636 100292
rect 286324 100240 286376 100292
rect 314752 100240 314804 100292
rect 327724 100240 327776 100292
rect 341800 100240 341852 100292
rect 376392 100240 376444 100292
rect 419448 100240 419500 100292
rect 440792 100240 440844 100292
rect 455512 100240 455564 100292
rect 456708 100240 456760 100292
rect 475384 100240 475436 100292
rect 509976 100240 510028 100292
rect 75828 100172 75880 100224
rect 112168 100172 112220 100224
rect 114560 100172 114612 100224
rect 115848 100172 115900 100224
rect 124864 100172 124916 100224
rect 126888 100172 126940 100224
rect 240784 100172 240836 100224
rect 356704 100172 356756 100224
rect 370596 100172 370648 100224
rect 408592 100172 408644 100224
rect 81348 100104 81400 100156
rect 89904 100104 89956 100156
rect 91008 100104 91060 100156
rect 99656 100104 99708 100156
rect 100668 100104 100720 100156
rect 117964 100104 118016 100156
rect 159088 100104 159140 100156
rect 186964 100104 187016 100156
rect 213368 100104 213420 100156
rect 261484 100104 261536 100156
rect 393688 100104 393740 100156
rect 83556 100036 83608 100088
rect 99472 100036 99524 100088
rect 142804 100036 142856 100088
rect 198648 100036 198700 100088
rect 225604 100036 225656 100088
rect 240600 100036 240652 100088
rect 251824 100036 251876 100088
rect 406200 100036 406252 100088
rect 478788 100036 478840 100088
rect 505744 100036 505796 100088
rect 81440 99968 81492 100020
rect 110420 99968 110472 100020
rect 131764 99968 131816 100020
rect 139216 99968 139268 100020
rect 149704 99968 149756 100020
rect 260288 99968 260340 100020
rect 302148 99968 302200 100020
rect 521844 99968 521896 100020
rect 477776 99900 477828 99952
rect 478696 99900 478748 99952
rect 102232 99832 102284 99884
rect 103428 99832 103480 99884
rect 121920 99696 121972 99748
rect 122748 99696 122800 99748
rect 265256 99628 265308 99680
rect 266268 99628 266320 99680
rect 287520 99356 287572 99408
rect 288348 99356 288400 99408
rect 315304 99356 315356 99408
rect 317144 99356 317196 99408
rect 323584 99356 323636 99408
rect 324504 99356 324556 99408
rect 334440 99356 334492 99408
rect 335268 99356 335320 99408
rect 374000 99356 374052 99408
rect 375288 99356 375340 99408
rect 381360 99356 381412 99408
rect 382188 99356 382240 99408
rect 383936 99356 383988 99408
rect 384948 99356 385000 99408
rect 494704 99356 494756 99408
rect 500040 99356 500092 99408
rect 183744 99288 183796 99340
rect 184848 99288 184900 99340
rect 280528 99331 280580 99340
rect 280528 99297 280537 99331
rect 280537 99297 280571 99331
rect 280571 99297 280580 99331
rect 280528 99288 280580 99297
rect 469128 99288 469180 99340
rect 502892 99288 502944 99340
rect 503076 99288 503128 99340
rect 513288 99288 513340 99340
rect 78404 99220 78456 99272
rect 132592 99220 132644 99272
rect 486976 99220 487028 99272
rect 523316 99220 523368 99272
rect 70216 99152 70268 99204
rect 142160 99152 142212 99204
rect 419448 99152 419500 99204
rect 518992 99152 519044 99204
rect 75644 99084 75696 99136
rect 149060 99084 149112 99136
rect 354588 99084 354640 99136
rect 512276 99084 512328 99136
rect 71412 99016 71464 99068
rect 146300 99016 146352 99068
rect 331128 99016 331180 99068
rect 520648 99016 520700 99068
rect 66168 98948 66220 99000
rect 167000 98948 167052 99000
rect 306288 98948 306340 99000
rect 510804 98948 510856 99000
rect 80704 98880 80756 98932
rect 193220 98880 193272 98932
rect 284208 98880 284260 98932
rect 512552 98880 512604 98932
rect 61752 98812 61804 98864
rect 179420 98812 179472 98864
rect 251088 98812 251140 98864
rect 503996 98812 504048 98864
rect 77944 98744 77996 98796
rect 195980 98744 196032 98796
rect 241428 98744 241480 98796
rect 515128 98744 515180 98796
rect 67272 98676 67324 98728
rect 218060 98676 218112 98728
rect 227628 98676 227680 98728
rect 509700 98676 509752 98728
rect 81164 98608 81216 98660
rect 207020 98608 207072 98660
rect 216588 98608 216640 98660
rect 519084 98608 519136 98660
rect 187700 97996 187752 98048
rect 188436 97996 188488 98048
rect 25504 97928 25556 97980
rect 129464 97928 129516 97980
rect 146760 97928 146812 97980
rect 567844 97928 567896 97980
rect 43444 97860 43496 97912
rect 346768 97860 346820 97912
rect 69848 97792 69900 97844
rect 178776 97792 178828 97844
rect 491300 97588 491352 97640
rect 503076 97588 503128 97640
rect 487804 97520 487856 97572
rect 523224 97520 523276 97572
rect 463608 97452 463660 97504
rect 505376 97452 505428 97504
rect 61844 97384 61896 97436
rect 81900 97384 81952 97436
rect 365628 97384 365680 97436
rect 517796 97384 517848 97436
rect 57888 97316 57940 97368
rect 81440 97316 81492 97368
rect 355968 97316 356020 97368
rect 520556 97316 520608 97368
rect 79784 97248 79836 97300
rect 212540 97248 212592 97300
rect 329748 97248 329800 97300
rect 516416 97248 516468 97300
rect 212264 96636 212316 96688
rect 212356 96636 212408 96688
rect 356520 96679 356572 96688
rect 356520 96645 356529 96679
rect 356529 96645 356563 96679
rect 356563 96645 356572 96679
rect 356520 96636 356572 96645
rect 168840 96568 168892 96620
rect 176752 96568 176804 96620
rect 565084 96568 565136 96620
rect 32404 96500 32456 96552
rect 413560 96500 413612 96552
rect 456616 96500 456668 96552
rect 191104 96432 191156 96484
rect 512644 96432 512696 96484
rect 440148 96364 440200 96416
rect 516324 96364 516376 96416
rect 398748 96296 398800 96348
rect 501788 96296 501840 96348
rect 519268 96296 519320 96348
rect 389088 96228 389140 96280
rect 510988 96228 511040 96280
rect 349068 96160 349120 96212
rect 508412 96160 508464 96212
rect 326988 96092 327040 96144
rect 515036 96092 515088 96144
rect 275928 96024 275980 96076
rect 510712 96024 510764 96076
rect 195888 95956 195940 96008
rect 516508 95956 516560 96008
rect 83372 95888 83424 95940
rect 151728 95888 151780 95940
rect 520832 95888 520884 95940
rect 512736 95208 512788 95260
rect 484216 95004 484268 95056
rect 487804 95004 487856 95056
rect 481732 94936 481784 94988
rect 484492 94936 484544 94988
rect 83464 94664 83516 94716
rect 492772 94664 492824 94716
rect 523132 94664 523184 94716
rect 83096 94528 83148 94580
rect 83464 94528 83516 94580
rect 393228 94596 393280 94648
rect 505560 94596 505612 94648
rect 367008 94528 367060 94580
rect 501604 94528 501656 94580
rect 79140 94460 79192 94512
rect 567200 94460 567252 94512
rect 487804 93848 487856 93900
rect 491300 93848 491352 93900
rect 3424 93780 3476 93832
rect 15936 93780 15988 93832
rect 433248 93712 433300 93764
rect 507124 93712 507176 93764
rect 522120 93644 522172 93696
rect 386328 93576 386380 93628
rect 521752 93576 521804 93628
rect 249708 93508 249760 93560
rect 516692 93508 516744 93560
rect 220728 93440 220780 93492
rect 505192 93440 505244 93492
rect 217968 93372 218020 93424
rect 521936 93372 521988 93424
rect 173808 93304 173860 93356
rect 196072 93304 196124 93356
rect 200028 93304 200080 93356
rect 520740 93304 520792 93356
rect 122840 93236 122892 93288
rect 186228 93236 186280 93288
rect 515312 93236 515364 93288
rect 183468 93168 183520 93220
rect 518072 93168 518124 93220
rect 59268 93100 59320 93152
rect 78680 93100 78732 93152
rect 146208 93100 146260 93152
rect 522028 93100 522080 93152
rect 488540 91944 488592 91996
rect 492772 91944 492824 91996
rect 436008 91876 436060 91928
rect 507952 91876 508004 91928
rect 278688 91808 278740 91860
rect 505100 91808 505152 91860
rect 79416 91740 79468 91792
rect 444380 91740 444432 91792
rect 480720 91060 480772 91112
rect 481732 91060 481784 91112
rect 483020 91060 483072 91112
rect 488632 91060 488684 91112
rect 298008 90380 298060 90432
rect 519360 90380 519412 90432
rect 76656 90312 76708 90364
rect 335360 90312 335412 90364
rect 356520 89700 356572 89752
rect 176752 89675 176804 89684
rect 176752 89641 176761 89675
rect 176761 89641 176795 89675
rect 176795 89641 176804 89675
rect 176752 89632 176804 89641
rect 356612 89564 356664 89616
rect 83280 89403 83332 89412
rect 83280 89369 83289 89403
rect 83289 89369 83323 89403
rect 83323 89369 83332 89403
rect 83280 89360 83332 89369
rect 78128 89020 78180 89072
rect 305000 89020 305052 89072
rect 280068 88952 280120 89004
rect 508044 88952 508096 89004
rect 484492 88612 484544 88664
rect 487804 88612 487856 88664
rect 482284 88476 482336 88528
rect 484216 88476 484268 88528
rect 84936 87592 84988 87644
rect 138020 87592 138072 87644
rect 176476 87592 176528 87644
rect 187700 87592 187752 87644
rect 293868 87592 293920 87644
rect 506756 87592 506808 87644
rect 151544 86980 151596 87032
rect 151636 86980 151688 87032
rect 411168 87023 411220 87032
rect 411168 86989 411177 87023
rect 411177 86989 411211 87023
rect 411211 86989 411220 87023
rect 411168 86980 411220 86989
rect 512736 86980 512788 87032
rect 512828 86980 512880 87032
rect 176660 86912 176712 86964
rect 176752 86912 176804 86964
rect 198556 86912 198608 86964
rect 280528 86912 280580 86964
rect 483756 86912 483808 86964
rect 484492 86912 484544 86964
rect 487252 86640 487304 86692
rect 488540 86640 488592 86692
rect 201408 86368 201460 86420
rect 274640 86368 274692 86420
rect 253848 86300 253900 86352
rect 504272 86300 504324 86352
rect 75460 86232 75512 86284
rect 342260 86232 342312 86284
rect 473268 86232 473320 86284
rect 528560 86232 528612 86284
rect 477500 85552 477552 85604
rect 480720 85552 480772 85604
rect 79784 85527 79836 85536
rect 79784 85493 79793 85527
rect 79793 85493 79827 85527
rect 79827 85493 79836 85527
rect 79784 85484 79836 85493
rect 512828 85527 512880 85536
rect 512828 85493 512837 85527
rect 512837 85493 512871 85527
rect 512871 85493 512880 85527
rect 512828 85484 512880 85493
rect 558184 85484 558236 85536
rect 564440 85484 564492 85536
rect 77024 84872 77076 84924
rect 155960 84872 156012 84924
rect 102048 84804 102100 84856
rect 261484 84804 261536 84856
rect 314568 84804 314620 84856
rect 508228 84804 508280 84856
rect 476120 84124 476172 84176
rect 482928 84192 482980 84244
rect 78220 83580 78272 83632
rect 287060 83580 287112 83632
rect 210884 83512 210936 83564
rect 502708 83512 502760 83564
rect 79232 83444 79284 83496
rect 451280 83444 451332 83496
rect 481088 82832 481140 82884
rect 483756 82832 483808 82884
rect 485504 82832 485556 82884
rect 487252 82832 487304 82884
rect 89904 82084 89956 82136
rect 90088 82084 90140 82136
rect 211068 82084 211120 82136
rect 396080 82084 396132 82136
rect 478880 81404 478932 81456
rect 481088 81404 481140 81456
rect 151544 81107 151596 81116
rect 151544 81073 151553 81107
rect 151553 81073 151587 81107
rect 151587 81073 151596 81107
rect 151544 81064 151596 81073
rect 228916 80656 228968 80708
rect 505468 80656 505520 80708
rect 356612 80044 356664 80096
rect 474648 80044 474700 80096
rect 476120 80044 476172 80096
rect 356704 79908 356756 79960
rect 271788 79364 271840 79416
rect 506480 79364 506532 79416
rect 76840 79296 76892 79348
rect 378140 79296 378192 79348
rect 473268 79296 473320 79348
rect 477408 79296 477460 79348
rect 483664 78208 483716 78260
rect 485504 78208 485556 78260
rect 75368 78072 75420 78124
rect 263600 78072 263652 78124
rect 471244 78072 471296 78124
rect 474648 78072 474700 78124
rect 157248 78004 157300 78056
rect 230480 78004 230532 78056
rect 245568 78004 245620 78056
rect 501880 78004 501932 78056
rect 194508 77936 194560 77988
rect 481640 77936 481692 77988
rect 475384 77528 475436 77580
rect 478880 77528 478932 77580
rect 151544 77367 151596 77376
rect 151544 77333 151553 77367
rect 151553 77333 151587 77367
rect 151587 77333 151596 77367
rect 151544 77324 151596 77333
rect 198464 77299 198516 77308
rect 198464 77265 198473 77299
rect 198473 77265 198507 77299
rect 198507 77265 198516 77299
rect 198464 77256 198516 77265
rect 280436 77299 280488 77308
rect 280436 77265 280445 77299
rect 280445 77265 280479 77299
rect 280479 77265 280488 77299
rect 280436 77256 280488 77265
rect 72516 77188 72568 77240
rect 580172 77188 580224 77240
rect 151452 77163 151504 77172
rect 151452 77129 151461 77163
rect 151461 77129 151495 77163
rect 151495 77129 151504 77163
rect 151452 77120 151504 77129
rect 176844 77120 176896 77172
rect 198464 77163 198516 77172
rect 198464 77129 198473 77163
rect 198473 77129 198507 77163
rect 198507 77129 198516 77163
rect 198464 77120 198516 77129
rect 356704 77163 356756 77172
rect 356704 77129 356713 77163
rect 356713 77129 356747 77163
rect 356747 77129 356756 77163
rect 356704 77120 356756 77129
rect 411168 77163 411220 77172
rect 411168 77129 411177 77163
rect 411177 77129 411211 77163
rect 411211 77129 411220 77163
rect 411168 77120 411220 77129
rect 470600 76712 470652 76764
rect 473268 76712 473320 76764
rect 85488 76576 85540 76628
rect 242900 76576 242952 76628
rect 184848 76508 184900 76560
rect 360200 76508 360252 76560
rect 79968 75896 80020 75948
rect 512828 75939 512880 75948
rect 512828 75905 512837 75939
rect 512837 75905 512871 75939
rect 512871 75905 512880 75939
rect 512828 75896 512880 75905
rect 480904 75828 480956 75880
rect 482284 75828 482336 75880
rect 119988 75148 120040 75200
rect 204260 75148 204312 75200
rect 233148 75148 233200 75200
rect 309232 75148 309284 75200
rect 107568 73924 107620 73976
rect 133880 73924 133932 73976
rect 240048 73924 240100 73976
rect 385040 73924 385092 73976
rect 76564 73856 76616 73908
rect 171140 73856 171192 73908
rect 332508 73856 332560 73908
rect 501696 73856 501748 73908
rect 19248 73788 19300 73840
rect 338120 73788 338172 73840
rect 342168 72496 342220 72548
rect 489920 72496 489972 72548
rect 84016 72428 84068 72480
rect 553400 72428 553452 72480
rect 469312 71952 469364 72004
rect 471244 71952 471296 72004
rect 226248 71068 226300 71120
rect 284300 71068 284352 71120
rect 364156 71068 364208 71120
rect 371240 71068 371292 71120
rect 93768 71000 93820 71052
rect 365720 71000 365772 71052
rect 375196 71000 375248 71052
rect 418160 71000 418212 71052
rect 472440 70592 472492 70644
rect 475384 70592 475436 70644
rect 83648 70456 83700 70508
rect 83648 70320 83700 70372
rect 89904 70388 89956 70440
rect 280252 70388 280304 70440
rect 280344 70320 280396 70372
rect 356796 70252 356848 70304
rect 89812 70184 89864 70236
rect 338028 69708 338080 69760
rect 496820 69708 496872 69760
rect 74080 69640 74132 69692
rect 445760 69640 445812 69692
rect 469864 69232 469916 69284
rect 472440 69232 472492 69284
rect 468944 69028 468996 69080
rect 470508 69028 470560 69080
rect 128268 68416 128320 68468
rect 289820 68416 289872 68468
rect 81716 68348 81768 68400
rect 320180 68348 320232 68400
rect 348976 68348 349028 68400
rect 502616 68348 502668 68400
rect 96528 68280 96580 68332
rect 504180 68280 504232 68332
rect 79784 67600 79836 67652
rect 79968 67600 80020 67652
rect 151544 67600 151596 67652
rect 176752 67643 176804 67652
rect 176752 67609 176761 67643
rect 176761 67609 176795 67643
rect 176795 67609 176804 67643
rect 176752 67600 176804 67609
rect 198556 67600 198608 67652
rect 411168 67643 411220 67652
rect 411168 67609 411177 67643
rect 411177 67609 411211 67643
rect 411211 67609 411220 67643
rect 411168 67600 411220 67609
rect 140780 67532 140832 67584
rect 140872 67532 140924 67584
rect 467104 67464 467156 67516
rect 469312 67464 469364 67516
rect 467196 67192 467248 67244
rect 468944 67192 468996 67244
rect 256516 66920 256568 66972
rect 303620 66920 303672 66972
rect 371148 66920 371200 66972
rect 378232 66920 378284 66972
rect 119988 66852 120040 66904
rect 508320 66852 508372 66904
rect 83372 66215 83424 66224
rect 83372 66181 83381 66215
rect 83381 66181 83415 66215
rect 83415 66181 83424 66215
rect 83372 66172 83424 66181
rect 512828 66215 512880 66224
rect 512828 66181 512837 66215
rect 512837 66181 512871 66215
rect 512871 66181 512880 66215
rect 512828 66172 512880 66181
rect 360108 65628 360160 65680
rect 433340 65628 433392 65680
rect 315948 65560 316000 65612
rect 505284 65560 505336 65612
rect 106188 65492 106240 65544
rect 208400 65492 208452 65544
rect 210976 65492 211028 65544
rect 504088 65492 504140 65544
rect 3332 64812 3384 64864
rect 33784 64812 33836 64864
rect 519544 64812 519596 64864
rect 579804 64812 579856 64864
rect 88248 64132 88300 64184
rect 509608 64132 509660 64184
rect 22008 62840 22060 62892
rect 240784 62840 240836 62892
rect 165528 62772 165580 62824
rect 506664 62772 506716 62824
rect 476764 62636 476816 62688
rect 480904 62636 480956 62688
rect 465172 62092 465224 62144
rect 467196 62092 467248 62144
rect 222108 61616 222160 61668
rect 269120 61616 269172 61668
rect 75276 61548 75328 61600
rect 267740 61548 267792 61600
rect 107476 61480 107528 61532
rect 311992 61480 312044 61532
rect 260748 61412 260800 61464
rect 502340 61412 502392 61464
rect 99288 61344 99340 61396
rect 509516 61344 509568 61396
rect 89812 60732 89864 60784
rect 79692 60664 79744 60716
rect 79876 60664 79928 60716
rect 151544 60800 151596 60852
rect 198556 60800 198608 60852
rect 482008 60732 482060 60784
rect 483664 60732 483716 60784
rect 89996 60664 90048 60716
rect 151452 60664 151504 60716
rect 198464 60664 198516 60716
rect 333888 60120 333940 60172
rect 456800 60120 456852 60172
rect 45468 60052 45520 60104
rect 370596 60052 370648 60104
rect 467748 60052 467800 60104
rect 494060 60052 494112 60104
rect 97908 59984 97960 60036
rect 504364 59984 504416 60036
rect 144644 58760 144696 58812
rect 396172 58760 396224 58812
rect 68836 58692 68888 58744
rect 323584 58692 323636 58744
rect 219256 58624 219308 58676
rect 506572 58624 506624 58676
rect 445576 57944 445628 57996
rect 445668 57944 445720 57996
rect 79876 57919 79928 57928
rect 79876 57885 79885 57919
rect 79885 57885 79919 57919
rect 79919 57885 79928 57919
rect 79876 57876 79928 57885
rect 89996 57876 90048 57928
rect 140688 57876 140740 57928
rect 140780 57876 140832 57928
rect 144736 57919 144788 57928
rect 144736 57885 144745 57919
rect 144745 57885 144779 57919
rect 144779 57885 144788 57919
rect 144736 57876 144788 57885
rect 176844 57876 176896 57928
rect 198464 57919 198516 57928
rect 198464 57885 198473 57919
rect 198473 57885 198507 57919
rect 198507 57885 198516 57919
rect 198464 57876 198516 57885
rect 212448 57919 212500 57928
rect 212448 57885 212457 57919
rect 212457 57885 212491 57919
rect 212491 57885 212500 57919
rect 212448 57876 212500 57885
rect 280436 57876 280488 57928
rect 333888 57919 333940 57928
rect 333888 57885 333897 57919
rect 333897 57885 333931 57919
rect 333931 57885 333940 57919
rect 333888 57876 333940 57885
rect 356612 57919 356664 57928
rect 356612 57885 356621 57919
rect 356621 57885 356655 57919
rect 356655 57885 356664 57919
rect 356612 57876 356664 57885
rect 411168 57919 411220 57928
rect 411168 57885 411177 57919
rect 411177 57885 411211 57919
rect 411211 57885 411220 57919
rect 411168 57876 411220 57885
rect 83556 57808 83608 57860
rect 462412 57808 462464 57860
rect 465172 57808 465224 57860
rect 467840 57740 467892 57792
rect 469864 57740 469916 57792
rect 344836 57264 344888 57316
rect 527180 57264 527232 57316
rect 83648 57196 83700 57248
rect 376760 57196 376812 57248
rect 380808 57196 380860 57248
rect 431960 57196 432012 57248
rect 512828 56627 512880 56636
rect 512828 56593 512837 56627
rect 512837 56593 512871 56627
rect 512871 56593 512880 56627
rect 512828 56584 512880 56593
rect 140688 56559 140740 56568
rect 140688 56525 140697 56559
rect 140697 56525 140731 56559
rect 140731 56525 140740 56559
rect 140688 56516 140740 56525
rect 81532 55972 81584 56024
rect 350632 55972 350684 56024
rect 354496 55972 354548 56024
rect 419540 55972 419592 56024
rect 478880 55972 478932 56024
rect 482008 55972 482060 56024
rect 220636 55904 220688 55956
rect 505100 55904 505152 55956
rect 15108 55836 15160 55888
rect 131764 55836 131816 55888
rect 136548 55836 136600 55888
rect 503812 55836 503864 55888
rect 472900 53864 472952 53916
rect 478880 53864 478932 53916
rect 464344 53796 464396 53848
rect 467840 53796 467892 53848
rect 391756 53048 391808 53100
rect 487160 53048 487212 53100
rect 467840 52436 467892 52488
rect 472900 52436 472952 52488
rect 474004 52436 474056 52488
rect 476764 52436 476816 52488
rect 80888 51688 80940 51740
rect 382280 51688 382332 51740
rect 384948 51688 385000 51740
rect 476120 51688 476172 51740
rect 3424 51008 3476 51060
rect 71044 51008 71096 51060
rect 151452 51008 151504 51060
rect 151636 51008 151688 51060
rect 79876 50915 79928 50924
rect 79876 50881 79885 50915
rect 79885 50881 79919 50915
rect 79919 50881 79928 50915
rect 79876 50872 79928 50881
rect 357256 50396 357308 50448
rect 415400 50396 415452 50448
rect 78496 50328 78548 50380
rect 234620 50328 234672 50380
rect 250996 50328 251048 50380
rect 393320 50328 393372 50380
rect 461584 49648 461636 49700
rect 462412 49648 462464 49700
rect 382188 49104 382240 49156
rect 540980 49104 541032 49156
rect 81624 49036 81676 49088
rect 404360 49036 404412 49088
rect 153108 48968 153160 49020
rect 507032 48968 507084 49020
rect 89904 48331 89956 48340
rect 89904 48297 89913 48331
rect 89913 48297 89947 48331
rect 89947 48297 89956 48331
rect 89904 48288 89956 48297
rect 144736 48331 144788 48340
rect 144736 48297 144745 48331
rect 144745 48297 144779 48331
rect 144779 48297 144788 48331
rect 144736 48288 144788 48297
rect 176752 48331 176804 48340
rect 176752 48297 176761 48331
rect 176761 48297 176795 48331
rect 176795 48297 176804 48331
rect 176752 48288 176804 48297
rect 198556 48288 198608 48340
rect 210976 48331 211028 48340
rect 210976 48297 210985 48331
rect 210985 48297 211019 48331
rect 211019 48297 211028 48331
rect 210976 48288 211028 48297
rect 212448 48331 212500 48340
rect 212448 48297 212457 48331
rect 212457 48297 212491 48331
rect 212491 48297 212500 48331
rect 212448 48288 212500 48297
rect 280344 48331 280396 48340
rect 280344 48297 280353 48331
rect 280353 48297 280387 48331
rect 280387 48297 280396 48331
rect 280344 48288 280396 48297
rect 333888 48331 333940 48340
rect 333888 48297 333897 48331
rect 333897 48297 333931 48331
rect 333931 48297 333940 48331
rect 333888 48288 333940 48297
rect 356704 48288 356756 48340
rect 411168 48331 411220 48340
rect 411168 48297 411177 48331
rect 411177 48297 411211 48331
rect 411211 48297 411220 48331
rect 411168 48288 411220 48297
rect 151636 48220 151688 48272
rect 465816 47880 465868 47932
rect 467840 47880 467892 47932
rect 90916 47540 90968 47592
rect 200120 47540 200172 47592
rect 140780 46928 140832 46980
rect 210976 46971 211028 46980
rect 210976 46937 210985 46971
rect 210985 46937 211019 46971
rect 211019 46937 211028 46971
rect 210976 46928 211028 46937
rect 512828 46903 512880 46912
rect 512828 46869 512837 46903
rect 512837 46869 512871 46903
rect 512871 46869 512880 46903
rect 512828 46860 512880 46869
rect 83372 46248 83424 46300
rect 237472 46248 237524 46300
rect 281448 46248 281500 46300
rect 333980 46248 334032 46300
rect 335268 46248 335320 46300
rect 429200 46248 429252 46300
rect 155868 46180 155920 46232
rect 492680 46180 492732 46232
rect 140780 45543 140832 45552
rect 140780 45509 140789 45543
rect 140789 45509 140823 45543
rect 140823 45509 140832 45543
rect 140780 45500 140832 45509
rect 103428 44888 103480 44940
rect 425060 44888 425112 44940
rect 223488 44820 223540 44872
rect 565820 44820 565872 44872
rect 456064 44004 456116 44056
rect 461584 44140 461636 44192
rect 462688 43528 462740 43580
rect 464344 43528 464396 43580
rect 110236 43460 110288 43512
rect 506940 43460 506992 43512
rect 78036 43392 78088 43444
rect 538220 43392 538272 43444
rect 463792 42780 463844 42832
rect 465816 42780 465868 42832
rect 235908 42100 235960 42152
rect 492680 42100 492732 42152
rect 79508 42032 79560 42084
rect 358820 42032 358872 42084
rect 469312 42032 469364 42084
rect 474004 42032 474056 42084
rect 198556 41420 198608 41472
rect 460204 41420 460256 41472
rect 462688 41420 462740 41472
rect 89812 41352 89864 41404
rect 89996 41352 90048 41404
rect 198464 41352 198516 41404
rect 549904 41352 549956 41404
rect 580172 41352 580224 41404
rect 76748 40740 76800 40792
rect 367100 40740 367152 40792
rect 391848 40740 391900 40792
rect 441620 40740 441672 40792
rect 104808 40672 104860 40724
rect 494060 40672 494112 40724
rect 465724 40060 465776 40112
rect 469312 40060 469364 40112
rect 461584 39856 461636 39908
rect 463792 39856 463844 39908
rect 360844 39380 360896 39432
rect 370504 39380 370556 39432
rect 307576 39312 307628 39364
rect 520464 39312 520516 39364
rect 151544 38675 151596 38684
rect 151544 38641 151553 38675
rect 151553 38641 151587 38675
rect 151587 38641 151596 38675
rect 151544 38632 151596 38641
rect 445576 38632 445628 38684
rect 445668 38632 445720 38684
rect 144736 38607 144788 38616
rect 144736 38573 144745 38607
rect 144745 38573 144779 38607
rect 144779 38573 144788 38607
rect 144736 38564 144788 38573
rect 176844 38564 176896 38616
rect 198464 38607 198516 38616
rect 198464 38573 198473 38607
rect 198473 38573 198507 38607
rect 198507 38573 198516 38607
rect 198464 38564 198516 38573
rect 280436 38564 280488 38616
rect 161388 38020 161440 38072
rect 356888 38020 356940 38072
rect 228824 37952 228876 38004
rect 501512 37952 501564 38004
rect 79876 37884 79928 37936
rect 436100 37884 436152 37936
rect 210976 37272 211028 37324
rect 211068 37272 211120 37324
rect 512828 37315 512880 37324
rect 512828 37281 512837 37315
rect 512837 37281 512871 37315
rect 512871 37281 512880 37315
rect 512828 37272 512880 37281
rect 140872 35912 140924 35964
rect 458272 34484 458324 34536
rect 461584 34484 461636 34536
rect 462964 34484 463016 34536
rect 465724 34484 465776 34536
rect 451188 33804 451240 33856
rect 574744 33804 574796 33856
rect 248236 33736 248288 33788
rect 495440 33736 495492 33788
rect 182088 32512 182140 32564
rect 252560 32512 252612 32564
rect 219348 32444 219400 32496
rect 294052 32444 294104 32496
rect 353300 32444 353352 32496
rect 360844 32444 360896 32496
rect 78588 32376 78640 32428
rect 223580 32376 223632 32428
rect 256608 32376 256660 32428
rect 460940 32376 460992 32428
rect 89996 31807 90048 31816
rect 89996 31773 90005 31807
rect 90005 31773 90039 31807
rect 90039 31773 90048 31807
rect 89996 31764 90048 31773
rect 176752 31739 176804 31748
rect 176752 31705 176761 31739
rect 176761 31705 176795 31739
rect 176795 31705 176804 31739
rect 176752 31696 176804 31705
rect 280344 31739 280396 31748
rect 280344 31705 280353 31739
rect 280353 31705 280387 31739
rect 280387 31705 280396 31739
rect 280344 31696 280396 31705
rect 198556 31628 198608 31680
rect 237196 31016 237248 31068
rect 311900 31016 311952 31068
rect 409788 31016 409840 31068
rect 469220 31016 469272 31068
rect 457444 30200 457496 30252
rect 458272 30200 458324 30252
rect 9588 29724 9640 29776
rect 207664 29724 207716 29776
rect 297824 29724 297876 29776
rect 430580 29724 430632 29776
rect 184848 29656 184900 29708
rect 484400 29656 484452 29708
rect 204076 29588 204128 29640
rect 506848 29588 506900 29640
rect 553124 29180 553176 29232
rect 560208 29180 560260 29232
rect 89904 29044 89956 29096
rect 144736 29019 144788 29028
rect 144736 28985 144745 29019
rect 144745 28985 144779 29019
rect 144779 28985 144788 29019
rect 144736 28976 144788 28985
rect 411168 28908 411220 28960
rect 411352 28908 411404 28960
rect 103428 28364 103480 28416
rect 420920 28364 420972 28416
rect 423588 28364 423640 28416
rect 440240 28364 440292 28416
rect 137928 28296 137980 28348
rect 491300 28296 491352 28348
rect 144828 28228 144880 28280
rect 581092 28228 581144 28280
rect 89812 27591 89864 27600
rect 89812 27557 89821 27591
rect 89821 27557 89855 27591
rect 89855 27557 89864 27591
rect 89812 27548 89864 27557
rect 210976 27591 211028 27600
rect 210976 27557 210985 27591
rect 210985 27557 211019 27591
rect 211019 27557 211028 27591
rect 210976 27548 211028 27557
rect 512828 27548 512880 27600
rect 351184 27208 351236 27260
rect 353300 27208 353352 27260
rect 38568 26936 38620 26988
rect 153200 26936 153252 26988
rect 266268 26936 266320 26988
rect 401600 26936 401652 26988
rect 151452 26868 151504 26920
rect 539600 26868 539652 26920
rect 97908 25712 97960 25764
rect 251824 25712 251876 25764
rect 246948 25644 247000 25696
rect 462320 25644 462372 25696
rect 100668 25576 100720 25628
rect 408500 25576 408552 25628
rect 20628 25508 20680 25560
rect 91100 25508 91152 25560
rect 110328 25508 110380 25560
rect 550640 25508 550692 25560
rect 216496 24148 216548 24200
rect 233332 24148 233384 24200
rect 75736 24080 75788 24132
rect 281540 24080 281592 24132
rect 465724 23468 465776 23520
rect 467104 23468 467156 23520
rect 26148 23128 26200 23180
rect 28264 23128 28316 23180
rect 28908 22788 28960 22840
rect 142804 22788 142856 22840
rect 269028 22788 269080 22840
rect 400220 22788 400272 22840
rect 81808 22720 81860 22772
rect 552020 22720 552072 22772
rect 140872 22652 140924 22704
rect 452568 22176 452620 22228
rect 456064 22176 456116 22228
rect 455420 22108 455472 22160
rect 457444 22108 457496 22160
rect 3148 22040 3200 22092
rect 514852 22040 514904 22092
rect 89996 21904 90048 21956
rect 297916 21428 297968 21480
rect 576860 21428 576912 21480
rect 95148 21360 95200 21412
rect 473360 21360 473412 21412
rect 478696 21360 478748 21412
rect 484400 21360 484452 21412
rect 282828 20068 282880 20120
rect 531320 20068 531372 20120
rect 79600 20000 79652 20052
rect 338212 20000 338264 20052
rect 449164 20000 449216 20052
rect 452568 20000 452620 20052
rect 21916 19932 21968 19984
rect 117964 19932 118016 19984
rect 122748 19932 122800 19984
rect 169760 19932 169812 19984
rect 173716 19932 173768 19984
rect 456800 19932 456852 19984
rect 445576 19320 445628 19372
rect 445668 19320 445720 19372
rect 144736 19295 144788 19304
rect 144736 19261 144745 19295
rect 144745 19261 144779 19295
rect 144779 19261 144788 19295
rect 144736 19252 144788 19261
rect 176844 19295 176896 19304
rect 176844 19261 176853 19295
rect 176853 19261 176887 19295
rect 176887 19261 176896 19295
rect 176844 19252 176896 19261
rect 211160 19252 211212 19304
rect 212448 19295 212500 19304
rect 212448 19261 212457 19295
rect 212457 19261 212491 19295
rect 212491 19261 212500 19295
rect 212448 19252 212500 19261
rect 333888 19295 333940 19304
rect 333888 19261 333897 19295
rect 333897 19261 333931 19295
rect 333931 19261 333940 19295
rect 333888 19252 333940 19261
rect 333980 19252 334032 19304
rect 334808 19252 334860 19304
rect 338120 19295 338172 19304
rect 338120 19261 338129 19295
rect 338129 19261 338163 19295
rect 338163 19261 338172 19295
rect 389180 19295 389232 19304
rect 338120 19252 338172 19261
rect 389180 19261 389189 19295
rect 389189 19261 389223 19295
rect 389223 19261 389232 19295
rect 389180 19252 389232 19261
rect 391756 19295 391808 19304
rect 391756 19261 391765 19295
rect 391765 19261 391799 19295
rect 391799 19261 391808 19295
rect 391756 19252 391808 19261
rect 411168 19295 411220 19304
rect 411168 19261 411177 19295
rect 411177 19261 411211 19295
rect 411211 19261 411220 19295
rect 411168 19252 411220 19261
rect 414020 19252 414072 19304
rect 414480 19252 414532 19304
rect 117228 18708 117280 18760
rect 136640 18708 136692 18760
rect 364248 18708 364300 18760
rect 546592 18708 546644 18760
rect 80796 18640 80848 18692
rect 502340 18640 502392 18692
rect 37188 18572 37240 18624
rect 64144 18572 64196 18624
rect 85488 18572 85540 18624
rect 509424 18572 509476 18624
rect 547144 17960 547196 18012
rect 549260 17960 549312 18012
rect 563704 17892 563756 17944
rect 579804 17892 579856 17944
rect 231768 17348 231820 17400
rect 365720 17348 365772 17400
rect 450544 17348 450596 17400
rect 455328 17348 455380 17400
rect 125508 17280 125560 17332
rect 452660 17280 452712 17332
rect 91008 17212 91060 17264
rect 518992 17212 519044 17264
rect 202788 16056 202840 16108
rect 368480 16056 368532 16108
rect 384948 16056 385000 16108
rect 459560 16056 459612 16108
rect 115848 15988 115900 16040
rect 186320 15988 186372 16040
rect 193128 15988 193180 16040
rect 397460 15988 397512 16040
rect 59268 15920 59320 15972
rect 233240 15920 233292 15972
rect 286968 15920 287020 15972
rect 502800 15920 502852 15972
rect 39948 15852 40000 15904
rect 327724 15852 327776 15904
rect 412548 15852 412600 15904
rect 427820 15852 427872 15904
rect 448428 15852 448480 15904
rect 525800 15852 525852 15904
rect 56508 15172 56560 15224
rect 57244 15172 57296 15224
rect 288348 14968 288400 15020
rect 310520 14968 310572 15020
rect 92388 14900 92440 14952
rect 186964 14900 187016 14952
rect 204168 14900 204220 14952
rect 351920 14900 351972 14952
rect 63132 14832 63184 14884
rect 371240 14832 371292 14884
rect 375288 14832 375340 14884
rect 528652 14832 528704 14884
rect 72700 14764 72752 14816
rect 412640 14764 412692 14816
rect 158628 14696 158680 14748
rect 503720 14696 503772 14748
rect 64604 14628 64656 14680
rect 416780 14628 416832 14680
rect 73896 14560 73948 14612
rect 427820 14560 427872 14612
rect 57796 14492 57848 14544
rect 459560 14492 459612 14544
rect 10968 14424 11020 14476
rect 37924 14424 37976 14476
rect 68744 14424 68796 14476
rect 560300 14424 560352 14476
rect 345020 13812 345072 13864
rect 351184 13812 351236 13864
rect 72884 13064 72936 13116
rect 124864 13064 124916 13116
rect 126888 13064 126940 13116
rect 293960 13064 294012 13116
rect 426348 13064 426400 13116
rect 500960 13064 501012 13116
rect 488448 12452 488500 12504
rect 65708 12384 65760 12436
rect 142068 12384 142120 12436
rect 169760 12384 169812 12436
rect 170588 12384 170640 12436
rect 204260 12384 204312 12436
rect 205088 12384 205140 12436
rect 212540 12384 212592 12436
rect 213460 12384 213512 12436
rect 213920 12384 213972 12436
rect 214656 12384 214708 12436
rect 280252 12384 280304 12436
rect 281172 12384 281224 12436
rect 281540 12384 281592 12436
rect 282460 12384 282512 12436
rect 335360 12384 335412 12436
rect 335912 12384 335964 12436
rect 350632 12384 350684 12436
rect 351368 12384 351420 12436
rect 351920 12384 351972 12436
rect 352564 12384 352616 12436
rect 404360 12384 404412 12436
rect 404912 12384 404964 12436
rect 412640 12384 412692 12436
rect 413284 12384 413336 12436
rect 448520 12384 448572 12436
rect 448980 12384 449032 12436
rect 454040 12384 454092 12436
rect 454868 12384 454920 12436
rect 473360 12384 473412 12436
rect 473912 12384 473964 12436
rect 486884 12384 486936 12436
rect 487068 12384 487120 12436
rect 502340 12384 502392 12436
rect 502524 12384 502576 12436
rect 81256 12316 81308 12368
rect 229100 12316 229152 12368
rect 61936 12248 61988 12300
rect 260840 12248 260892 12300
rect 63316 12180 63368 12232
rect 269120 12180 269172 12232
rect 68468 12112 68520 12164
rect 276480 12112 276532 12164
rect 61568 12044 61620 12096
rect 372620 12044 372672 12096
rect 61660 11976 61712 12028
rect 472716 11976 472768 12028
rect 46756 11908 46808 11960
rect 465080 11908 465132 11960
rect 50988 11840 51040 11892
rect 494704 11840 494756 11892
rect 511356 11840 511408 11892
rect 571340 11840 571392 11892
rect 64512 11772 64564 11824
rect 516324 11772 516376 11824
rect 65892 11704 65944 11756
rect 529940 11704 529992 11756
rect 457444 10956 457496 11008
rect 462964 10956 463016 11008
rect 77116 10412 77168 10464
rect 253940 10412 253992 10464
rect 34428 10344 34480 10396
rect 350540 10344 350592 10396
rect 17868 10276 17920 10328
rect 437480 10276 437532 10328
rect 411168 9775 411220 9784
rect 411168 9741 411177 9775
rect 411177 9741 411211 9775
rect 411211 9741 411220 9775
rect 411168 9732 411220 9741
rect 140780 9707 140832 9716
rect 140780 9673 140789 9707
rect 140789 9673 140823 9707
rect 140823 9673 140832 9707
rect 140780 9664 140832 9673
rect 144736 9707 144788 9716
rect 144736 9673 144745 9707
rect 144745 9673 144779 9707
rect 144779 9673 144788 9707
rect 144736 9664 144788 9673
rect 176936 9664 176988 9716
rect 212448 9707 212500 9716
rect 212448 9673 212457 9707
rect 212457 9673 212491 9707
rect 212491 9673 212500 9707
rect 212448 9664 212500 9673
rect 333888 9707 333940 9716
rect 333888 9673 333897 9707
rect 333897 9673 333931 9707
rect 333931 9673 333940 9707
rect 333888 9664 333940 9673
rect 338304 9664 338356 9716
rect 389456 9664 389508 9716
rect 391848 9664 391900 9716
rect 488172 9707 488224 9716
rect 488172 9673 488181 9707
rect 488181 9673 488215 9707
rect 488215 9673 488224 9707
rect 488172 9664 488224 9673
rect 512460 9707 512512 9716
rect 512460 9673 512469 9707
rect 512469 9673 512503 9707
rect 512503 9673 512512 9707
rect 512460 9664 512512 9673
rect 61476 9596 61528 9648
rect 121828 9596 121880 9648
rect 411168 9596 411220 9648
rect 502524 9596 502576 9648
rect 64788 9528 64840 9580
rect 190828 9528 190880 9580
rect 445668 9571 445720 9580
rect 445668 9537 445677 9571
rect 445677 9537 445711 9571
rect 445711 9537 445720 9571
rect 445668 9528 445720 9537
rect 59084 9460 59136 9512
rect 206284 9460 206336 9512
rect 63408 9392 63460 9444
rect 279976 9392 280028 9444
rect 113548 9324 113600 9376
rect 336740 9324 336792 9376
rect 60464 9256 60516 9308
rect 290740 9256 290792 9308
rect 65616 9188 65668 9240
rect 244372 9188 244424 9240
rect 273168 9188 273220 9240
rect 510804 9188 510856 9240
rect 68560 9120 68612 9172
rect 308588 9120 308640 9172
rect 30196 9052 30248 9104
rect 286324 9052 286376 9104
rect 444196 9052 444248 9104
rect 518900 9052 518952 9104
rect 70032 8984 70084 9036
rect 340696 8984 340748 9036
rect 376392 8984 376444 9036
rect 512092 8984 512144 9036
rect 71228 8916 71280 8968
rect 358544 8916 358596 8968
rect 382372 8916 382424 8968
rect 521660 8916 521712 8968
rect 540244 8916 540296 8968
rect 573824 8916 573876 8968
rect 462320 8848 462372 8900
rect 465724 8848 465776 8900
rect 3424 8236 3476 8288
rect 513748 8236 513800 8288
rect 54024 7624 54076 7676
rect 299480 7624 299532 7676
rect 331220 7624 331272 7676
rect 332416 7624 332468 7676
rect 408500 7624 408552 7676
rect 409696 7624 409748 7676
rect 416780 7624 416832 7676
rect 417976 7624 418028 7676
rect 447416 7624 447468 7676
rect 449164 7624 449216 7676
rect 117136 7556 117188 7608
rect 149704 7556 149756 7608
rect 178960 7556 179012 7608
rect 443000 7556 443052 7608
rect 451280 7556 451332 7608
rect 452476 7556 452528 7608
rect 494060 7556 494112 7608
rect 495348 7556 495400 7608
rect 552756 7556 552808 7608
rect 564348 7556 564400 7608
rect 201500 7488 201552 7540
rect 202696 7488 202748 7540
rect 71136 6808 71188 6860
rect 153936 6808 153988 6860
rect 60556 6740 60608 6792
rect 159916 6740 159968 6792
rect 72424 6672 72476 6724
rect 183744 6672 183796 6724
rect 475108 6672 475160 6724
rect 481088 6672 481140 6724
rect 515220 6672 515272 6724
rect 68928 6604 68980 6656
rect 125416 6604 125468 6656
rect 138480 6604 138532 6656
rect 256700 6604 256752 6656
rect 406108 6604 406160 6656
rect 434720 6604 434772 6656
rect 459652 6604 459704 6656
rect 510620 6604 510672 6656
rect 70676 6536 70728 6588
rect 225604 6536 225656 6588
rect 229008 6536 229060 6588
rect 416872 6536 416924 6588
rect 447784 6536 447836 6588
rect 514760 6536 514812 6588
rect 67364 6468 67416 6520
rect 258632 6468 258684 6520
rect 263508 6468 263560 6520
rect 313372 6468 313424 6520
rect 423956 6468 424008 6520
rect 513564 6468 513616 6520
rect 67548 6400 67600 6452
rect 318064 6400 318116 6452
rect 422760 6400 422812 6452
rect 516232 6400 516284 6452
rect 531964 6400 532016 6452
rect 572628 6400 572680 6452
rect 73988 6332 74040 6384
rect 554872 6332 554924 6384
rect 66076 6264 66128 6316
rect 558368 6264 558420 6316
rect 65984 6196 66036 6248
rect 561956 6196 562008 6248
rect 11244 6128 11296 6180
rect 19984 6128 20036 6180
rect 38476 6128 38528 6180
rect 46204 6128 46256 6180
rect 66904 6128 66956 6180
rect 569040 6128 569092 6180
rect 432328 5992 432380 6044
rect 433248 5992 433300 6044
rect 201592 5924 201644 5976
rect 211068 5924 211120 5976
rect 481824 5924 481876 5976
rect 491208 5924 491260 5976
rect 259828 5856 259880 5908
rect 260748 5856 260800 5908
rect 135260 5720 135312 5772
rect 144828 5720 144880 5772
rect 438124 5720 438176 5772
rect 442908 5720 442960 5772
rect 182180 5652 182232 5704
rect 199936 5652 199988 5704
rect 46940 5516 46992 5568
rect 50344 5516 50396 5568
rect 571984 5516 572036 5568
rect 576216 5516 576268 5568
rect 320088 5108 320140 5160
rect 350264 5040 350316 5092
rect 378692 5040 378744 5092
rect 462228 5040 462280 5092
rect 327632 4972 327684 5024
rect 457444 4972 457496 5024
rect 291936 4904 291988 4956
rect 447416 4904 447468 4956
rect 456708 4904 456760 4956
rect 467932 4904 467984 4956
rect 206928 4836 206980 4888
rect 225328 4836 225380 4888
rect 287152 4836 287204 4888
rect 450544 4836 450596 4888
rect 6460 4768 6512 4820
rect 14464 4768 14516 4820
rect 40960 4768 41012 4820
rect 55864 4768 55916 4820
rect 112352 4768 112404 4820
rect 237380 4768 237432 4820
rect 272892 4768 272944 4820
rect 460204 4768 460256 4820
rect 527824 4768 527876 4820
rect 548892 4768 548944 4820
rect 554044 4768 554096 4820
rect 578608 4768 578660 4820
rect 502432 4632 502484 4684
rect 503628 4632 503680 4684
rect 12440 4360 12492 4412
rect 17224 4360 17276 4412
rect 133696 4156 133748 4208
rect 64420 4088 64472 4140
rect 133788 4088 133840 4140
rect 572 4020 624 4072
rect 9036 4020 9088 4072
rect 64328 4020 64380 4072
rect 80244 4020 80296 4072
rect 84844 4020 84896 4072
rect 142160 4020 142212 4072
rect 143264 4020 143316 4072
rect 145656 4020 145708 4072
rect 146208 4020 146260 4072
rect 146300 4020 146352 4072
rect 146852 4020 146904 4072
rect 157524 4020 157576 4072
rect 158628 4020 158680 4072
rect 167000 4020 167052 4072
rect 168196 4020 168248 4072
rect 176936 4020 176988 4072
rect 177764 4020 177816 4072
rect 179420 4020 179472 4072
rect 180156 4020 180208 4072
rect 198004 4020 198056 4072
rect 198648 4020 198700 4072
rect 199200 4020 199252 4072
rect 200028 4020 200080 4072
rect 201500 4020 201552 4072
rect 202788 4020 202840 4072
rect 207020 4020 207072 4072
rect 207480 4020 207532 4072
rect 208676 4020 208728 4072
rect 209688 4020 209740 4072
rect 209872 4020 209924 4072
rect 210884 4020 210936 4072
rect 217048 4020 217100 4072
rect 217968 4020 218020 4072
rect 218060 4020 218112 4072
rect 219348 4020 219400 4072
rect 274088 4020 274140 4072
rect 274548 4020 274600 4072
rect 275284 4020 275336 4072
rect 275928 4020 275980 4072
rect 278872 4020 278924 4072
rect 280068 4020 280120 4072
rect 331220 4020 331272 4072
rect 332508 4020 332560 4072
rect 337108 4020 337160 4072
rect 338028 4020 338080 4072
rect 356152 4020 356204 4072
rect 357348 4020 357400 4072
rect 397828 4020 397880 4072
rect 398748 4020 398800 4072
rect 399024 4020 399076 4072
rect 400128 4020 400180 4072
rect 408500 4020 408552 4072
rect 409788 4020 409840 4072
rect 412088 4020 412140 4072
rect 412548 4020 412600 4072
rect 456064 4020 456116 4072
rect 456616 4020 456668 4072
rect 466828 4020 466880 4072
rect 467748 4020 467800 4072
rect 485780 4020 485832 4072
rect 486976 4020 487028 4072
rect 498936 4020 498988 4072
rect 499488 4020 499540 4072
rect 511448 4088 511500 4140
rect 513196 4088 513248 4140
rect 512184 4020 512236 4072
rect 69940 3952 69992 4004
rect 150440 3952 150492 4004
rect 470324 3952 470376 4004
rect 494152 3952 494204 4004
rect 497740 3952 497792 4004
rect 517704 3952 517756 4004
rect 68652 3884 68704 3936
rect 162308 3884 162360 3936
rect 477500 3884 477552 3936
rect 500132 3884 500184 3936
rect 500868 3884 500920 3936
rect 513472 3884 513524 3936
rect 64696 3816 64748 3868
rect 165896 3816 165948 3868
rect 60372 3748 60424 3800
rect 167092 3748 167144 3800
rect 66996 3680 67048 3732
rect 74448 3680 74500 3732
rect 257436 3816 257488 3868
rect 375288 3816 375340 3868
rect 406384 3816 406436 3868
rect 431132 3816 431184 3868
rect 439504 3816 439556 3868
rect 443000 3816 443052 3868
rect 502984 3816 503036 3868
rect 300308 3748 300360 3800
rect 378692 3748 378744 3800
rect 401324 3748 401376 3800
rect 512368 3748 512420 3800
rect 270500 3680 270552 3732
rect 513380 3680 513432 3732
rect 63224 3612 63276 3664
rect 222936 3612 222988 3664
rect 227720 3612 227772 3664
rect 228916 3612 228968 3664
rect 236000 3612 236052 3664
rect 237196 3612 237248 3664
rect 252652 3612 252704 3664
rect 253848 3612 253900 3664
rect 520372 3612 520424 3664
rect 7656 3544 7708 3596
rect 15844 3544 15896 3596
rect 20720 3544 20772 3596
rect 21916 3544 21968 3596
rect 29092 3544 29144 3596
rect 30288 3544 30340 3596
rect 43352 3544 43404 3596
rect 315304 3544 315356 3596
rect 321652 3544 321704 3596
rect 322848 3544 322900 3596
rect 322940 3544 322992 3596
rect 517612 3544 517664 3596
rect 520280 3544 520332 3596
rect 521476 3544 521528 3596
rect 574744 3544 574796 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 17224 3476 17276 3528
rect 17868 3476 17920 3528
rect 18328 3476 18380 3528
rect 19248 3476 19300 3528
rect 19524 3476 19576 3528
rect 20628 3476 20680 3528
rect 25504 3476 25556 3528
rect 26148 3476 26200 3528
rect 26700 3476 26752 3528
rect 27528 3476 27580 3528
rect 27896 3476 27948 3528
rect 28908 3476 28960 3528
rect 33876 3476 33928 3528
rect 34428 3476 34480 3528
rect 34980 3476 35032 3528
rect 35808 3476 35860 3528
rect 36176 3476 36228 3528
rect 37188 3476 37240 3528
rect 37372 3476 37424 3528
rect 38568 3476 38620 3528
rect 42156 3476 42208 3528
rect 42708 3476 42760 3528
rect 44548 3476 44600 3528
rect 45468 3476 45520 3528
rect 45744 3476 45796 3528
rect 46756 3476 46808 3528
rect 51632 3476 51684 3528
rect 52368 3476 52420 3528
rect 52828 3476 52880 3528
rect 53748 3476 53800 3528
rect 60004 3476 60056 3528
rect 60648 3476 60700 3528
rect 61200 3476 61252 3528
rect 62028 3476 62080 3528
rect 62396 3476 62448 3528
rect 63040 3476 63092 3528
rect 63592 3476 63644 3528
rect 64236 3476 64288 3528
rect 68284 3476 68336 3528
rect 68836 3476 68888 3528
rect 71872 3476 71924 3528
rect 72884 3476 72936 3528
rect 2872 3408 2924 3460
rect 13084 3408 13136 3460
rect 58808 3408 58860 3460
rect 59268 3408 59320 3460
rect 72792 3408 72844 3460
rect 515588 3476 515640 3528
rect 518164 3476 518216 3528
rect 542912 3476 542964 3528
rect 554780 3476 554832 3528
rect 555976 3476 556028 3528
rect 581000 3476 581052 3528
rect 522672 3408 522724 3460
rect 528560 3408 528612 3460
rect 529848 3408 529900 3460
rect 573364 3408 573416 3460
rect 579804 3408 579856 3460
rect 76656 3340 76708 3392
rect 77208 3340 77260 3392
rect 77852 3340 77904 3392
rect 78312 3340 78364 3392
rect 81900 3340 81952 3392
rect 82636 3340 82688 3392
rect 87328 3340 87380 3392
rect 88248 3340 88300 3392
rect 89720 3340 89772 3392
rect 90916 3340 90968 3392
rect 93308 3340 93360 3392
rect 93768 3340 93820 3392
rect 93952 3340 94004 3392
rect 94504 3340 94556 3392
rect 95700 3340 95752 3392
rect 96528 3340 96580 3392
rect 96896 3340 96948 3392
rect 97908 3340 97960 3392
rect 98092 3340 98144 3392
rect 99380 3340 99432 3392
rect 101588 3340 101640 3392
rect 102048 3340 102100 3392
rect 102784 3340 102836 3392
rect 103428 3340 103480 3392
rect 105176 3340 105228 3392
rect 106188 3340 106240 3392
rect 106372 3340 106424 3392
rect 107660 3340 107712 3392
rect 114744 3340 114796 3392
rect 115756 3340 115808 3392
rect 117320 3340 117372 3392
rect 118240 3340 118292 3392
rect 119436 3340 119488 3392
rect 119988 3340 120040 3392
rect 124220 3340 124272 3392
rect 125508 3340 125560 3392
rect 127808 3340 127860 3392
rect 128268 3340 128320 3392
rect 129740 3340 129792 3392
rect 130200 3340 130252 3392
rect 136088 3340 136140 3392
rect 136548 3340 136600 3392
rect 148048 3340 148100 3392
rect 148968 3340 149020 3392
rect 158720 3340 158772 3392
rect 187792 3340 187844 3392
rect 188436 3340 188488 3392
rect 189632 3340 189684 3392
rect 190368 3340 190420 3392
rect 192024 3340 192076 3392
rect 193128 3340 193180 3392
rect 226524 3340 226576 3392
rect 227628 3340 227680 3392
rect 232504 3340 232556 3392
rect 233148 3340 233200 3392
rect 239588 3340 239640 3392
rect 240048 3340 240100 3392
rect 240784 3340 240836 3392
rect 241428 3340 241480 3392
rect 249156 3340 249208 3392
rect 249708 3340 249760 3392
rect 250352 3340 250404 3392
rect 251088 3340 251140 3392
rect 251456 3340 251508 3392
rect 262220 3340 262272 3392
rect 263416 3340 263468 3392
rect 283656 3340 283708 3392
rect 284208 3340 284260 3392
rect 285956 3340 286008 3392
rect 286968 3340 287020 3392
rect 287060 3340 287112 3392
rect 288348 3340 288400 3392
rect 293132 3340 293184 3392
rect 293868 3340 293920 3392
rect 296720 3340 296772 3392
rect 298008 3340 298060 3392
rect 301412 3340 301464 3392
rect 302148 3340 302200 3392
rect 303804 3340 303856 3392
rect 304908 3340 304960 3392
rect 305000 3340 305052 3392
rect 306196 3340 306248 3392
rect 326436 3340 326488 3392
rect 326988 3340 327040 3392
rect 330024 3340 330076 3392
rect 331128 3340 331180 3392
rect 344284 3340 344336 3392
rect 344928 3340 344980 3392
rect 361580 3340 361632 3392
rect 362132 3340 362184 3392
rect 363328 3340 363380 3392
rect 364156 3340 364208 3392
rect 364524 3340 364576 3392
rect 365628 3340 365680 3392
rect 365720 3340 365772 3392
rect 366916 3340 366968 3392
rect 370412 3340 370464 3392
rect 371148 3340 371200 3392
rect 374000 3340 374052 3392
rect 375196 3340 375248 3392
rect 379980 3340 380032 3392
rect 380808 3340 380860 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 385868 3340 385920 3392
rect 386328 3340 386380 3392
rect 388260 3340 388312 3392
rect 389088 3340 389140 3392
rect 421564 3340 421616 3392
rect 422208 3340 422260 3392
rect 425060 3340 425112 3392
rect 426348 3340 426400 3392
rect 433340 3340 433392 3392
rect 434628 3340 434680 3392
rect 439412 3340 439464 3392
rect 440148 3340 440200 3392
rect 459560 3340 459612 3392
rect 460848 3340 460900 3392
rect 483480 3340 483532 3392
rect 484308 3340 484360 3392
rect 507860 3340 507912 3392
rect 155132 3272 155184 3324
rect 155868 3272 155920 3324
rect 175372 3272 175424 3324
rect 176568 3272 176620 3324
rect 182548 3272 182600 3324
rect 183468 3272 183520 3324
rect 241980 3272 242032 3324
rect 242808 3272 242860 3324
rect 339500 3272 339552 3324
rect 340788 3272 340840 3324
rect 494152 3272 494204 3324
rect 543004 3272 543056 3324
rect 546500 3272 546552 3324
rect 89996 3204 90048 3256
rect 90916 3204 90968 3256
rect 218152 3204 218204 3256
rect 219256 3204 219308 3256
rect 277676 3204 277728 3256
rect 278688 3204 278740 3256
rect 305000 3204 305052 3256
rect 306288 3204 306340 3256
rect 365720 3204 365772 3256
rect 367008 3204 367060 3256
rect 200396 3136 200448 3188
rect 201408 3136 201460 3188
rect 215852 3136 215904 3188
rect 216588 3136 216640 3188
rect 328828 3136 328880 3188
rect 329748 3136 329800 3188
rect 353760 3136 353812 3188
rect 354588 3136 354640 3188
rect 354956 3136 355008 3188
rect 355968 3136 356020 3188
rect 172980 3068 173032 3120
rect 173808 3068 173860 3120
rect 415676 3068 415728 3120
rect 416688 3068 416740 3120
rect 84936 3000 84988 3052
rect 85488 3000 85540 3052
rect 163504 3000 163556 3052
rect 164148 3000 164200 3052
rect 164700 3000 164752 3052
rect 165528 3000 165580 3052
rect 319260 3000 319312 3052
rect 319996 3000 320048 3052
rect 347872 3000 347924 3052
rect 349068 3000 349120 3052
rect 504364 3000 504416 3052
rect 507216 3000 507268 3052
rect 181352 2932 181404 2984
rect 182088 2932 182140 2984
rect 4068 2864 4120 2916
rect 8944 2864 8996 2916
rect 50528 2864 50580 2916
rect 50988 2864 51040 2916
rect 69480 2864 69532 2916
rect 70124 2864 70176 2916
rect 139676 2864 139728 2916
rect 140688 2864 140740 2916
rect 144736 2796 144788 2848
rect 161112 2796 161164 2848
rect 161388 2796 161440 2848
rect 204076 2796 204128 2848
rect 212448 2796 212500 2848
rect 333888 2796 333940 2848
rect 393228 2796 393280 2848
rect 453672 2796 453724 2848
rect 453948 2796 454000 2848
rect 144460 2728 144512 2780
rect 212264 2728 212316 2780
rect 333612 2728 333664 2780
rect 512000 2728 512052 2780
rect 512552 2728 512604 2780
rect 536840 2320 536892 2372
rect 538128 2320 538180 2372
rect 445760 2184 445812 2236
rect 446588 2184 446640 2236
rect 99472 552 99524 604
rect 100484 552 100536 604
rect 120080 552 120132 604
rect 120632 552 120684 604
rect 128360 552 128412 604
rect 129004 552 129056 604
rect 171140 552 171192 604
rect 171784 552 171836 604
rect 186320 552 186372 604
rect 187240 552 187292 604
rect 195980 552 196032 604
rect 196808 552 196860 604
rect 203892 595 203944 604
rect 203892 561 203901 595
rect 203901 561 203935 595
rect 203935 561 203944 595
rect 203892 552 203944 561
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 223580 552 223632 604
rect 224132 552 224184 604
rect 247960 552 248012 604
rect 248328 552 248380 604
rect 358820 552 358872 604
rect 359740 552 359792 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 393044 595 393096 604
rect 393044 561 393053 595
rect 393053 561 393087 595
rect 393087 561 393096 595
rect 393044 552 393096 561
rect 393320 552 393372 604
rect 394240 552 394292 604
rect 396080 552 396132 604
rect 396632 552 396684 604
rect 401600 552 401652 604
rect 402520 552 402572 604
rect 410892 595 410944 604
rect 410892 561 410901 595
rect 410901 561 410935 595
rect 410935 561 410944 595
rect 410892 552 410944 561
rect 492680 552 492732 604
rect 492956 552 493008 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 500960 552 501012 604
rect 501236 552 501288 604
rect 502432 595 502484 604
rect 502432 561 502441 595
rect 502441 561 502475 595
rect 502475 561 502484 595
rect 502432 552 502484 561
rect 505100 552 505152 604
rect 506020 552 506072 604
rect 508136 552 508188 604
rect 508412 552 508464 604
rect 513656 552 513708 604
rect 514392 552 514444 604
rect 576860 552 576912 604
rect 577412 552 577464 604
rect 581092 552 581144 604
rect 582196 552 582248 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700262 8156 703520
rect 8116 700256 8168 700262
rect 8116 700198 8168 700204
rect 14464 700256 14516 700262
rect 14464 700198 14516 700204
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 8944 602540 8996 602546
rect 8944 602482 8996 602488
rect 2688 599276 2740 599282
rect 2688 599218 2740 599224
rect 572 4072 624 4078
rect 572 4014 624 4020
rect 584 480 612 4014
rect 2700 3534 2728 599218
rect 2870 596048 2926 596057
rect 2870 595983 2926 595992
rect 2884 594862 2912 595983
rect 2872 594856 2924 594862
rect 2872 594798 2924 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 538286 3464 538591
rect 3424 538280 3476 538286
rect 3424 538222 3476 538228
rect 3146 509960 3202 509969
rect 3146 509895 3202 509904
rect 3160 509318 3188 509895
rect 3148 509312 3200 509318
rect 3148 509254 3200 509260
rect 3424 496800 3476 496806
rect 3424 496742 3476 496748
rect 3436 495553 3464 496742
rect 3422 495544 3478 495553
rect 3422 495479 3478 495488
rect 3792 481636 3844 481642
rect 3792 481578 3844 481584
rect 3804 481137 3832 481578
rect 3790 481128 3846 481137
rect 3790 481063 3846 481072
rect 3422 438016 3478 438025
rect 3422 437951 3478 437960
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 3436 417450 3464 437951
rect 3424 417444 3476 417450
rect 3424 417386 3476 417392
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3344 394738 3372 394975
rect 3332 394732 3384 394738
rect 3332 394674 3384 394680
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3436 379574 3464 380559
rect 3424 379568 3476 379574
rect 3424 379510 3476 379516
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3436 336802 3464 337447
rect 3424 336796 3476 336802
rect 3424 336738 3476 336744
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 3424 308984 3476 308990
rect 3424 308926 3476 308932
rect 3436 308825 3464 308926
rect 3422 308816 3478 308825
rect 3422 308751 3478 308760
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 278905 3464 280055
rect 3422 278896 3478 278905
rect 3422 278831 3478 278840
rect 3422 265704 3478 265713
rect 3422 265639 3478 265648
rect 3436 264994 3464 265639
rect 3424 264988 3476 264994
rect 3424 264930 3476 264936
rect 3422 251288 3478 251297
rect 3422 251223 3424 251232
rect 3476 251223 3478 251232
rect 3424 251194 3476 251200
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3514 136368 3570 136377
rect 3514 136303 3570 136312
rect 3528 135862 3556 136303
rect 3516 135856 3568 135862
rect 3516 135798 3568 135804
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3436 121514 3464 122023
rect 3424 121508 3476 121514
rect 3424 121450 3476 121456
rect 4068 107704 4120 107710
rect 4066 107672 4068 107681
rect 4120 107672 4122 107681
rect 4066 107607 4122 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3422 80064 3478 80073
rect 3422 79999 3478 80008
rect 3436 78985 3464 79999
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 480 4108 2858
rect 5262 2816 5318 2825
rect 5262 2751 5318 2760
rect 5276 480 5304 2751
rect 6472 480 6500 4762
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 480 7696 3538
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 480 8892 3470
rect 8956 2922 8984 602482
rect 9036 602132 9088 602138
rect 9036 602074 9088 602080
rect 9048 4078 9076 602074
rect 13082 600536 13138 600545
rect 13082 600471 13138 600480
rect 9128 509312 9180 509318
rect 9128 509254 9180 509260
rect 9140 322930 9168 509254
rect 9128 322924 9180 322930
rect 9128 322866 9180 322872
rect 9128 317484 9180 317490
rect 9128 317426 9180 317432
rect 9140 308990 9168 317426
rect 9128 308984 9180 308990
rect 9128 308926 9180 308932
rect 9128 135856 9180 135862
rect 9128 135798 9180 135804
rect 9140 102746 9168 135798
rect 11704 121508 11756 121514
rect 11704 121450 11756 121456
rect 9128 102740 9180 102746
rect 9128 102682 9180 102688
rect 11716 100706 11744 121450
rect 11704 100700 11756 100706
rect 11704 100642 11756 100648
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9600 3534 9628 29718
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10980 3534 11008 14418
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 10060 480 10088 3470
rect 11256 480 11284 6122
rect 12440 4412 12492 4418
rect 12440 4354 12492 4360
rect 12452 480 12480 4354
rect 13096 3466 13124 600471
rect 13176 379568 13228 379574
rect 13176 379510 13228 379516
rect 13188 351898 13216 379510
rect 13176 351892 13228 351898
rect 13176 351834 13228 351840
rect 14476 158710 14504 700198
rect 24320 699718 24348 703520
rect 40512 699718 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 70308 700664 70360 700670
rect 70308 700606 70360 700612
rect 67456 700392 67508 700398
rect 67456 700334 67508 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 40500 699712 40552 699718
rect 40500 699654 40552 699660
rect 43444 699712 43496 699718
rect 43444 699654 43496 699660
rect 17224 652792 17276 652798
rect 17224 652734 17276 652740
rect 15844 600364 15896 600370
rect 15844 600306 15896 600312
rect 14464 158704 14516 158710
rect 14464 158646 14516 158652
rect 14464 149116 14516 149122
rect 14464 149058 14516 149064
rect 13634 30968 13690 30977
rect 13634 30903 13690 30912
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 13648 480 13676 30903
rect 14476 4826 14504 149058
rect 15108 55888 15160 55894
rect 15108 55830 15160 55836
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 15120 3482 15148 55830
rect 15856 3602 15884 600306
rect 15936 346452 15988 346458
rect 15936 346394 15988 346400
rect 15948 93838 15976 346394
rect 17236 329798 17264 652734
rect 21364 604852 21416 604858
rect 21364 604794 21416 604800
rect 20076 594108 20128 594114
rect 20076 594050 20128 594056
rect 19984 427848 20036 427854
rect 19984 427790 20036 427796
rect 17224 329792 17276 329798
rect 17224 329734 17276 329740
rect 17224 146328 17276 146334
rect 17224 146270 17276 146276
rect 15936 93832 15988 93838
rect 15936 93774 15988 93780
rect 16026 8936 16082 8945
rect 16026 8871 16082 8880
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 14844 3454 15148 3482
rect 14844 480 14872 3454
rect 16040 480 16068 8871
rect 17236 4418 17264 146270
rect 19248 73840 19300 73846
rect 19248 73782 19300 73788
rect 17868 10328 17920 10334
rect 17868 10270 17920 10276
rect 17224 4412 17276 4418
rect 17224 4354 17276 4360
rect 17880 3534 17908 10270
rect 19260 3534 19288 73782
rect 19996 6186 20024 427790
rect 20088 180810 20116 594050
rect 21376 295322 21404 604794
rect 24674 600672 24730 600681
rect 24674 600607 24730 600616
rect 21364 295316 21416 295322
rect 21364 295258 21416 295264
rect 20076 180804 20128 180810
rect 20076 180746 20128 180752
rect 22008 62892 22060 62898
rect 22008 62834 22060 62840
rect 20628 25560 20680 25566
rect 20628 25502 20680 25508
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 20640 3534 20668 25502
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21928 3602 21956 19926
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 17236 480 17264 3470
rect 18340 480 18368 3470
rect 19536 480 19564 3470
rect 20732 480 20760 3538
rect 22020 3482 22048 62834
rect 23110 3768 23166 3777
rect 23110 3703 23166 3712
rect 21928 3454 22048 3482
rect 21928 480 21956 3454
rect 23124 480 23152 3703
rect 24688 3482 24716 600607
rect 24780 102105 24808 699654
rect 43456 616146 43484 699654
rect 55864 623824 55916 623830
rect 55864 623766 55916 623772
rect 43444 616140 43496 616146
rect 43444 616082 43496 616088
rect 48964 610020 49016 610026
rect 48964 609962 49016 609968
rect 39396 605872 39448 605878
rect 39396 605814 39448 605820
rect 28264 603220 28316 603226
rect 28264 603162 28316 603168
rect 27528 601996 27580 602002
rect 27528 601938 27580 601944
rect 25504 567248 25556 567254
rect 25504 567190 25556 567196
rect 24766 102096 24822 102105
rect 24766 102031 24822 102040
rect 25516 97986 25544 567190
rect 25504 97980 25556 97986
rect 25504 97922 25556 97928
rect 26148 23180 26200 23186
rect 26148 23122 26200 23128
rect 26160 3534 26188 23122
rect 27540 3534 27568 601938
rect 28276 23186 28304 603162
rect 31668 602676 31720 602682
rect 31668 602618 31720 602624
rect 30288 596828 30340 596834
rect 30288 596770 30340 596776
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28908 22840 28960 22846
rect 28908 22782 28960 22788
rect 28920 3534 28948 22782
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 24320 3454 24716 3482
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 24320 480 24348 3454
rect 25516 480 25544 3470
rect 26712 480 26740 3470
rect 27908 480 27936 3470
rect 29104 480 29132 3538
rect 30208 3482 30236 9046
rect 30300 3602 30328 596770
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 31680 3482 31708 602618
rect 35806 595504 35862 595513
rect 35806 595439 35862 595448
rect 32404 594856 32456 594862
rect 32404 594798 32456 594804
rect 32416 96558 32444 594798
rect 33784 397520 33836 397526
rect 33784 397462 33836 397468
rect 32404 96552 32456 96558
rect 32404 96494 32456 96500
rect 33796 64870 33824 397462
rect 33784 64864 33836 64870
rect 33784 64806 33836 64812
rect 33046 24168 33102 24177
rect 33046 24103 33102 24112
rect 33060 3482 33088 24103
rect 34428 10396 34480 10402
rect 34428 10338 34480 10344
rect 34440 3534 34468 10338
rect 35820 3534 35848 595439
rect 39304 552084 39356 552090
rect 39304 552026 39356 552032
rect 37924 361616 37976 361622
rect 37924 361558 37976 361564
rect 37188 18624 37240 18630
rect 37188 18566 37240 18572
rect 37200 3534 37228 18566
rect 37936 14482 37964 361558
rect 39316 100842 39344 552026
rect 39408 481642 39436 605814
rect 48226 601896 48282 601905
rect 48226 601831 48282 601840
rect 42708 592680 42760 592686
rect 42708 592622 42760 592628
rect 39396 481636 39448 481642
rect 39396 481578 39448 481584
rect 39304 100836 39356 100842
rect 39304 100778 39356 100784
rect 38568 26988 38620 26994
rect 38568 26930 38620 26936
rect 37924 14476 37976 14482
rect 37924 14418 37976 14424
rect 38476 6180 38528 6186
rect 38476 6122 38528 6128
rect 30208 3454 30328 3482
rect 30300 480 30328 3454
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34980 3528 35032 3534
rect 34980 3470 35032 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 33888 480 33916 3470
rect 34992 480 35020 3470
rect 36188 480 36216 3470
rect 37384 480 37412 3470
rect 38488 3074 38516 6122
rect 38580 3534 38608 26930
rect 39948 15904 40000 15910
rect 39948 15846 40000 15852
rect 38568 3528 38620 3534
rect 39960 3482 39988 15846
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 38568 3470 38620 3476
rect 39776 3454 39988 3482
rect 38488 3046 38608 3074
rect 38580 480 38608 3046
rect 39776 480 39804 3454
rect 40972 480 41000 4762
rect 42720 3534 42748 592622
rect 46848 565888 46900 565894
rect 46848 565830 46900 565836
rect 43444 538280 43496 538286
rect 43444 538222 43496 538228
rect 43456 97918 43484 538222
rect 46204 419552 46256 419558
rect 46204 419494 46256 419500
rect 43444 97912 43496 97918
rect 43444 97854 43496 97860
rect 45468 60104 45520 60110
rect 45468 60046 45520 60052
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42168 480 42196 3470
rect 43364 480 43392 3538
rect 45480 3534 45508 60046
rect 46216 6186 46244 419494
rect 46756 11960 46808 11966
rect 46756 11902 46808 11908
rect 46204 6180 46256 6186
rect 46204 6122 46256 6128
rect 46768 3534 46796 11902
rect 46860 9081 46888 565830
rect 46846 9072 46902 9081
rect 46846 9007 46902 9016
rect 46940 5568 46992 5574
rect 46940 5510 46992 5516
rect 44548 3528 44600 3534
rect 44548 3470 44600 3476
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 44560 480 44588 3470
rect 45756 480 45784 3470
rect 46952 480 46980 5510
rect 48240 3482 48268 601831
rect 48976 471986 49004 609962
rect 52366 601760 52422 601769
rect 52366 601695 52422 601704
rect 50344 569968 50396 569974
rect 50344 569910 50396 569916
rect 48964 471980 49016 471986
rect 48964 471922 49016 471928
rect 49608 368552 49660 368558
rect 49608 368494 49660 368500
rect 49620 3482 49648 368494
rect 50356 5574 50384 569910
rect 50988 11892 51040 11898
rect 50988 11834 51040 11840
rect 50344 5568 50396 5574
rect 50344 5510 50396 5516
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 51000 2922 51028 11834
rect 52380 3534 52408 601695
rect 53746 600400 53802 600409
rect 53746 600335 53802 600344
rect 53760 3534 53788 600335
rect 55876 263566 55904 623766
rect 57888 608660 57940 608666
rect 57888 608602 57940 608608
rect 57244 604920 57296 604926
rect 57244 604862 57296 604868
rect 56508 603560 56560 603566
rect 56508 603502 56560 603508
rect 55864 263560 55916 263566
rect 55864 263502 55916 263508
rect 55864 233300 55916 233306
rect 55864 233242 55916 233248
rect 54024 7676 54076 7682
rect 54024 7618 54076 7624
rect 51632 3528 51684 3534
rect 51632 3470 51684 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52828 3528 52880 3534
rect 52828 3470 52880 3476
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 50528 2916 50580 2922
rect 50528 2858 50580 2864
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50540 480 50568 2858
rect 51644 480 51672 3470
rect 52840 480 52868 3470
rect 54036 480 54064 7618
rect 55218 4856 55274 4865
rect 55876 4826 55904 233242
rect 56520 101726 56548 603502
rect 57256 208350 57284 604862
rect 57796 335368 57848 335374
rect 57796 335310 57848 335316
rect 57704 266416 57756 266422
rect 57704 266358 57756 266364
rect 57244 208344 57296 208350
rect 57244 208286 57296 208292
rect 57244 131164 57296 131170
rect 57244 131106 57296 131112
rect 56508 101720 56560 101726
rect 56508 101662 56560 101668
rect 57256 15230 57284 131106
rect 56508 15224 56560 15230
rect 56508 15166 56560 15172
rect 57244 15224 57296 15230
rect 57244 15166 57296 15172
rect 55218 4791 55274 4800
rect 55864 4820 55916 4826
rect 55232 480 55260 4791
rect 55864 4762 55916 4768
rect 56520 626 56548 15166
rect 57716 626 57744 266358
rect 57808 14550 57836 335310
rect 57900 97374 57928 608602
rect 64788 607300 64840 607306
rect 64788 607242 64840 607248
rect 61844 606484 61896 606490
rect 61844 606426 61896 606432
rect 61752 606416 61804 606422
rect 61752 606358 61804 606364
rect 60556 603152 60608 603158
rect 60556 603094 60608 603100
rect 59268 602472 59320 602478
rect 59268 602414 59320 602420
rect 59174 601080 59230 601089
rect 59174 601015 59230 601024
rect 59084 430636 59136 430642
rect 59084 430578 59136 430584
rect 57888 97368 57940 97374
rect 57888 97310 57940 97316
rect 57796 14544 57848 14550
rect 57796 14486 57848 14492
rect 59096 9518 59124 430578
rect 59188 101697 59216 601015
rect 59174 101688 59230 101697
rect 59174 101623 59230 101632
rect 59280 93158 59308 602414
rect 60464 592068 60516 592074
rect 60464 592010 60516 592016
rect 60372 445800 60424 445806
rect 60372 445742 60424 445748
rect 59268 93152 59320 93158
rect 59268 93094 59320 93100
rect 59268 15972 59320 15978
rect 59268 15914 59320 15920
rect 59084 9512 59136 9518
rect 59084 9454 59136 9460
rect 59280 3466 59308 15914
rect 60384 3806 60412 445742
rect 60476 9314 60504 592010
rect 60464 9308 60516 9314
rect 60464 9250 60516 9256
rect 60568 6798 60596 603094
rect 60646 602304 60702 602313
rect 60646 602239 60702 602248
rect 60556 6792 60608 6798
rect 60556 6734 60608 6740
rect 60372 3800 60424 3806
rect 60372 3742 60424 3748
rect 60660 3534 60688 602239
rect 61660 496868 61712 496874
rect 61660 496810 61712 496816
rect 61568 478916 61620 478922
rect 61568 478858 61620 478864
rect 61476 229152 61528 229158
rect 61476 229094 61528 229100
rect 61488 9654 61516 229094
rect 61580 12102 61608 478858
rect 61568 12096 61620 12102
rect 61568 12038 61620 12044
rect 61672 12034 61700 496810
rect 61764 98870 61792 606358
rect 61752 98864 61804 98870
rect 61752 98806 61804 98812
rect 61856 97442 61884 606426
rect 64604 603900 64656 603906
rect 64604 603842 64656 603848
rect 64144 603356 64196 603362
rect 64144 603298 64196 603304
rect 62028 600568 62080 600574
rect 62028 600510 62080 600516
rect 61936 600432 61988 600438
rect 61936 600374 61988 600380
rect 61844 97436 61896 97442
rect 61844 97378 61896 97384
rect 61948 12306 61976 600374
rect 61936 12300 61988 12306
rect 61936 12242 61988 12248
rect 61660 12028 61712 12034
rect 61660 11970 61712 11976
rect 61476 9648 61528 9654
rect 61476 9590 61528 9596
rect 62040 3534 62068 600510
rect 63408 554804 63460 554810
rect 63408 554746 63460 554752
rect 63316 510672 63368 510678
rect 63316 510614 63368 510620
rect 63224 405748 63276 405754
rect 63224 405690 63276 405696
rect 63132 386436 63184 386442
rect 63132 386378 63184 386384
rect 63040 332648 63092 332654
rect 63040 332590 63092 332596
rect 63052 3534 63080 332590
rect 63144 14890 63172 386378
rect 63132 14884 63184 14890
rect 63132 14826 63184 14832
rect 63236 3670 63264 405690
rect 63328 12238 63356 510614
rect 63316 12232 63368 12238
rect 63316 12174 63368 12180
rect 63420 9450 63448 554746
rect 64156 18630 64184 603298
rect 64512 507884 64564 507890
rect 64512 507826 64564 507832
rect 64420 441652 64472 441658
rect 64420 441594 64472 441600
rect 64328 401668 64380 401674
rect 64328 401610 64380 401616
rect 64234 39264 64290 39273
rect 64234 39199 64290 39208
rect 64144 18624 64196 18630
rect 64144 18566 64196 18572
rect 63408 9444 63460 9450
rect 63408 9386 63460 9392
rect 63224 3664 63276 3670
rect 63224 3606 63276 3612
rect 64248 3534 64276 39199
rect 64340 4078 64368 401610
rect 64432 4146 64460 441594
rect 64524 11830 64552 507826
rect 64616 14686 64644 603842
rect 64696 599004 64748 599010
rect 64696 598946 64748 598952
rect 64604 14680 64656 14686
rect 64604 14622 64656 14628
rect 64512 11824 64564 11830
rect 64512 11766 64564 11772
rect 64602 11656 64658 11665
rect 64602 11591 64658 11600
rect 64420 4140 64472 4146
rect 64420 4082 64472 4088
rect 64328 4072 64380 4078
rect 64328 4014 64380 4020
rect 60004 3528 60056 3534
rect 60004 3470 60056 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 61200 3528 61252 3534
rect 61200 3470 61252 3476
rect 62028 3528 62080 3534
rect 62028 3470 62080 3476
rect 62396 3528 62448 3534
rect 62396 3470 62448 3476
rect 63040 3528 63092 3534
rect 63040 3470 63092 3476
rect 63592 3528 63644 3534
rect 63592 3470 63644 3476
rect 64236 3528 64288 3534
rect 64236 3470 64288 3476
rect 64616 3482 64644 11591
rect 64708 3874 64736 598946
rect 64800 9586 64828 607242
rect 66168 606552 66220 606558
rect 66168 606494 66220 606500
rect 66076 503736 66128 503742
rect 66076 503678 66128 503684
rect 65984 485852 66036 485858
rect 65984 485794 66036 485800
rect 65892 412684 65944 412690
rect 65892 412626 65944 412632
rect 65800 383716 65852 383722
rect 65800 383658 65852 383664
rect 65708 178084 65760 178090
rect 65708 178026 65760 178032
rect 65616 171148 65668 171154
rect 65616 171090 65668 171096
rect 64788 9580 64840 9586
rect 64788 9522 64840 9528
rect 65628 9246 65656 171090
rect 65720 12442 65748 178026
rect 65708 12436 65760 12442
rect 65708 12378 65760 12384
rect 65616 9240 65668 9246
rect 65616 9182 65668 9188
rect 64696 3868 64748 3874
rect 64696 3810 64748 3816
rect 58808 3460 58860 3466
rect 58808 3402 58860 3408
rect 59268 3460 59320 3466
rect 59268 3402 59320 3408
rect 56428 598 56548 626
rect 57624 598 57744 626
rect 56428 480 56456 598
rect 57624 480 57652 598
rect 58820 480 58848 3402
rect 60016 480 60044 3470
rect 61212 480 61240 3470
rect 62408 480 62436 3470
rect 63604 480 63632 3470
rect 64616 3454 64828 3482
rect 64800 480 64828 3454
rect 65812 3346 65840 383658
rect 65904 11762 65932 412626
rect 65892 11756 65944 11762
rect 65892 11698 65944 11704
rect 65996 6254 66024 485794
rect 66088 6322 66116 503678
rect 66180 99006 66208 606494
rect 67272 604988 67324 604994
rect 67272 604930 67324 604936
rect 67086 604072 67142 604081
rect 67086 604007 67142 604016
rect 66994 578232 67050 578241
rect 66994 578167 67050 578176
rect 67008 572665 67036 578167
rect 66994 572656 67050 572665
rect 66994 572591 67050 572600
rect 66994 534304 67050 534313
rect 66994 534239 67050 534248
rect 67008 531593 67036 534239
rect 66994 531584 67050 531593
rect 66994 531519 67050 531528
rect 66534 521656 66590 521665
rect 66534 521591 66590 521600
rect 66548 512281 66576 521591
rect 66534 512272 66590 512281
rect 66534 512207 66590 512216
rect 66626 510368 66682 510377
rect 66626 510303 66682 510312
rect 66640 500993 66668 510303
rect 66626 500984 66682 500993
rect 66626 500919 66682 500928
rect 66994 491192 67050 491201
rect 66994 491127 67050 491136
rect 67008 483721 67036 491127
rect 66994 483712 67050 483721
rect 66994 483647 67050 483656
rect 66994 478816 67050 478825
rect 66994 478751 67050 478760
rect 67008 469441 67036 478751
rect 66994 469432 67050 469441
rect 66994 469367 67050 469376
rect 66902 469160 66958 469169
rect 66902 469095 66958 469104
rect 66916 459785 66944 469095
rect 66902 459776 66958 459785
rect 66902 459711 66958 459720
rect 66718 446448 66774 446457
rect 66718 446383 66774 446392
rect 66732 434761 66760 446383
rect 66718 434752 66774 434761
rect 66718 434687 66774 434696
rect 66994 434616 67050 434625
rect 66994 434551 67050 434560
rect 67008 429865 67036 434551
rect 66994 429856 67050 429865
rect 66994 429791 67050 429800
rect 66902 398984 66958 398993
rect 66902 398919 66958 398928
rect 66916 396137 66944 398919
rect 66902 396128 66958 396137
rect 66902 396063 66958 396072
rect 66994 383480 67050 383489
rect 66994 383415 67050 383424
rect 67008 374105 67036 383415
rect 66994 374096 67050 374105
rect 66994 374031 67050 374040
rect 66718 336560 66774 336569
rect 66718 336495 66774 336504
rect 66732 327321 66760 336495
rect 66902 328400 66958 328409
rect 66902 328335 66958 328344
rect 66718 327312 66774 327321
rect 66718 327247 66774 327256
rect 66916 323649 66944 328335
rect 66902 323640 66958 323649
rect 66902 323575 66958 323584
rect 66994 299296 67050 299305
rect 66994 299231 67050 299240
rect 67008 290057 67036 299231
rect 66994 290048 67050 290057
rect 66994 289983 67050 289992
rect 66902 280120 66958 280129
rect 66902 280055 66958 280064
rect 66916 270745 66944 280055
rect 66996 277432 67048 277438
rect 66996 277374 67048 277380
rect 66902 270736 66958 270745
rect 66902 270671 66958 270680
rect 66904 251320 66956 251326
rect 66904 251262 66956 251268
rect 66718 201376 66774 201385
rect 66718 201311 66774 201320
rect 66732 195537 66760 201311
rect 66718 195528 66774 195537
rect 66718 195463 66774 195472
rect 66168 99000 66220 99006
rect 66168 98942 66220 98948
rect 66076 6316 66128 6322
rect 66076 6258 66128 6264
rect 65984 6248 66036 6254
rect 65984 6190 66036 6196
rect 66916 6186 66944 251262
rect 66904 6180 66956 6186
rect 66904 6122 66956 6128
rect 67008 3738 67036 277374
rect 67100 249762 67128 604007
rect 67180 603424 67232 603430
rect 67180 603366 67232 603372
rect 67088 249756 67140 249762
rect 67088 249698 67140 249704
rect 67086 240136 67142 240145
rect 67086 240071 67142 240080
rect 67100 222465 67128 240071
rect 67086 222456 67142 222465
rect 67086 222391 67142 222400
rect 67086 206000 67142 206009
rect 67086 205935 67142 205944
rect 67100 205465 67128 205935
rect 67086 205456 67142 205465
rect 67086 205391 67142 205400
rect 67086 191584 67142 191593
rect 67086 191519 67142 191528
rect 67100 174185 67128 191519
rect 67086 174176 67142 174185
rect 67086 174111 67142 174120
rect 67086 114472 67142 114481
rect 67086 114407 67142 114416
rect 67100 113393 67128 114407
rect 67086 113384 67142 113393
rect 67086 113319 67142 113328
rect 67086 103320 67142 103329
rect 67086 103255 67142 103264
rect 67100 89729 67128 103255
rect 67192 101794 67220 603366
rect 67180 101788 67232 101794
rect 67180 101730 67232 101736
rect 67284 98734 67312 604930
rect 67364 561740 67416 561746
rect 67364 561682 67416 561688
rect 67272 98728 67324 98734
rect 67272 98670 67324 98676
rect 67086 89720 67142 89729
rect 67086 89655 67142 89664
rect 67270 72448 67326 72457
rect 67270 72383 67326 72392
rect 67284 67697 67312 72383
rect 67270 67688 67326 67697
rect 67270 67623 67326 67632
rect 67086 57896 67142 57905
rect 67086 57831 67142 57840
rect 67100 50969 67128 57831
rect 67086 50960 67142 50969
rect 67086 50895 67142 50904
rect 67376 6526 67404 561682
rect 67468 100473 67496 700334
rect 68744 700324 68796 700330
rect 68744 700266 68796 700272
rect 67548 607368 67600 607374
rect 67548 607310 67600 607316
rect 67454 100464 67510 100473
rect 67454 100399 67510 100408
rect 67364 6520 67416 6526
rect 67364 6462 67416 6468
rect 67560 6458 67588 607310
rect 68284 604580 68336 604586
rect 68284 604522 68336 604528
rect 68296 151774 68324 604522
rect 68652 459604 68704 459610
rect 68652 459546 68704 459552
rect 68560 292596 68612 292602
rect 68560 292538 68612 292544
rect 68376 264988 68428 264994
rect 68376 264930 68428 264936
rect 68284 151768 68336 151774
rect 68284 151710 68336 151716
rect 68388 100638 68416 264930
rect 68468 251252 68520 251258
rect 68468 251194 68520 251200
rect 68480 165510 68508 251194
rect 68468 165504 68520 165510
rect 68468 165446 68520 165452
rect 68468 153264 68520 153270
rect 68468 153206 68520 153212
rect 68376 100632 68428 100638
rect 68376 100574 68428 100580
rect 68480 12170 68508 153206
rect 68468 12164 68520 12170
rect 68468 12106 68520 12112
rect 68572 9178 68600 292538
rect 68560 9172 68612 9178
rect 68560 9114 68612 9120
rect 67548 6452 67600 6458
rect 67548 6394 67600 6400
rect 68664 3942 68692 459546
rect 68756 223514 68784 700266
rect 69756 606620 69808 606626
rect 69756 606562 69808 606568
rect 68928 604716 68980 604722
rect 68928 604658 68980 604664
rect 68836 602472 68888 602478
rect 68836 602414 68888 602420
rect 68744 223508 68796 223514
rect 68744 223450 68796 223456
rect 68744 190528 68796 190534
rect 68744 190470 68796 190476
rect 68756 14482 68784 190470
rect 68848 100502 68876 602414
rect 68836 100496 68888 100502
rect 68836 100438 68888 100444
rect 68836 58744 68888 58750
rect 68836 58686 68888 58692
rect 68744 14476 68796 14482
rect 68744 14418 68796 14424
rect 68652 3936 68704 3942
rect 68652 3878 68704 3884
rect 66996 3732 67048 3738
rect 66996 3674 67048 3680
rect 68848 3534 68876 58686
rect 68940 6662 68968 604658
rect 69664 600636 69716 600642
rect 69664 600578 69716 600584
rect 69676 237386 69704 600578
rect 69768 425066 69796 606562
rect 70216 602608 70268 602614
rect 70216 602550 70268 602556
rect 69756 425060 69808 425066
rect 69756 425002 69808 425008
rect 69756 417444 69808 417450
rect 69756 417386 69808 417392
rect 69664 237380 69716 237386
rect 69664 237322 69716 237328
rect 69664 155236 69716 155242
rect 69664 155178 69716 155184
rect 68928 6656 68980 6662
rect 68928 6598 68980 6604
rect 69676 3913 69704 155178
rect 69768 100434 69796 417386
rect 69848 394732 69900 394738
rect 69848 394674 69900 394680
rect 69756 100428 69808 100434
rect 69756 100370 69808 100376
rect 69860 97850 69888 394674
rect 70124 295384 70176 295390
rect 70124 295326 70176 295332
rect 70032 273284 70084 273290
rect 70032 273226 70084 273232
rect 69940 237448 69992 237454
rect 69940 237390 69992 237396
rect 69848 97844 69900 97850
rect 69848 97786 69900 97792
rect 69952 4010 69980 237390
rect 70044 9042 70072 273226
rect 70032 9036 70084 9042
rect 70032 8978 70084 8984
rect 69940 4004 69992 4010
rect 69940 3946 69992 3952
rect 69662 3904 69718 3913
rect 69662 3839 69718 3848
rect 68284 3528 68336 3534
rect 67178 3496 67234 3505
rect 68284 3470 68336 3476
rect 68836 3528 68888 3534
rect 68836 3470 68888 3476
rect 67178 3431 67234 3440
rect 65812 3318 66024 3346
rect 65996 480 66024 3318
rect 67192 480 67220 3431
rect 68296 480 68324 3470
rect 70136 2922 70164 295326
rect 70228 99210 70256 602550
rect 70320 100298 70348 700606
rect 72804 698306 72832 703446
rect 81348 700596 81400 700602
rect 81348 700538 81400 700544
rect 75828 700528 75880 700534
rect 75828 700470 75880 700476
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659666 72924 659682
rect 72804 659660 72936 659666
rect 72804 659654 72884 659660
rect 72884 659602 72936 659608
rect 73068 659660 73120 659666
rect 73068 659602 73120 659608
rect 73080 656878 73108 659602
rect 73068 656872 73120 656878
rect 73068 656814 73120 656820
rect 72976 647284 73028 647290
rect 72976 647226 73028 647232
rect 72988 640422 73016 647226
rect 72976 640416 73028 640422
rect 72976 640358 73028 640364
rect 72792 640280 72844 640286
rect 72792 640222 72844 640228
rect 72804 637566 72832 640222
rect 72792 637560 72844 637566
rect 72792 637502 72844 637508
rect 73068 627972 73120 627978
rect 73068 627914 73120 627920
rect 73080 618322 73108 627914
rect 72976 618316 73028 618322
rect 72976 618258 73028 618264
rect 73068 618316 73120 618322
rect 73068 618258 73120 618264
rect 72988 618186 73016 618258
rect 72976 618180 73028 618186
rect 72976 618122 73028 618128
rect 73068 608728 73120 608734
rect 73068 608670 73120 608676
rect 71596 606212 71648 606218
rect 71596 606154 71648 606160
rect 71044 603764 71096 603770
rect 71044 603706 71096 603712
rect 70308 100292 70360 100298
rect 70308 100234 70360 100240
rect 70216 99204 70268 99210
rect 70216 99146 70268 99152
rect 71056 51066 71084 603706
rect 71504 602404 71556 602410
rect 71504 602346 71556 602352
rect 71136 600840 71188 600846
rect 71136 600782 71188 600788
rect 71148 194546 71176 600782
rect 71410 599992 71466 600001
rect 71410 599927 71466 599936
rect 71320 310548 71372 310554
rect 71320 310490 71372 310496
rect 71136 194540 71188 194546
rect 71136 194482 71188 194488
rect 71228 182232 71280 182238
rect 71228 182174 71280 182180
rect 71136 140072 71188 140078
rect 71136 140014 71188 140020
rect 71044 51060 71096 51066
rect 71044 51002 71096 51008
rect 71148 6866 71176 140014
rect 71240 8974 71268 182174
rect 71228 8968 71280 8974
rect 71228 8910 71280 8916
rect 71136 6860 71188 6866
rect 71136 6802 71188 6808
rect 70676 6588 70728 6594
rect 70676 6530 70728 6536
rect 69480 2916 69532 2922
rect 69480 2858 69532 2864
rect 70124 2916 70176 2922
rect 70124 2858 70176 2864
rect 69492 480 69520 2858
rect 70688 480 70716 6530
rect 71332 3369 71360 310490
rect 71424 99074 71452 599927
rect 71516 100366 71544 602346
rect 71608 101658 71636 606154
rect 72424 605328 72476 605334
rect 72424 605270 72476 605276
rect 71688 603628 71740 603634
rect 71688 603570 71740 603576
rect 71596 101652 71648 101658
rect 71596 101594 71648 101600
rect 71504 100360 71556 100366
rect 71504 100302 71556 100308
rect 71412 99068 71464 99074
rect 71412 99010 71464 99016
rect 71700 3641 71728 603570
rect 72332 200796 72384 200802
rect 72332 200738 72384 200744
rect 72344 190505 72372 200738
rect 72330 190496 72386 190505
rect 72330 190431 72386 190440
rect 72332 180804 72384 180810
rect 72332 180746 72384 180752
rect 72344 171222 72372 180746
rect 72332 171216 72384 171222
rect 72332 171158 72384 171164
rect 72436 165578 72464 605270
rect 72976 605260 73028 605266
rect 72976 605202 73028 605208
rect 72516 601792 72568 601798
rect 72516 601734 72568 601740
rect 72528 223582 72556 601734
rect 72884 600772 72936 600778
rect 72884 600714 72936 600720
rect 72792 586492 72844 586498
rect 72792 586434 72844 586440
rect 72804 576910 72832 586434
rect 72792 576904 72844 576910
rect 72792 576846 72844 576852
rect 72792 547868 72844 547874
rect 72792 547810 72844 547816
rect 72804 538286 72832 547810
rect 72792 538280 72844 538286
rect 72792 538222 72844 538228
rect 72792 489864 72844 489870
rect 72792 489806 72844 489812
rect 72804 480282 72832 489806
rect 72792 480276 72844 480282
rect 72792 480218 72844 480224
rect 72792 451240 72844 451246
rect 72792 451182 72844 451188
rect 72804 441726 72832 451182
rect 72792 441720 72844 441726
rect 72792 441662 72844 441668
rect 72792 431928 72844 431934
rect 72792 431870 72844 431876
rect 72804 422346 72832 431870
rect 72792 422340 72844 422346
rect 72792 422282 72844 422288
rect 72792 412616 72844 412622
rect 72792 412558 72844 412564
rect 72804 403034 72832 412558
rect 72792 403028 72844 403034
rect 72792 402970 72844 402976
rect 72792 393304 72844 393310
rect 72792 393246 72844 393252
rect 72804 383790 72832 393246
rect 72792 383784 72844 383790
rect 72792 383726 72844 383732
rect 72792 373992 72844 373998
rect 72792 373934 72844 373940
rect 72804 364410 72832 373934
rect 72792 364404 72844 364410
rect 72792 364346 72844 364352
rect 72608 336796 72660 336802
rect 72608 336738 72660 336744
rect 72516 223576 72568 223582
rect 72516 223518 72568 223524
rect 72516 211200 72568 211206
rect 72516 211142 72568 211148
rect 72424 165572 72476 165578
rect 72424 165514 72476 165520
rect 72424 161424 72476 161430
rect 72424 161366 72476 161372
rect 72436 151842 72464 161366
rect 72424 151836 72476 151842
rect 72424 151778 72476 151784
rect 72424 142112 72476 142118
rect 72424 142054 72476 142060
rect 72436 132530 72464 142054
rect 72424 132524 72476 132530
rect 72424 132466 72476 132472
rect 72424 127016 72476 127022
rect 72424 126958 72476 126964
rect 72332 122800 72384 122806
rect 72332 122742 72384 122748
rect 72344 113218 72372 122742
rect 72332 113212 72384 113218
rect 72332 113154 72384 113160
rect 72436 6730 72464 126958
rect 72528 77246 72556 211142
rect 72620 100774 72648 336738
rect 72792 315988 72844 315994
rect 72792 315930 72844 315936
rect 72804 306406 72832 315930
rect 72792 306400 72844 306406
rect 72792 306342 72844 306348
rect 72792 296676 72844 296682
rect 72792 296618 72844 296624
rect 72804 287094 72832 296618
rect 72792 287088 72844 287094
rect 72792 287030 72844 287036
rect 72792 281580 72844 281586
rect 72792 281522 72844 281528
rect 72700 277364 72752 277370
rect 72700 277306 72752 277312
rect 72712 267782 72740 277306
rect 72700 267776 72752 267782
rect 72700 267718 72752 267724
rect 72700 258800 72752 258806
rect 72700 258742 72752 258748
rect 72712 249150 72740 258742
rect 72700 249144 72752 249150
rect 72700 249086 72752 249092
rect 72700 239488 72752 239494
rect 72700 239430 72752 239436
rect 72712 229770 72740 239430
rect 72700 229764 72752 229770
rect 72700 229706 72752 229712
rect 72700 216980 72752 216986
rect 72700 216922 72752 216928
rect 72712 210458 72740 216922
rect 72700 210452 72752 210458
rect 72700 210394 72752 210400
rect 72700 193248 72752 193254
rect 72700 193190 72752 193196
rect 72608 100768 72660 100774
rect 72608 100710 72660 100716
rect 72516 77240 72568 77246
rect 72516 77182 72568 77188
rect 72712 14822 72740 193190
rect 72700 14816 72752 14822
rect 72700 14758 72752 14764
rect 72424 6724 72476 6730
rect 72424 6666 72476 6672
rect 71686 3632 71742 3641
rect 71686 3567 71742 3576
rect 71872 3528 71924 3534
rect 71872 3470 71924 3476
rect 71318 3360 71374 3369
rect 71318 3295 71374 3304
rect 71884 480 71912 3470
rect 72804 3466 72832 281522
rect 72896 101425 72924 600714
rect 72988 102678 73016 605202
rect 73080 586498 73108 608670
rect 74264 606280 74316 606286
rect 74264 606222 74316 606228
rect 74170 600808 74226 600817
rect 74170 600743 74226 600752
rect 73068 586492 73120 586498
rect 73068 586434 73120 586440
rect 73068 576904 73120 576910
rect 73068 576846 73120 576852
rect 73080 547874 73108 576846
rect 73068 547868 73120 547874
rect 73068 547810 73120 547816
rect 73068 538280 73120 538286
rect 73068 538222 73120 538228
rect 73080 489870 73108 538222
rect 73068 489864 73120 489870
rect 73068 489806 73120 489812
rect 73068 480276 73120 480282
rect 73068 480218 73120 480224
rect 73080 451246 73108 480218
rect 73068 451240 73120 451246
rect 73068 451182 73120 451188
rect 74080 448588 74132 448594
rect 74080 448530 74132 448536
rect 73068 441720 73120 441726
rect 73068 441662 73120 441668
rect 73080 431934 73108 441662
rect 73068 431928 73120 431934
rect 73068 431870 73120 431876
rect 73068 422340 73120 422346
rect 73068 422282 73120 422288
rect 73080 412622 73108 422282
rect 73068 412616 73120 412622
rect 73068 412558 73120 412564
rect 73068 403028 73120 403034
rect 73068 402970 73120 402976
rect 73080 393310 73108 402970
rect 73068 393304 73120 393310
rect 73068 393246 73120 393252
rect 73068 383784 73120 383790
rect 73068 383726 73120 383732
rect 73080 373998 73108 383726
rect 73068 373992 73120 373998
rect 73068 373934 73120 373940
rect 73068 364404 73120 364410
rect 73068 364346 73120 364352
rect 73080 315994 73108 364346
rect 73068 315988 73120 315994
rect 73068 315930 73120 315936
rect 73068 306400 73120 306406
rect 73068 306342 73120 306348
rect 73080 296682 73108 306342
rect 73068 296676 73120 296682
rect 73068 296618 73120 296624
rect 73068 287088 73120 287094
rect 73068 287030 73120 287036
rect 73080 277370 73108 287030
rect 73068 277364 73120 277370
rect 73068 277306 73120 277312
rect 73068 267776 73120 267782
rect 73068 267718 73120 267724
rect 73080 258806 73108 267718
rect 73068 258800 73120 258806
rect 73068 258742 73120 258748
rect 73068 249144 73120 249150
rect 73068 249086 73120 249092
rect 73080 239494 73108 249086
rect 73988 241528 74040 241534
rect 73988 241470 74040 241476
rect 73068 239488 73120 239494
rect 73068 239430 73120 239436
rect 73068 229764 73120 229770
rect 73068 229706 73120 229712
rect 73080 216986 73108 229706
rect 73068 216980 73120 216986
rect 73068 216922 73120 216928
rect 73068 210452 73120 210458
rect 73068 210394 73120 210400
rect 73080 200802 73108 210394
rect 73896 208412 73948 208418
rect 73896 208354 73948 208360
rect 73068 200796 73120 200802
rect 73068 200738 73120 200744
rect 73066 190496 73122 190505
rect 73066 190431 73122 190440
rect 73080 180810 73108 190431
rect 73068 180804 73120 180810
rect 73068 180746 73120 180752
rect 73068 171216 73120 171222
rect 73068 171158 73120 171164
rect 73080 161430 73108 171158
rect 73068 161424 73120 161430
rect 73068 161366 73120 161372
rect 73068 151836 73120 151842
rect 73068 151778 73120 151784
rect 73080 142118 73108 151778
rect 73068 142112 73120 142118
rect 73068 142054 73120 142060
rect 73068 132524 73120 132530
rect 73068 132466 73120 132472
rect 73080 122806 73108 132466
rect 73804 126268 73856 126274
rect 73804 126210 73856 126216
rect 73068 122800 73120 122806
rect 73068 122742 73120 122748
rect 73068 113212 73120 113218
rect 73068 113154 73120 113160
rect 73080 110430 73108 113154
rect 73068 110424 73120 110430
rect 73068 110366 73120 110372
rect 73816 109070 73844 126210
rect 73068 109064 73120 109070
rect 73068 109006 73120 109012
rect 73804 109064 73856 109070
rect 73804 109006 73856 109012
rect 72976 102672 73028 102678
rect 72976 102614 73028 102620
rect 72882 101416 72938 101425
rect 72882 101351 72938 101360
rect 72884 13116 72936 13122
rect 72884 13058 72936 13064
rect 72896 3534 72924 13058
rect 73080 9217 73108 109006
rect 73804 107908 73856 107914
rect 73804 107850 73856 107856
rect 73816 101561 73844 107850
rect 73802 101552 73858 101561
rect 73802 101487 73858 101496
rect 73908 14618 73936 208354
rect 73896 14612 73948 14618
rect 73896 14554 73948 14560
rect 73066 9208 73122 9217
rect 73066 9143 73122 9152
rect 74000 6390 74028 241470
rect 74092 69698 74120 448530
rect 74184 107914 74212 600743
rect 74172 107908 74224 107914
rect 74172 107850 74224 107856
rect 74276 107794 74304 606222
rect 74448 602200 74500 602206
rect 74448 602142 74500 602148
rect 74356 600908 74408 600914
rect 74356 600850 74408 600856
rect 74184 107766 74304 107794
rect 74184 102610 74212 107766
rect 74264 107704 74316 107710
rect 74264 107646 74316 107652
rect 74172 102604 74224 102610
rect 74172 102546 74224 102552
rect 74276 102134 74304 107646
rect 74264 102128 74316 102134
rect 74264 102070 74316 102076
rect 74080 69692 74132 69698
rect 74080 69634 74132 69640
rect 73988 6384 74040 6390
rect 73988 6326 74040 6332
rect 73250 3904 73306 3913
rect 73250 3839 73306 3848
rect 72884 3528 72936 3534
rect 73264 3505 73292 3839
rect 72884 3470 72936 3476
rect 73066 3496 73122 3505
rect 72792 3460 72844 3466
rect 73066 3431 73122 3440
rect 73250 3496 73306 3505
rect 73250 3431 73306 3440
rect 72792 3402 72844 3408
rect 73080 480 73108 3431
rect 74368 626 74396 600850
rect 74460 3738 74488 602142
rect 75552 601044 75604 601050
rect 75552 600986 75604 600992
rect 75460 518968 75512 518974
rect 75460 518910 75512 518916
rect 75368 456816 75420 456822
rect 75368 456758 75420 456764
rect 75276 357468 75328 357474
rect 75276 357410 75328 357416
rect 75184 178152 75236 178158
rect 75184 178094 75236 178100
rect 75196 102785 75224 178094
rect 75182 102776 75238 102785
rect 75182 102711 75238 102720
rect 75288 61606 75316 357410
rect 75380 78130 75408 456758
rect 75472 86290 75500 518910
rect 75564 101590 75592 600986
rect 75644 599820 75696 599826
rect 75644 599762 75696 599768
rect 75552 101584 75604 101590
rect 75552 101526 75604 101532
rect 75656 99142 75684 599762
rect 75736 577176 75788 577182
rect 75736 577118 75788 577124
rect 75644 99136 75696 99142
rect 75644 99078 75696 99084
rect 75460 86284 75512 86290
rect 75460 86226 75512 86232
rect 75368 78124 75420 78130
rect 75368 78066 75420 78072
rect 75276 61600 75328 61606
rect 75276 61542 75328 61548
rect 75748 24138 75776 577118
rect 75840 100230 75868 700470
rect 77208 700460 77260 700466
rect 77208 700402 77260 700408
rect 76564 600704 76616 600710
rect 76564 600646 76616 600652
rect 76576 324290 76604 600646
rect 76932 572756 76984 572762
rect 76932 572698 76984 572704
rect 76840 525836 76892 525842
rect 76840 525778 76892 525784
rect 76748 416832 76800 416838
rect 76748 416774 76800 416780
rect 76656 324352 76708 324358
rect 76656 324294 76708 324300
rect 76564 324284 76616 324290
rect 76564 324226 76616 324232
rect 76564 299532 76616 299538
rect 76564 299474 76616 299480
rect 76470 206000 76526 206009
rect 76470 205935 76526 205944
rect 76484 205465 76512 205935
rect 76470 205456 76526 205465
rect 76470 205391 76526 205400
rect 75828 100224 75880 100230
rect 75828 100166 75880 100172
rect 76576 73914 76604 299474
rect 76668 90370 76696 324294
rect 76656 90364 76708 90370
rect 76656 90306 76708 90312
rect 76564 73908 76616 73914
rect 76564 73850 76616 73856
rect 76760 40798 76788 416774
rect 76852 79354 76880 525778
rect 76944 101969 76972 572698
rect 77024 558952 77076 558958
rect 77024 558894 77076 558900
rect 76930 101960 76986 101969
rect 76930 101895 76986 101904
rect 77036 84930 77064 558894
rect 77116 500064 77168 500070
rect 77116 500006 77168 500012
rect 77024 84924 77076 84930
rect 77024 84866 77076 84872
rect 76840 79348 76892 79354
rect 76840 79290 76892 79296
rect 76748 40792 76800 40798
rect 76748 40734 76800 40740
rect 75736 24132 75788 24138
rect 75736 24074 75788 24080
rect 77128 10470 77156 500006
rect 77220 100609 77248 700402
rect 79876 617568 79928 617574
rect 79876 617510 79928 617516
rect 79324 605056 79376 605062
rect 79324 604998 79376 605004
rect 78678 599584 78734 599593
rect 78678 599519 78734 599528
rect 78692 599010 78720 599519
rect 78680 599004 78732 599010
rect 78680 598946 78732 598952
rect 78678 595776 78734 595785
rect 78678 595711 78734 595720
rect 78692 594114 78720 595711
rect 78680 594108 78732 594114
rect 78680 594050 78732 594056
rect 78678 592240 78734 592249
rect 78678 592175 78734 592184
rect 78692 592074 78720 592175
rect 78680 592068 78732 592074
rect 78680 592010 78732 592016
rect 78954 577552 79010 577561
rect 78954 577487 79010 577496
rect 78968 577182 78996 577487
rect 78956 577176 79008 577182
rect 78956 577118 79008 577124
rect 78770 574016 78826 574025
rect 78770 573951 78826 573960
rect 78784 572762 78812 573951
rect 78772 572756 78824 572762
rect 78772 572698 78824 572704
rect 78678 570208 78734 570217
rect 78678 570143 78734 570152
rect 78692 569974 78720 570143
rect 78680 569968 78732 569974
rect 78680 569910 78732 569916
rect 78678 566672 78734 566681
rect 78678 566607 78734 566616
rect 78692 565894 78720 566607
rect 78680 565888 78732 565894
rect 78680 565830 78732 565836
rect 78678 562864 78734 562873
rect 78678 562799 78734 562808
rect 78692 561746 78720 562799
rect 78680 561740 78732 561746
rect 78680 561682 78732 561688
rect 78678 555792 78734 555801
rect 78678 555727 78734 555736
rect 78692 554810 78720 555727
rect 78680 554804 78732 554810
rect 78680 554746 78732 554752
rect 78678 526416 78734 526425
rect 78678 526351 78734 526360
rect 78692 525842 78720 526351
rect 78680 525836 78732 525842
rect 78680 525778 78732 525784
rect 78862 519072 78918 519081
rect 78862 519007 78918 519016
rect 78876 518974 78904 519007
rect 78864 518968 78916 518974
rect 78864 518910 78916 518916
rect 78678 511728 78734 511737
rect 78678 511663 78734 511672
rect 78692 510678 78720 511663
rect 78680 510672 78732 510678
rect 78680 510614 78732 510620
rect 78678 508192 78734 508201
rect 78678 508127 78734 508136
rect 78692 507890 78720 508127
rect 78680 507884 78732 507890
rect 78680 507826 78732 507832
rect 78678 504656 78734 504665
rect 78678 504591 78734 504600
rect 78692 503742 78720 504591
rect 78680 503736 78732 503742
rect 78680 503678 78732 503684
rect 79046 500848 79102 500857
rect 79046 500783 79102 500792
rect 79060 500070 79088 500783
rect 79048 500064 79100 500070
rect 79048 500006 79100 500012
rect 78678 497312 78734 497321
rect 78678 497247 78734 497256
rect 78692 496874 78720 497247
rect 78680 496868 78732 496874
rect 78680 496810 78732 496816
rect 78678 486160 78734 486169
rect 78678 486095 78734 486104
rect 78692 485858 78720 486095
rect 78680 485852 78732 485858
rect 78680 485794 78732 485800
rect 78678 479088 78734 479097
rect 78678 479023 78734 479032
rect 78692 478922 78720 479023
rect 78680 478916 78732 478922
rect 78680 478858 78732 478864
rect 78680 471980 78732 471986
rect 78680 471922 78732 471928
rect 78692 471753 78720 471922
rect 78678 471744 78734 471753
rect 78678 471679 78734 471688
rect 78678 460592 78734 460601
rect 78678 460527 78734 460536
rect 78692 459610 78720 460527
rect 78680 459604 78732 459610
rect 78680 459546 78732 459552
rect 78678 457056 78734 457065
rect 78678 456991 78734 457000
rect 78692 456822 78720 456991
rect 78680 456816 78732 456822
rect 78680 456758 78732 456764
rect 78678 449712 78734 449721
rect 78678 449647 78734 449656
rect 78692 448594 78720 449647
rect 78680 448588 78732 448594
rect 78680 448530 78732 448536
rect 78678 446176 78734 446185
rect 78678 446111 78734 446120
rect 78692 445806 78720 446111
rect 78680 445800 78732 445806
rect 78680 445742 78732 445748
rect 78678 442368 78734 442377
rect 78678 442303 78734 442312
rect 78692 441658 78720 442303
rect 78680 441652 78732 441658
rect 78680 441594 78732 441600
rect 78494 438832 78550 438841
rect 78494 438767 78550 438776
rect 78402 395040 78458 395049
rect 78402 394975 78458 394984
rect 78218 307184 78274 307193
rect 78218 307119 78274 307128
rect 78126 303648 78182 303657
rect 78126 303583 78182 303592
rect 77942 197840 77998 197849
rect 77942 197775 77998 197784
rect 77206 100600 77262 100609
rect 77206 100535 77262 100544
rect 77956 98802 77984 197775
rect 78034 161120 78090 161129
rect 78034 161055 78090 161064
rect 77944 98796 77996 98802
rect 77944 98738 77996 98744
rect 77206 90400 77262 90409
rect 77206 90335 77262 90344
rect 77116 10464 77168 10470
rect 77116 10406 77168 10412
rect 75458 3768 75514 3777
rect 74448 3732 74500 3738
rect 75458 3703 75514 3712
rect 74448 3674 74500 3680
rect 74276 598 74396 626
rect 74276 480 74304 598
rect 75472 480 75500 3703
rect 77220 3398 77248 90335
rect 78048 43450 78076 161055
rect 78140 89078 78168 303583
rect 78128 89072 78180 89078
rect 78128 89014 78180 89020
rect 78232 83638 78260 307119
rect 78312 245608 78364 245614
rect 78312 245550 78364 245556
rect 78220 83632 78272 83638
rect 78220 83574 78272 83580
rect 78036 43444 78088 43450
rect 78036 43386 78088 43392
rect 78324 3398 78352 245550
rect 78416 99278 78444 394975
rect 78404 99272 78456 99278
rect 78404 99214 78456 99220
rect 78508 50386 78536 438767
rect 78586 435024 78642 435033
rect 78586 434959 78642 434968
rect 78496 50380 78548 50386
rect 78496 50322 78548 50328
rect 78600 32434 78628 434959
rect 78678 431488 78734 431497
rect 78678 431423 78734 431432
rect 78692 430642 78720 431423
rect 78680 430636 78732 430642
rect 78680 430578 78732 430584
rect 78678 427952 78734 427961
rect 78678 427887 78734 427896
rect 78692 427854 78720 427887
rect 78680 427848 78732 427854
rect 78680 427790 78732 427796
rect 78678 420608 78734 420617
rect 78678 420543 78734 420552
rect 78692 419558 78720 420543
rect 78680 419552 78732 419558
rect 78680 419494 78732 419500
rect 78680 416832 78732 416838
rect 78678 416800 78680 416809
rect 78732 416800 78734 416809
rect 78678 416735 78734 416744
rect 78678 413264 78734 413273
rect 78678 413199 78734 413208
rect 78692 412690 78720 413199
rect 78680 412684 78732 412690
rect 78680 412626 78732 412632
rect 78678 405920 78734 405929
rect 78678 405855 78734 405864
rect 78692 405754 78720 405855
rect 78680 405748 78732 405754
rect 78680 405690 78732 405696
rect 78678 402384 78734 402393
rect 78678 402319 78734 402328
rect 78692 401674 78720 402319
rect 78680 401668 78732 401674
rect 78680 401610 78732 401616
rect 78678 398576 78734 398585
rect 78678 398511 78734 398520
rect 78692 397526 78720 398511
rect 78680 397520 78732 397526
rect 78680 397462 78732 397468
rect 78678 387696 78734 387705
rect 78678 387631 78734 387640
rect 78692 386442 78720 387631
rect 78680 386436 78732 386442
rect 78680 386378 78732 386384
rect 78678 383888 78734 383897
rect 78678 383823 78734 383832
rect 78692 383722 78720 383823
rect 78680 383716 78732 383722
rect 78680 383658 78732 383664
rect 78678 369472 78734 369481
rect 78678 369407 78734 369416
rect 78692 368558 78720 369407
rect 78680 368552 78732 368558
rect 78680 368494 78732 368500
rect 78678 362128 78734 362137
rect 78678 362063 78734 362072
rect 78692 361622 78720 362063
rect 78680 361616 78732 361622
rect 78680 361558 78732 361564
rect 78678 358320 78734 358329
rect 78678 358255 78734 358264
rect 78692 357474 78720 358255
rect 78680 357468 78732 357474
rect 78680 357410 78732 357416
rect 78680 351892 78732 351898
rect 78680 351834 78732 351840
rect 78692 351257 78720 351834
rect 78678 351248 78734 351257
rect 78678 351183 78734 351192
rect 78678 347440 78734 347449
rect 78678 347375 78734 347384
rect 78692 346458 78720 347375
rect 78680 346452 78732 346458
rect 78680 346394 78732 346400
rect 78678 336560 78734 336569
rect 78678 336495 78734 336504
rect 78692 335374 78720 336495
rect 78680 335368 78732 335374
rect 78680 335310 78732 335316
rect 78678 332752 78734 332761
rect 78678 332687 78734 332696
rect 78692 332654 78720 332687
rect 78680 332648 78732 332654
rect 78680 332590 78732 332596
rect 78680 329792 78732 329798
rect 78680 329734 78732 329740
rect 78692 329225 78720 329734
rect 78678 329216 78734 329225
rect 78678 329151 78734 329160
rect 78678 325680 78734 325689
rect 78678 325615 78734 325624
rect 78692 324358 78720 325615
rect 78680 324352 78732 324358
rect 78680 324294 78732 324300
rect 78680 322924 78732 322930
rect 78680 322866 78732 322872
rect 78692 321881 78720 322866
rect 78678 321872 78734 321881
rect 78678 321807 78734 321816
rect 78678 318336 78734 318345
rect 78678 318271 78734 318280
rect 78692 317490 78720 318271
rect 78680 317484 78732 317490
rect 78680 317426 78732 317432
rect 78678 310992 78734 311001
rect 78678 310927 78734 310936
rect 78692 310554 78720 310927
rect 78680 310548 78732 310554
rect 78680 310490 78732 310496
rect 79230 300112 79286 300121
rect 79230 300047 79286 300056
rect 79244 299538 79272 300047
rect 79232 299532 79284 299538
rect 79232 299474 79284 299480
rect 78678 296304 78734 296313
rect 78678 296239 78734 296248
rect 78692 295390 78720 296239
rect 78680 295384 78732 295390
rect 78680 295326 78732 295332
rect 78678 292768 78734 292777
rect 78678 292703 78734 292712
rect 78692 292602 78720 292703
rect 78680 292596 78732 292602
rect 78680 292538 78732 292544
rect 78678 281616 78734 281625
rect 78678 281551 78680 281560
rect 78732 281551 78734 281560
rect 78680 281522 78732 281528
rect 78678 278080 78734 278089
rect 78678 278015 78734 278024
rect 78692 277438 78720 278015
rect 78680 277432 78732 277438
rect 78680 277374 78732 277380
rect 78678 274544 78734 274553
rect 78678 274479 78734 274488
rect 78692 273290 78720 274479
rect 78680 273284 78732 273290
rect 78680 273226 78732 273232
rect 78678 267200 78734 267209
rect 78678 267135 78734 267144
rect 78692 266422 78720 267135
rect 78680 266416 78732 266422
rect 78680 266358 78732 266364
rect 78680 263560 78732 263566
rect 78680 263502 78732 263508
rect 78692 263401 78720 263502
rect 78678 263392 78734 263401
rect 78678 263327 78734 263336
rect 78678 252512 78734 252521
rect 78678 252447 78734 252456
rect 78692 251326 78720 252447
rect 78680 251320 78732 251326
rect 78680 251262 78732 251268
rect 78680 249756 78732 249762
rect 78680 249698 78732 249704
rect 78692 248985 78720 249698
rect 78678 248976 78734 248985
rect 78678 248911 78734 248920
rect 78678 241632 78734 241641
rect 78678 241567 78734 241576
rect 78692 241534 78720 241567
rect 78680 241528 78732 241534
rect 78680 241470 78732 241476
rect 78678 237824 78734 237833
rect 78678 237759 78734 237768
rect 78692 237454 78720 237759
rect 78680 237448 78732 237454
rect 78680 237390 78732 237396
rect 78678 234288 78734 234297
rect 78678 234223 78734 234232
rect 78692 233306 78720 234223
rect 78680 233300 78732 233306
rect 78680 233242 78732 233248
rect 78678 230480 78734 230489
rect 78678 230415 78734 230424
rect 78692 229158 78720 230415
rect 78680 229152 78732 229158
rect 78680 229094 78732 229100
rect 78680 223508 78732 223514
rect 78680 223450 78732 223456
rect 78692 223417 78720 223450
rect 78678 223408 78734 223417
rect 78678 223343 78734 223352
rect 78678 212256 78734 212265
rect 78678 212191 78734 212200
rect 78692 211206 78720 212191
rect 78680 211200 78732 211206
rect 78680 211142 78732 211148
rect 78678 208720 78734 208729
rect 78678 208655 78734 208664
rect 78692 208418 78720 208655
rect 78680 208412 78732 208418
rect 78680 208354 78732 208360
rect 78678 194032 78734 194041
rect 78678 193967 78734 193976
rect 78692 193254 78720 193967
rect 78680 193248 78732 193254
rect 78680 193190 78732 193196
rect 78680 190528 78732 190534
rect 78678 190496 78680 190505
rect 78732 190496 78734 190505
rect 78678 190431 78734 190440
rect 79230 186688 79286 186697
rect 79230 186623 79286 186632
rect 78678 183152 78734 183161
rect 78678 183087 78734 183096
rect 78692 182238 78720 183087
rect 78680 182232 78732 182238
rect 78680 182174 78732 182180
rect 78678 179344 78734 179353
rect 78678 179279 78734 179288
rect 78692 178090 78720 179279
rect 78680 178084 78732 178090
rect 78680 178026 78732 178032
rect 78678 172272 78734 172281
rect 78678 172207 78734 172216
rect 78692 171154 78720 172207
rect 78680 171148 78732 171154
rect 78680 171090 78732 171096
rect 78680 165504 78732 165510
rect 78680 165446 78732 165452
rect 78692 164937 78720 165446
rect 78678 164928 78734 164937
rect 78678 164863 78734 164872
rect 78680 158704 78732 158710
rect 78680 158646 78732 158652
rect 78692 157593 78720 158646
rect 78678 157584 78734 157593
rect 78678 157519 78734 157528
rect 78678 153776 78734 153785
rect 78678 153711 78734 153720
rect 78692 153270 78720 153711
rect 78680 153264 78732 153270
rect 78680 153206 78732 153212
rect 78678 150240 78734 150249
rect 78678 150175 78734 150184
rect 78692 149122 78720 150175
rect 78680 149116 78732 149122
rect 78680 149058 78732 149064
rect 78678 146704 78734 146713
rect 78678 146639 78734 146648
rect 78692 146334 78720 146639
rect 78680 146328 78732 146334
rect 78680 146270 78732 146276
rect 78678 132016 78734 132025
rect 78678 131951 78734 131960
rect 78692 131170 78720 131951
rect 78680 131164 78732 131170
rect 78680 131106 78732 131112
rect 78678 128208 78734 128217
rect 78678 128143 78734 128152
rect 78692 127022 78720 128143
rect 78680 127016 78732 127022
rect 78680 126958 78732 126964
rect 79138 113792 79194 113801
rect 79138 113727 79194 113736
rect 78680 110424 78732 110430
rect 78680 110366 78732 110372
rect 78692 109993 78720 110366
rect 78678 109984 78734 109993
rect 78678 109919 78734 109928
rect 79152 94518 79180 113727
rect 79140 94512 79192 94518
rect 79140 94454 79192 94460
rect 78680 93152 78732 93158
rect 78680 93094 78732 93100
rect 78588 32428 78640 32434
rect 78588 32370 78640 32376
rect 78692 3482 78720 93094
rect 79244 83502 79272 186623
rect 79336 126274 79364 604998
rect 79416 603696 79468 603702
rect 79416 603638 79468 603644
rect 79428 187785 79456 603638
rect 79598 559328 79654 559337
rect 79598 559263 79654 559272
rect 79612 558958 79640 559263
rect 79600 558952 79652 558958
rect 79600 558894 79652 558900
rect 79888 530233 79916 617510
rect 81256 607232 81308 607238
rect 81256 607174 81308 607180
rect 81164 606348 81216 606354
rect 81164 606290 81216 606296
rect 79968 604784 80020 604790
rect 79968 604726 80020 604732
rect 79874 530224 79930 530233
rect 79874 530159 79930 530168
rect 79506 493504 79562 493513
rect 79506 493439 79562 493448
rect 79520 245614 79548 493439
rect 79874 391232 79930 391241
rect 79874 391167 79930 391176
rect 79782 343904 79838 343913
rect 79782 343839 79838 343848
rect 79690 259856 79746 259865
rect 79690 259791 79746 259800
rect 79508 245608 79560 245614
rect 79508 245550 79560 245556
rect 79704 244202 79732 259791
rect 79612 244174 79732 244202
rect 79612 225026 79640 244174
rect 79520 224998 79640 225026
rect 79520 210458 79548 224998
rect 79598 219600 79654 219609
rect 79598 219535 79654 219544
rect 79508 210452 79560 210458
rect 79508 210394 79560 210400
rect 79508 199572 79560 199578
rect 79508 199514 79560 199520
rect 79520 190534 79548 199514
rect 79508 190528 79560 190534
rect 79508 190470 79560 190476
rect 79414 187776 79470 187785
rect 79414 187711 79470 187720
rect 79508 180804 79560 180810
rect 79508 180746 79560 180752
rect 79520 171154 79548 180746
rect 79508 171148 79560 171154
rect 79508 171090 79560 171096
rect 79508 166320 79560 166326
rect 79508 166262 79560 166268
rect 79520 151842 79548 166262
rect 79508 151836 79560 151842
rect 79508 151778 79560 151784
rect 79506 142896 79562 142905
rect 79506 142831 79562 142840
rect 79324 126268 79376 126274
rect 79324 126210 79376 126216
rect 79414 124672 79470 124681
rect 79414 124607 79470 124616
rect 79428 91798 79456 124607
rect 79416 91792 79468 91798
rect 79416 91734 79468 91740
rect 79232 83496 79284 83502
rect 79232 83438 79284 83444
rect 79520 42090 79548 142831
rect 79508 42084 79560 42090
rect 79508 42026 79560 42032
rect 79612 20058 79640 219535
rect 79692 210452 79744 210458
rect 79692 210394 79744 210400
rect 79704 199578 79732 210394
rect 79692 199572 79744 199578
rect 79692 199514 79744 199520
rect 79692 190528 79744 190534
rect 79692 190470 79744 190476
rect 79704 180810 79732 190470
rect 79692 180804 79744 180810
rect 79692 180746 79744 180752
rect 79692 171148 79744 171154
rect 79692 171090 79744 171096
rect 79704 166326 79732 171090
rect 79692 166320 79744 166326
rect 79692 166262 79744 166268
rect 79692 151836 79744 151842
rect 79692 151778 79744 151784
rect 79704 142118 79732 151778
rect 79692 142112 79744 142118
rect 79692 142054 79744 142060
rect 79692 132524 79744 132530
rect 79692 132466 79744 132472
rect 79704 122806 79732 132466
rect 79692 122800 79744 122806
rect 79692 122742 79744 122748
rect 79692 113212 79744 113218
rect 79692 113154 79744 113160
rect 79704 102270 79732 113154
rect 79692 102264 79744 102270
rect 79692 102206 79744 102212
rect 79796 97306 79824 343839
rect 79888 102406 79916 391167
rect 79980 176730 80008 604726
rect 80702 601352 80758 601361
rect 80702 601287 80758 601296
rect 80716 600953 80744 601287
rect 81072 600976 81124 600982
rect 80702 600944 80758 600953
rect 81072 600918 81124 600924
rect 80702 600879 80758 600888
rect 80978 482624 81034 482633
rect 80978 482559 81034 482568
rect 80886 340096 80942 340105
rect 80886 340031 80942 340040
rect 80794 201376 80850 201385
rect 80794 201311 80850 201320
rect 79968 176724 80020 176730
rect 79968 176666 80020 176672
rect 80704 176724 80756 176730
rect 80704 176666 80756 176672
rect 79968 142112 80020 142118
rect 79968 142054 80020 142060
rect 79980 132530 80008 142054
rect 79968 132524 80020 132530
rect 79968 132466 80020 132472
rect 79968 122800 80020 122806
rect 79968 122742 80020 122748
rect 79980 113218 80008 122742
rect 79968 113212 80020 113218
rect 79968 113154 80020 113160
rect 79876 102400 79928 102406
rect 79876 102342 79928 102348
rect 79876 102264 79928 102270
rect 79876 102206 79928 102212
rect 79784 97300 79836 97306
rect 79784 97242 79836 97248
rect 79888 86986 79916 102206
rect 80716 98938 80744 176666
rect 80704 98932 80756 98938
rect 80704 98874 80756 98880
rect 79796 86958 79916 86986
rect 79796 85542 79824 86958
rect 79784 85536 79836 85542
rect 79784 85478 79836 85484
rect 79968 75948 80020 75954
rect 79968 75890 80020 75896
rect 79980 67658 80008 75890
rect 79784 67652 79836 67658
rect 79784 67594 79836 67600
rect 79968 67652 80020 67658
rect 79968 67594 80020 67600
rect 79796 60738 79824 67594
rect 79704 60722 79824 60738
rect 79692 60716 79824 60722
rect 79744 60710 79824 60716
rect 79876 60716 79928 60722
rect 79692 60658 79744 60664
rect 79876 60658 79928 60664
rect 79888 57934 79916 60658
rect 79876 57928 79928 57934
rect 79876 57870 79928 57876
rect 79876 50924 79928 50930
rect 79876 50866 79928 50872
rect 79888 37942 79916 50866
rect 79876 37936 79928 37942
rect 79876 37878 79928 37884
rect 79600 20052 79652 20058
rect 79600 19994 79652 20000
rect 80808 18698 80836 201311
rect 80900 51746 80928 340031
rect 80992 101522 81020 482559
rect 81084 179382 81112 600918
rect 81072 179376 81124 179382
rect 81072 179318 81124 179324
rect 81072 120080 81124 120086
rect 81072 120022 81124 120028
rect 81084 102746 81112 120022
rect 81072 102740 81124 102746
rect 81072 102682 81124 102688
rect 80980 101516 81032 101522
rect 80980 101458 81032 101464
rect 81176 98666 81204 606290
rect 81164 98660 81216 98666
rect 81164 98602 81216 98608
rect 80888 51740 80940 51746
rect 80888 51682 80940 51688
rect 80796 18692 80848 18698
rect 80796 18634 80848 18640
rect 81268 12374 81296 607174
rect 81360 100162 81388 700538
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 700738 137876 703520
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 138664 700732 138716 700738
rect 138664 700674 138716 700680
rect 88340 699712 88392 699718
rect 88340 699654 88392 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 104900 699712 104952 699718
rect 104900 699654 104952 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 81716 626612 81768 626618
rect 81716 626554 81768 626560
rect 81624 607912 81676 607918
rect 81624 607854 81676 607860
rect 81440 603832 81492 603838
rect 81440 603774 81492 603780
rect 81452 596834 81480 603774
rect 81440 596828 81492 596834
rect 81440 596770 81492 596776
rect 81438 464400 81494 464409
rect 81438 464335 81494 464344
rect 81348 100156 81400 100162
rect 81348 100098 81400 100104
rect 81452 100026 81480 464335
rect 81530 409456 81586 409465
rect 81530 409391 81586 409400
rect 81440 100020 81492 100026
rect 81440 99962 81492 99968
rect 81440 97368 81492 97374
rect 81440 97310 81492 97316
rect 81256 12368 81308 12374
rect 81256 12310 81308 12316
rect 80244 4072 80296 4078
rect 80244 4014 80296 4020
rect 78692 3454 79088 3482
rect 76656 3392 76708 3398
rect 76656 3334 76708 3340
rect 77208 3392 77260 3398
rect 77208 3334 77260 3340
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 78312 3392 78364 3398
rect 78312 3334 78364 3340
rect 76668 480 76696 3334
rect 77864 480 77892 3334
rect 79060 480 79088 3454
rect 80256 480 80284 4014
rect 81452 480 81480 97310
rect 81544 56030 81572 409391
rect 81636 314537 81664 607854
rect 81728 380361 81756 626554
rect 82084 606144 82136 606150
rect 82084 606086 82136 606092
rect 81714 380352 81770 380361
rect 81714 380287 81770 380296
rect 81622 314528 81678 314537
rect 81622 314463 81678 314472
rect 81622 270736 81678 270745
rect 81622 270671 81678 270680
rect 81532 56024 81584 56030
rect 81532 55966 81584 55972
rect 81636 49094 81664 270671
rect 81714 216064 81770 216073
rect 81714 215999 81770 216008
rect 81728 68406 81756 215999
rect 81900 179376 81952 179382
rect 81900 179318 81952 179324
rect 81806 168464 81862 168473
rect 81806 168399 81862 168408
rect 81716 68400 81768 68406
rect 81716 68342 81768 68348
rect 81624 49088 81676 49094
rect 81624 49030 81676 49036
rect 81820 22778 81848 168399
rect 81912 120086 81940 179318
rect 82096 155281 82124 606086
rect 86408 605940 86460 605946
rect 86408 605882 86460 605888
rect 82268 605192 82320 605198
rect 82268 605134 82320 605140
rect 82176 602268 82228 602274
rect 82176 602210 82228 602216
rect 82082 155272 82138 155281
rect 82188 155242 82216 602210
rect 82280 178158 82308 605134
rect 83280 605124 83332 605130
rect 83280 605066 83332 605072
rect 83188 603288 83240 603294
rect 83188 603230 83240 603236
rect 83200 592770 83228 603230
rect 83292 596850 83320 605066
rect 83464 602064 83516 602070
rect 83464 602006 83516 602012
rect 83370 601352 83426 601361
rect 83370 601287 83426 601296
rect 83384 600409 83412 601287
rect 83476 601202 83504 602006
rect 86420 601868 86448 605882
rect 88352 603242 88380 699654
rect 93766 605976 93822 605985
rect 93766 605911 93822 605920
rect 88260 603214 88380 603242
rect 88260 602478 88288 603214
rect 88800 603152 88852 603158
rect 88800 603094 88852 603100
rect 88340 603084 88392 603090
rect 88340 603026 88392 603032
rect 88248 602472 88300 602478
rect 88248 602414 88300 602420
rect 88352 602313 88380 603026
rect 88338 602304 88394 602313
rect 88338 602239 88394 602248
rect 88812 601868 88840 603094
rect 93780 601868 93808 605911
rect 101128 604716 101180 604722
rect 101128 604658 101180 604664
rect 98736 603900 98788 603906
rect 98736 603842 98788 603848
rect 96160 603764 96212 603770
rect 96160 603706 96212 603712
rect 96172 601868 96200 603706
rect 97908 603492 97960 603498
rect 97908 603434 97960 603440
rect 92388 601656 92440 601662
rect 92388 601598 92440 601604
rect 92400 601361 92428 601598
rect 92386 601352 92442 601361
rect 83660 601310 83858 601338
rect 91112 601322 91218 601338
rect 91100 601316 91218 601322
rect 83476 601174 83596 601202
rect 83464 601112 83516 601118
rect 83464 601054 83516 601060
rect 83370 600400 83426 600409
rect 83370 600335 83426 600344
rect 83476 600030 83504 601054
rect 83464 600024 83516 600030
rect 83464 599966 83516 599972
rect 83292 596822 83504 596850
rect 82924 592742 83228 592770
rect 82924 592686 82952 592742
rect 82912 592680 82964 592686
rect 82912 592622 82964 592628
rect 83476 591954 83504 596822
rect 83384 591926 83504 591954
rect 83384 584474 83412 591926
rect 83292 584446 83412 584474
rect 83292 579578 83320 584446
rect 83108 579550 83320 579578
rect 83108 569956 83136 579550
rect 83108 569928 83412 569956
rect 83384 563122 83412 569928
rect 83292 563094 83412 563122
rect 83292 553466 83320 563094
rect 83292 553438 83412 553466
rect 83384 543810 83412 553438
rect 83292 543782 83412 543810
rect 83292 534154 83320 543782
rect 83292 534126 83412 534154
rect 83384 524498 83412 534126
rect 83292 524470 83412 524498
rect 83292 514842 83320 524470
rect 83292 514814 83412 514842
rect 82912 507884 82964 507890
rect 83384 507872 83412 514814
rect 82964 507844 83412 507872
rect 82912 507826 82964 507832
rect 83568 506274 83596 601174
rect 83660 601118 83688 601310
rect 91152 601310 91218 601316
rect 97920 601322 97948 603434
rect 98748 601868 98776 603842
rect 101140 601868 101168 604658
rect 103702 604480 103758 604489
rect 103702 604415 103758 604424
rect 103716 601868 103744 604415
rect 104912 602426 104940 699654
rect 138676 614786 138704 700674
rect 154132 700670 154160 703520
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 170324 695502 170352 703520
rect 202800 697610 202828 703520
rect 218992 700602 219020 703520
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 235184 700534 235212 703520
rect 235172 700528 235224 700534
rect 235172 700470 235224 700476
rect 267660 700369 267688 703520
rect 283852 700534 283880 703520
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 298744 700528 298796 700534
rect 298744 700470 298796 700476
rect 267646 700360 267702 700369
rect 267646 700295 267702 700304
rect 259368 698964 259420 698970
rect 259368 698906 259420 698912
rect 202788 697604 202840 697610
rect 202788 697546 202840 697552
rect 169944 695496 169996 695502
rect 169944 695438 169996 695444
rect 170312 695496 170364 695502
rect 170312 695438 170364 695444
rect 169956 687954 169984 695438
rect 169944 687948 169996 687954
rect 169944 687890 169996 687896
rect 170128 687948 170180 687954
rect 170128 687890 170180 687896
rect 170140 683233 170168 687890
rect 169758 683224 169814 683233
rect 169758 683159 169814 683168
rect 170126 683224 170182 683233
rect 170126 683159 170182 683168
rect 169772 683126 169800 683159
rect 169760 683120 169812 683126
rect 169760 683062 169812 683068
rect 188342 674112 188398 674121
rect 188342 674047 188398 674056
rect 173900 674008 173952 674014
rect 173898 673976 173900 673985
rect 178316 674008 178368 674014
rect 173952 673976 173954 673985
rect 178316 673950 178368 673956
rect 173898 673911 173954 673920
rect 178328 673849 178356 673950
rect 188356 673849 188384 674047
rect 154578 673840 154634 673849
rect 166906 673840 166962 673849
rect 154578 673775 154580 673784
rect 154632 673775 154634 673784
rect 162216 673804 162268 673810
rect 154580 673746 154632 673752
rect 166906 673775 166962 673784
rect 178314 673840 178370 673849
rect 178314 673775 178370 673784
rect 188342 673840 188398 673849
rect 188342 673775 188398 673784
rect 162216 673746 162268 673752
rect 162228 673577 162256 673746
rect 166920 673577 166948 673775
rect 162214 673568 162270 673577
rect 162214 673503 162270 673512
rect 166906 673568 166962 673577
rect 166906 673503 166962 673512
rect 170220 666596 170272 666602
rect 170220 666538 170272 666544
rect 170232 659682 170260 666538
rect 170048 659654 170260 659682
rect 170048 647290 170076 659654
rect 177948 650072 178000 650078
rect 177948 650014 178000 650020
rect 169944 647284 169996 647290
rect 169944 647226 169996 647232
rect 170036 647284 170088 647290
rect 170036 647226 170088 647232
rect 169956 640422 169984 647226
rect 169944 640416 169996 640422
rect 169944 640358 169996 640364
rect 170036 640416 170088 640422
rect 170036 640358 170088 640364
rect 170048 630698 170076 640358
rect 169852 630692 169904 630698
rect 169852 630634 169904 630640
rect 170036 630692 170088 630698
rect 170036 630634 170088 630640
rect 169864 630578 169892 630634
rect 169864 630550 169984 630578
rect 169956 621058 169984 630550
rect 169956 621030 170076 621058
rect 138664 614780 138716 614786
rect 138664 614722 138716 614728
rect 170048 611386 170076 621030
rect 169760 611380 169812 611386
rect 169760 611322 169812 611328
rect 170036 611380 170088 611386
rect 170036 611322 170088 611328
rect 128360 610632 128412 610638
rect 128360 610574 128412 610580
rect 118790 603936 118846 603945
rect 118620 603894 118790 603922
rect 118620 603809 118648 603894
rect 118790 603871 118846 603880
rect 118606 603800 118662 603809
rect 118606 603735 118662 603744
rect 108488 603696 108540 603702
rect 108488 603638 108540 603644
rect 104820 602410 104940 602426
rect 104808 602404 104940 602410
rect 104860 602398 104940 602404
rect 104808 602346 104860 602352
rect 104900 602336 104952 602342
rect 104900 602278 104952 602284
rect 104912 601905 104940 602278
rect 104898 601896 104954 601905
rect 108500 601868 108528 603638
rect 125784 603628 125836 603634
rect 125784 603570 125836 603576
rect 111064 603560 111116 603566
rect 111064 603502 111116 603508
rect 111076 601868 111104 603502
rect 121000 602132 121052 602138
rect 121000 602074 121052 602080
rect 121012 601868 121040 602074
rect 125796 601868 125824 603570
rect 128372 601868 128400 610574
rect 169772 607918 169800 611322
rect 169760 607912 169812 607918
rect 169760 607854 169812 607860
rect 155592 607368 155644 607374
rect 155592 607310 155644 607316
rect 145656 605124 145708 605130
rect 145656 605066 145708 605072
rect 138294 604616 138350 604625
rect 138294 604551 138350 604560
rect 138110 603936 138166 603945
rect 138110 603871 138166 603880
rect 137926 603800 137982 603809
rect 138124 603786 138152 603871
rect 137982 603758 138152 603786
rect 137926 603735 137982 603744
rect 133328 602540 133380 602546
rect 133328 602482 133380 602488
rect 133340 601868 133368 602482
rect 135720 602200 135772 602206
rect 135720 602142 135772 602148
rect 135732 601868 135760 602142
rect 138308 601868 138336 604551
rect 140688 604512 140740 604518
rect 140688 604454 140740 604460
rect 140700 601868 140728 604454
rect 143080 602268 143132 602274
rect 143080 602210 143132 602216
rect 143092 601868 143120 602210
rect 145668 601868 145696 605066
rect 153016 604580 153068 604586
rect 153016 604522 153068 604528
rect 149610 603936 149666 603945
rect 149666 603894 149744 603922
rect 149610 603871 149666 603880
rect 149716 603809 149744 603894
rect 149702 603800 149758 603809
rect 149702 603735 149758 603744
rect 148048 603696 148100 603702
rect 148048 603638 148100 603644
rect 148060 601868 148088 603638
rect 150624 603356 150676 603362
rect 150624 603298 150676 603304
rect 150636 601868 150664 603298
rect 153028 601868 153056 604522
rect 155604 601868 155632 607310
rect 165344 606144 165396 606150
rect 165344 606086 165396 606092
rect 160376 605056 160428 605062
rect 160376 604998 160428 605004
rect 157982 604752 158038 604761
rect 157982 604687 158038 604696
rect 157996 601868 158024 604687
rect 160388 601868 160416 604998
rect 165356 601868 165384 606086
rect 167920 606076 167972 606082
rect 167920 606018 167972 606024
rect 167932 601868 167960 606018
rect 168288 606008 168340 606014
rect 168286 605976 168288 605985
rect 168340 605976 168342 605985
rect 168286 605911 168342 605920
rect 172888 604580 172940 604586
rect 172888 604522 172940 604528
rect 170310 603528 170366 603537
rect 170310 603463 170366 603472
rect 170324 601868 170352 603463
rect 172900 601868 172928 604522
rect 175280 603356 175332 603362
rect 175280 603298 175332 603304
rect 175292 601868 175320 603298
rect 177960 601882 177988 650014
rect 180248 607300 180300 607306
rect 180248 607242 180300 607248
rect 177698 601854 177988 601882
rect 180260 601868 180288 607242
rect 204904 607232 204956 607238
rect 204904 607174 204956 607180
rect 190184 606552 190236 606558
rect 190184 606494 190236 606500
rect 185214 605976 185270 605985
rect 185214 605911 185270 605920
rect 185228 601868 185256 605911
rect 190090 604888 190146 604897
rect 190090 604823 190146 604832
rect 190104 603770 190132 604823
rect 190092 603764 190144 603770
rect 190092 603706 190144 603712
rect 190196 601868 190224 606494
rect 199936 606212 199988 606218
rect 199936 606154 199988 606160
rect 192576 605260 192628 605266
rect 192576 605202 192628 605208
rect 192588 601868 192616 605202
rect 196070 604072 196126 604081
rect 196070 604007 196126 604016
rect 195886 603800 195942 603809
rect 196084 603786 196112 604007
rect 195942 603758 196112 603786
rect 195886 603735 195942 603744
rect 197544 603492 197596 603498
rect 197544 603434 197596 603440
rect 197556 601868 197584 603434
rect 199948 601868 199976 606154
rect 202512 603424 202564 603430
rect 202512 603366 202564 603372
rect 202524 601868 202552 603366
rect 204916 601868 204944 607174
rect 224776 606484 224828 606490
rect 224776 606426 224828 606432
rect 209872 606212 209924 606218
rect 209872 606154 209924 606160
rect 209884 601868 209912 606154
rect 219806 606112 219862 606121
rect 219806 606047 219862 606056
rect 212262 603528 212318 603537
rect 212262 603463 212318 603472
rect 212276 601868 212304 603463
rect 219820 601868 219848 606047
rect 222200 604988 222252 604994
rect 222200 604930 222252 604936
rect 222212 601868 222240 604930
rect 224788 601868 224816 606426
rect 244464 606416 244516 606422
rect 244464 606358 244516 606364
rect 242072 604648 242124 604654
rect 242072 604590 242124 604596
rect 239496 602676 239548 602682
rect 239496 602618 239548 602624
rect 232136 602608 232188 602614
rect 232136 602550 232188 602556
rect 226892 602064 226944 602070
rect 226892 602006 226944 602012
rect 226904 601882 226932 602006
rect 226904 601854 227194 601882
rect 229586 601866 229968 601882
rect 232148 601868 232176 602550
rect 237288 601928 237340 601934
rect 237130 601876 237288 601882
rect 237130 601870 237340 601876
rect 229586 601860 229980 601866
rect 229586 601854 229928 601860
rect 104898 601831 104954 601840
rect 237130 601854 237328 601870
rect 239508 601868 239536 602618
rect 242084 601868 242112 604590
rect 244476 601868 244504 606358
rect 246856 605328 246908 605334
rect 246856 605270 246908 605276
rect 246868 601868 246896 605270
rect 256792 604852 256844 604858
rect 256792 604794 256844 604800
rect 256804 601868 256832 604794
rect 259380 601868 259408 698906
rect 298756 607918 298784 700470
rect 300136 698970 300164 703520
rect 332520 700534 332548 703520
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 348804 700466 348832 703520
rect 364996 700466 365024 703520
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 397472 699990 397500 703520
rect 413664 700398 413692 703520
rect 429856 703474 429884 703520
rect 429856 703446 429976 703474
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 397460 699984 397512 699990
rect 397460 699926 397512 699932
rect 398748 699984 398800 699990
rect 398748 699926 398800 699932
rect 300124 698964 300176 698970
rect 300124 698906 300176 698912
rect 398760 628590 398788 699926
rect 429948 692850 429976 703446
rect 462332 700330 462360 703520
rect 478524 703474 478552 703520
rect 478524 703446 478644 703474
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 478616 692850 478644 703446
rect 494808 700369 494836 703520
rect 520464 700528 520516 700534
rect 520464 700470 520516 700476
rect 509976 700460 510028 700466
rect 509976 700402 510028 700408
rect 494794 700360 494850 700369
rect 494794 700295 494850 700304
rect 502340 697604 502392 697610
rect 502340 697546 502392 697552
rect 429200 692844 429252 692850
rect 429200 692786 429252 692792
rect 429936 692844 429988 692850
rect 429936 692786 429988 692792
rect 477500 692844 477552 692850
rect 477500 692786 477552 692792
rect 478604 692844 478656 692850
rect 478604 692786 478656 692792
rect 429212 673470 429240 692786
rect 477512 683074 477540 692786
rect 477512 683046 477724 683074
rect 477696 673538 477724 683046
rect 477500 673532 477552 673538
rect 477500 673474 477552 673480
rect 477684 673532 477736 673538
rect 477684 673474 477736 673480
rect 429200 673464 429252 673470
rect 429200 673406 429252 673412
rect 429476 673464 429528 673470
rect 429476 673406 429528 673412
rect 429488 647290 429516 673406
rect 477512 663762 477540 673474
rect 477512 663734 477724 663762
rect 477696 654158 477724 663734
rect 477500 654152 477552 654158
rect 477500 654094 477552 654100
rect 477684 654152 477736 654158
rect 477684 654094 477736 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 477512 644450 477540 654094
rect 477512 644422 477724 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 477696 634846 477724 644422
rect 477500 634840 477552 634846
rect 477500 634782 477552 634788
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 398748 628584 398800 628590
rect 398748 628526 398800 628532
rect 429396 621058 429424 630550
rect 477512 625138 477540 634782
rect 501604 628584 501656 628590
rect 501604 628526 501656 628532
rect 477512 625110 477724 625138
rect 429396 621030 429516 621058
rect 398840 616140 398892 616146
rect 398840 616082 398892 616088
rect 382280 614780 382332 614786
rect 382280 614722 382332 614728
rect 380440 608728 380492 608734
rect 380440 608670 380492 608676
rect 313648 608660 313700 608666
rect 313648 608602 313700 608608
rect 375472 608660 375524 608666
rect 375472 608602 375524 608608
rect 298744 607912 298796 607918
rect 298744 607854 298796 607860
rect 293958 607472 294014 607481
rect 293958 607407 294014 607416
rect 281446 607336 281502 607345
rect 281446 607271 281502 607280
rect 276664 604920 276716 604926
rect 276664 604862 276716 604868
rect 261760 603288 261812 603294
rect 261760 603230 261812 603236
rect 261772 601868 261800 603230
rect 269488 602064 269540 602070
rect 269488 602006 269540 602012
rect 263876 601996 263928 602002
rect 263876 601938 263928 601944
rect 263888 601882 263916 601938
rect 267094 601896 267150 601905
rect 263888 601854 264178 601882
rect 266754 601854 267094 601882
rect 269500 601882 269528 602006
rect 269146 601854 269528 601882
rect 276676 601868 276704 604862
rect 281460 601868 281488 607271
rect 289820 604104 289872 604110
rect 289818 604072 289820 604081
rect 289872 604072 289874 604081
rect 289818 604007 289874 604016
rect 286414 602168 286470 602177
rect 286414 602103 286470 602112
rect 288990 602168 289046 602177
rect 288990 602103 289046 602112
rect 286428 601868 286456 602103
rect 289004 601868 289032 602103
rect 293972 601868 294000 607407
rect 298742 604888 298798 604897
rect 298742 604823 298798 604832
rect 298756 601868 298784 604823
rect 309152 604166 309272 604194
rect 299388 604104 299440 604110
rect 309152 604081 309180 604166
rect 299388 604046 299440 604052
rect 309138 604072 309194 604081
rect 299400 603809 299428 604046
rect 309138 604007 309194 604016
rect 299386 603800 299442 603809
rect 299386 603735 299442 603744
rect 309244 603702 309272 604166
rect 309232 603696 309284 603702
rect 309232 603638 309284 603644
rect 303712 603220 303764 603226
rect 303712 603162 303764 603168
rect 311256 603220 311308 603226
rect 311256 603162 311308 603168
rect 301320 603152 301372 603158
rect 301320 603094 301372 603100
rect 301332 601868 301360 603094
rect 303724 601868 303752 603162
rect 309048 601996 309100 602002
rect 309048 601938 309100 601944
rect 309060 601882 309088 601938
rect 308706 601854 309088 601882
rect 311268 601868 311296 603162
rect 313660 601868 313688 608602
rect 338304 607912 338356 607918
rect 338304 607854 338356 607860
rect 330942 607608 330998 607617
rect 330942 607543 330998 607552
rect 328552 606484 328604 606490
rect 328552 606426 328604 606432
rect 318616 606348 318668 606354
rect 318616 606290 318668 606296
rect 315946 602032 316002 602041
rect 315946 601967 316002 601976
rect 315960 601882 315988 601967
rect 315960 601854 316066 601882
rect 318628 601868 318656 606290
rect 323584 606280 323636 606286
rect 323584 606222 323636 606228
rect 318706 603800 318762 603809
rect 318706 603735 318762 603744
rect 318720 603702 318748 603735
rect 318708 603696 318760 603702
rect 318708 603638 318760 603644
rect 321008 603560 321060 603566
rect 321008 603502 321060 603508
rect 318800 603356 318852 603362
rect 318800 603298 318852 603304
rect 318812 602313 318840 603298
rect 318798 602304 318854 602313
rect 318798 602239 318854 602248
rect 321020 601868 321048 603502
rect 323596 601868 323624 606222
rect 325976 604784 326028 604790
rect 325976 604726 326028 604732
rect 325988 601868 326016 604726
rect 328460 604104 328512 604110
rect 328458 604072 328460 604081
rect 328512 604072 328514 604081
rect 328458 604007 328514 604016
rect 328564 601868 328592 606426
rect 330956 601868 330984 607543
rect 335910 606248 335966 606257
rect 335910 606183 335966 606192
rect 333336 604784 333388 604790
rect 333336 604726 333388 604732
rect 333348 601868 333376 604726
rect 335924 601868 335952 606183
rect 338028 604104 338080 604110
rect 338028 604046 338080 604052
rect 338040 603809 338068 604046
rect 338026 603800 338082 603809
rect 338026 603735 338082 603744
rect 338316 601868 338344 607854
rect 372896 607368 372948 607374
rect 372896 607310 372948 607316
rect 353208 607300 353260 607306
rect 353208 607242 353260 607248
rect 340880 607232 340932 607238
rect 340880 607174 340932 607180
rect 340892 601868 340920 607174
rect 347780 604104 347832 604110
rect 347778 604072 347780 604081
rect 347832 604072 347834 604081
rect 347778 604007 347834 604016
rect 345848 603968 345900 603974
rect 345848 603910 345900 603916
rect 343272 603288 343324 603294
rect 343272 603230 343324 603236
rect 343284 601868 343312 603230
rect 345860 601868 345888 603910
rect 350630 603664 350686 603673
rect 350630 603599 350686 603608
rect 346400 603152 346452 603158
rect 346400 603094 346452 603100
rect 346412 602449 346440 603094
rect 346398 602440 346454 602449
rect 346398 602375 346454 602384
rect 350644 601868 350672 603599
rect 351828 603492 351880 603498
rect 351828 603434 351880 603440
rect 351840 603090 351868 603434
rect 351828 603084 351880 603090
rect 351828 603026 351880 603032
rect 353220 601868 353248 607242
rect 360568 605192 360620 605198
rect 360568 605134 360620 605140
rect 358176 604716 358228 604722
rect 358176 604658 358228 604664
rect 357348 604104 357400 604110
rect 357348 604046 357400 604052
rect 357360 603945 357388 604046
rect 357346 603936 357402 603945
rect 357346 603871 357402 603880
rect 358188 601868 358216 604658
rect 360580 601868 360608 605134
rect 363144 603900 363196 603906
rect 363144 603842 363196 603848
rect 363156 601868 363184 603842
rect 369674 603800 369730 603809
rect 369950 603800 370006 603809
rect 369730 603758 369950 603786
rect 369674 603735 369730 603744
rect 369950 603735 370006 603744
rect 370504 602132 370556 602138
rect 370504 602074 370556 602080
rect 370516 601868 370544 602074
rect 372908 601868 372936 607310
rect 375484 601868 375512 608602
rect 379426 603800 379482 603809
rect 379426 603735 379482 603744
rect 379440 603650 379468 603735
rect 379610 603664 379666 603673
rect 379440 603622 379610 603650
rect 379610 603599 379666 603608
rect 377864 602200 377916 602206
rect 377864 602142 377916 602148
rect 377876 601868 377904 602142
rect 380452 601868 380480 608670
rect 381452 603560 381504 603566
rect 381452 603502 381504 603508
rect 381464 602410 381492 603502
rect 381452 602404 381504 602410
rect 381452 602346 381504 602352
rect 382292 602154 382320 614722
rect 397734 606520 397790 606529
rect 397734 606455 397790 606464
rect 385222 606384 385278 606393
rect 385222 606319 385278 606328
rect 382292 602126 382596 602154
rect 382568 601882 382596 602126
rect 382568 601854 382858 601882
rect 385236 601868 385264 606319
rect 390192 606280 390244 606286
rect 390192 606222 390244 606228
rect 387800 604852 387852 604858
rect 387800 604794 387852 604800
rect 387812 601868 387840 604794
rect 390204 601868 390232 606222
rect 392766 605024 392822 605033
rect 392766 604959 392822 604968
rect 392780 601868 392808 604959
rect 395160 603152 395212 603158
rect 395160 603094 395212 603100
rect 395172 601868 395200 603094
rect 397748 601868 397776 606455
rect 398852 604194 398880 616082
rect 429488 611386 429516 621030
rect 477696 617574 477724 625110
rect 501616 620922 501644 628526
rect 501616 620894 501736 620922
rect 477684 617568 477736 617574
rect 477684 617510 477736 617516
rect 501708 611402 501736 620894
rect 429200 611380 429252 611386
rect 429200 611322 429252 611328
rect 429476 611380 429528 611386
rect 501708 611374 501828 611402
rect 429476 611322 429528 611328
rect 429212 606490 429240 611322
rect 501800 608598 501828 611374
rect 501788 608592 501840 608598
rect 501788 608534 501840 608540
rect 501972 608592 502024 608598
rect 501972 608534 502024 608540
rect 461952 606620 462004 606626
rect 461952 606562 462004 606568
rect 429200 606484 429252 606490
rect 429200 606426 429252 606432
rect 456984 606076 457036 606082
rect 456984 606018 457036 606024
rect 444656 605056 444708 605062
rect 444656 604998 444708 605004
rect 419816 604988 419868 604994
rect 419816 604930 419868 604936
rect 412456 604920 412508 604926
rect 412456 604862 412508 604868
rect 398852 604166 399892 604194
rect 399864 601882 399892 604166
rect 410064 603832 410116 603838
rect 410064 603774 410116 603780
rect 407488 603152 407540 603158
rect 407488 603094 407540 603100
rect 399864 601854 400154 601882
rect 407500 601868 407528 603094
rect 410076 601868 410104 603774
rect 412468 601868 412496 604862
rect 417424 603764 417476 603770
rect 417424 603706 417476 603712
rect 417436 601868 417464 603706
rect 419828 601868 419856 604930
rect 439686 604208 439742 604217
rect 439686 604143 439742 604152
rect 422392 603628 422444 603634
rect 422392 603570 422444 603576
rect 422404 601868 422432 603570
rect 432328 603560 432380 603566
rect 432328 603502 432380 603508
rect 429750 603392 429806 603401
rect 429750 603327 429806 603336
rect 429764 601868 429792 603327
rect 432340 601868 432368 603502
rect 439700 601868 439728 604143
rect 444472 603764 444524 603770
rect 444472 603706 444524 603712
rect 444378 603664 444434 603673
rect 444378 603599 444434 603608
rect 444392 603514 444420 603599
rect 444484 603514 444512 603706
rect 444392 603486 444512 603514
rect 442078 603392 442134 603401
rect 442078 603327 442134 603336
rect 442092 601868 442120 603327
rect 444668 601868 444696 604998
rect 452016 603832 452068 603838
rect 449162 603800 449218 603809
rect 452016 603774 452068 603780
rect 449162 603735 449164 603744
rect 449216 603735 449218 603744
rect 449164 603706 449216 603712
rect 447046 603256 447102 603265
rect 447046 603191 447102 603200
rect 449622 603256 449678 603265
rect 449622 603191 449678 603200
rect 447060 601868 447088 603191
rect 449636 601868 449664 603191
rect 452028 601868 452056 603774
rect 454408 603764 454460 603770
rect 454408 603706 454460 603712
rect 454420 601868 454448 603706
rect 456996 601868 457024 606018
rect 461964 601868 461992 606562
rect 471704 606348 471756 606354
rect 471704 606290 471756 606296
rect 463606 604208 463662 604217
rect 463606 604143 463662 604152
rect 463620 603945 463648 604143
rect 463606 603936 463662 603945
rect 463606 603871 463662 603880
rect 469312 603696 469364 603702
rect 469312 603638 469364 603644
rect 466920 603492 466972 603498
rect 466920 603434 466972 603440
rect 464344 602336 464396 602342
rect 464344 602278 464396 602284
rect 464356 601868 464384 602278
rect 466932 601868 466960 603434
rect 469324 601868 469352 603638
rect 471716 601868 471744 606290
rect 488998 604072 489054 604081
rect 488998 604007 489054 604016
rect 483018 603936 483074 603945
rect 481732 603900 481784 603906
rect 483018 603871 483020 603880
rect 481732 603842 481784 603848
rect 483072 603871 483074 603880
rect 483020 603842 483072 603848
rect 473266 603800 473322 603809
rect 473266 603735 473322 603744
rect 473280 603673 473308 603735
rect 479248 603696 479300 603702
rect 473266 603664 473322 603673
rect 479248 603638 479300 603644
rect 473266 603599 473322 603608
rect 474280 602268 474332 602274
rect 474280 602210 474332 602216
rect 474292 601868 474320 602210
rect 479260 601868 479288 603638
rect 481640 603424 481692 603430
rect 481640 603366 481692 603372
rect 481652 601868 481680 603366
rect 481744 602478 481772 603842
rect 484216 603492 484268 603498
rect 484216 603434 484268 603440
rect 481732 602472 481784 602478
rect 481732 602414 481784 602420
rect 481824 602064 481876 602070
rect 481822 602032 481824 602041
rect 481876 602032 481878 602041
rect 481822 601967 481878 601976
rect 484228 601868 484256 603434
rect 489012 601868 489040 604007
rect 492680 603968 492732 603974
rect 492680 603910 492732 603916
rect 492770 603936 492826 603945
rect 491574 603392 491630 603401
rect 491574 603327 491630 603336
rect 491588 601868 491616 603327
rect 492692 602818 492720 603910
rect 492770 603871 492772 603880
rect 492824 603871 492826 603880
rect 492772 603842 492824 603848
rect 493968 603356 494020 603362
rect 493968 603298 494020 603304
rect 492680 602812 492732 602818
rect 492680 602754 492732 602760
rect 493980 601868 494008 603298
rect 498934 603120 498990 603129
rect 498934 603055 498990 603064
rect 498200 602812 498252 602818
rect 498200 602754 498252 602760
rect 267094 601831 267150 601840
rect 229928 601802 229980 601808
rect 115940 601792 115992 601798
rect 459560 601792 459612 601798
rect 367650 601760 367706 601769
rect 115992 601740 116058 601746
rect 115940 601734 116058 601740
rect 115952 601718 116058 601734
rect 118450 601730 118648 601746
rect 118450 601724 118660 601730
rect 118450 601718 118608 601724
rect 427726 601760 427782 601769
rect 367706 601718 367954 601746
rect 427386 601718 427726 601746
rect 367650 601695 367706 601704
rect 459402 601740 459560 601746
rect 459402 601734 459612 601740
rect 459402 601718 459600 601734
rect 427726 601695 427782 601704
rect 118608 601666 118660 601672
rect 162858 601352 162914 601361
rect 105832 601322 106122 601338
rect 113192 601322 113482 601338
rect 123128 601322 123418 601338
rect 92386 601287 92442 601296
rect 97908 601316 97960 601322
rect 91100 601258 91152 601264
rect 97908 601258 97960 601264
rect 105820 601316 106122 601322
rect 105872 601310 106122 601316
rect 113180 601316 113482 601322
rect 105820 601258 105872 601264
rect 113232 601310 113482 601316
rect 123116 601316 123418 601322
rect 113180 601258 113232 601264
rect 123168 601310 123418 601316
rect 130778 601322 131068 601338
rect 130778 601316 131080 601322
rect 130778 601310 131028 601316
rect 123116 601258 123168 601264
rect 195334 601352 195390 601361
rect 162914 601310 162978 601338
rect 182666 601322 183048 601338
rect 187344 601322 187634 601338
rect 182666 601316 183060 601322
rect 182666 601310 183008 601316
rect 162858 601287 162914 601296
rect 131028 601258 131080 601264
rect 183008 601258 183060 601264
rect 187332 601316 187634 601322
rect 187384 601310 187634 601316
rect 194994 601310 195334 601338
rect 195334 601287 195390 601296
rect 207202 601352 207258 601361
rect 249706 601352 249762 601361
rect 207258 601310 207506 601338
rect 214866 601322 215064 601338
rect 217258 601322 217640 601338
rect 234264 601322 234554 601338
rect 214866 601316 215076 601322
rect 214866 601310 215024 601316
rect 207202 601287 207258 601296
rect 187332 601258 187384 601264
rect 217258 601316 217652 601322
rect 217258 601310 217600 601316
rect 215024 601258 215076 601264
rect 217600 601258 217652 601264
rect 234252 601316 234554 601322
rect 234304 601310 234554 601316
rect 249458 601310 249706 601338
rect 278778 601352 278834 601361
rect 254228 601322 254426 601338
rect 271432 601322 271722 601338
rect 249706 601287 249762 601296
rect 254216 601316 254426 601322
rect 234252 601258 234304 601264
rect 254268 601310 254426 601316
rect 271420 601316 271722 601322
rect 254216 601258 254268 601264
rect 271472 601310 271722 601316
rect 274114 601322 274496 601338
rect 274114 601316 274508 601322
rect 274114 601310 274456 601316
rect 271420 601258 271472 601264
rect 296074 601352 296130 601361
rect 278834 601310 279082 601338
rect 283760 601322 284050 601338
rect 291212 601322 291410 601338
rect 283748 601316 284050 601322
rect 278778 601287 278834 601296
rect 274456 601258 274508 601264
rect 283800 601310 284050 601316
rect 291200 601316 291410 601322
rect 283748 601258 283800 601264
rect 291252 601310 291410 601316
rect 306010 601352 306066 601361
rect 296130 601310 296378 601338
rect 296074 601287 296130 601296
rect 402886 601352 402942 601361
rect 306066 601310 306314 601338
rect 347976 601322 348266 601338
rect 347964 601316 348266 601322
rect 306010 601287 306066 601296
rect 291200 601258 291252 601264
rect 348016 601310 348266 601316
rect 355626 601322 355916 601338
rect 365562 601322 365760 601338
rect 355626 601316 355928 601322
rect 355626 601310 355876 601316
rect 347964 601258 348016 601264
rect 365562 601316 365772 601322
rect 365562 601310 365720 601316
rect 355876 601258 355928 601264
rect 402546 601310 402886 601338
rect 405462 601352 405518 601361
rect 405122 601310 405462 601338
rect 402886 601287 402942 601296
rect 415398 601352 415454 601361
rect 415058 601310 415398 601338
rect 405462 601287 405518 601296
rect 435086 601352 435142 601361
rect 424810 601322 425192 601338
rect 424810 601316 425204 601322
rect 424810 601310 425152 601316
rect 415398 601287 415454 601296
rect 365720 601258 365772 601264
rect 434746 601310 435086 601338
rect 476946 601352 477002 601361
rect 437138 601322 437336 601338
rect 437138 601316 437348 601322
rect 437138 601310 437296 601316
rect 435086 601287 435142 601296
rect 425152 601258 425204 601264
rect 476698 601310 476946 601338
rect 476946 601287 477002 601296
rect 486330 601352 486386 601361
rect 496266 601352 496322 601361
rect 486386 601310 486634 601338
rect 486330 601287 486386 601296
rect 496322 601310 496570 601338
rect 498212 601322 498240 602754
rect 498948 601868 498976 603055
rect 498200 601316 498252 601322
rect 496266 601287 496322 601296
rect 437296 601258 437348 601264
rect 501354 601310 501736 601338
rect 498200 601258 498252 601264
rect 83648 601112 83700 601118
rect 83648 601054 83700 601060
rect 83648 600500 83700 600506
rect 83648 600442 83700 600448
rect 82832 506246 83596 506274
rect 82832 499202 82860 506246
rect 83660 501922 83688 600442
rect 501512 600296 501564 600302
rect 501510 600264 501512 600273
rect 501564 600264 501566 600273
rect 501510 600199 501566 600208
rect 501708 599690 501736 601310
rect 501696 599684 501748 599690
rect 501696 599626 501748 599632
rect 501510 589520 501566 589529
rect 501510 589455 501566 589464
rect 501524 556170 501552 589455
rect 501984 574122 502012 608534
rect 502064 603832 502116 603838
rect 502064 603774 502116 603780
rect 502076 598262 502104 603774
rect 502248 603696 502300 603702
rect 502248 603638 502300 603644
rect 502064 598256 502116 598262
rect 502064 598198 502116 598204
rect 502260 596834 502288 603638
rect 502248 596828 502300 596834
rect 502248 596770 502300 596776
rect 501696 574116 501748 574122
rect 501696 574058 501748 574064
rect 501972 574116 502024 574122
rect 501972 574058 502024 574064
rect 501512 556164 501564 556170
rect 501512 556106 501564 556112
rect 501512 556028 501564 556034
rect 501512 555970 501564 555976
rect 82924 501894 83688 501922
rect 82924 501770 82952 501894
rect 82912 501764 82964 501770
rect 82912 501706 82964 501712
rect 82912 501628 82964 501634
rect 82912 501570 82964 501576
rect 82924 501514 82952 501570
rect 82924 501486 83596 501514
rect 82832 499174 83228 499202
rect 83200 493218 83228 499174
rect 82924 493190 83228 493218
rect 82924 474858 82952 493190
rect 83568 488594 83596 501486
rect 83568 488566 83688 488594
rect 83660 474994 83688 488566
rect 83016 474978 83688 474994
rect 83004 474972 83688 474978
rect 83056 474966 83688 474972
rect 83004 474914 83056 474920
rect 82924 474830 83688 474858
rect 83004 469260 83056 469266
rect 83004 469202 83056 469208
rect 83016 463706 83044 469202
rect 83660 466426 83688 474830
rect 83568 466398 83688 466426
rect 83016 463678 83320 463706
rect 83292 458810 83320 463678
rect 83568 463570 83596 466398
rect 83200 458782 83320 458810
rect 83384 463542 83596 463570
rect 82634 452976 82690 452985
rect 82690 452934 83136 452962
rect 82634 452911 82690 452920
rect 83108 451194 83136 452934
rect 83200 452010 83228 458782
rect 83384 454050 83412 463542
rect 83384 454022 83596 454050
rect 83200 451982 83320 452010
rect 82832 451166 83136 451194
rect 82832 442218 82860 451166
rect 82912 448588 82964 448594
rect 83292 448576 83320 451982
rect 83568 451194 83596 454022
rect 83568 451166 83688 451194
rect 82964 448548 83320 448576
rect 82912 448530 82964 448536
rect 83660 447658 83688 451166
rect 82924 447630 83688 447658
rect 82924 444378 82952 447630
rect 82912 444372 82964 444378
rect 82912 444314 82964 444320
rect 82832 442190 83412 442218
rect 82912 441992 82964 441998
rect 82964 441940 83228 441946
rect 82912 441934 83228 441940
rect 82924 441918 83228 441934
rect 82912 441720 82964 441726
rect 82912 441662 82964 441668
rect 82924 440230 82952 441662
rect 82820 440224 82872 440230
rect 82820 440166 82872 440172
rect 82912 440224 82964 440230
rect 82912 440166 82964 440172
rect 82832 431882 82860 440166
rect 83200 432018 83228 441918
rect 83384 434738 83412 442190
rect 83384 434710 83688 434738
rect 83200 431990 83504 432018
rect 82832 431854 83044 431882
rect 83016 430574 83044 431854
rect 82820 430568 82872 430574
rect 82820 430510 82872 430516
rect 83004 430568 83056 430574
rect 83004 430510 83056 430516
rect 82832 421410 82860 430510
rect 83476 423042 83504 431990
rect 83384 423014 83504 423042
rect 83384 421818 83412 423014
rect 83660 422362 83688 434710
rect 83476 422334 83688 422362
rect 83476 421954 83504 422334
rect 83476 421926 83688 421954
rect 83384 421790 83504 421818
rect 82832 421382 83320 421410
rect 83292 419642 83320 421382
rect 83200 419614 83320 419642
rect 83200 418418 83228 419614
rect 83476 418418 83504 421790
rect 83200 418390 83320 418418
rect 83292 417330 83320 418390
rect 82924 417302 83320 417330
rect 83384 418390 83504 418418
rect 82924 407946 82952 417302
rect 83384 412672 83412 418390
rect 83384 412644 83504 412672
rect 83476 410938 83504 412644
rect 83200 410910 83504 410938
rect 83200 410394 83228 410910
rect 83200 410366 83412 410394
rect 82924 407918 83136 407946
rect 83108 405736 83136 407918
rect 83384 405770 83412 410366
rect 83384 405742 83596 405770
rect 83108 405708 83320 405736
rect 83292 404274 83320 405708
rect 83200 404246 83320 404274
rect 83200 393666 83228 404246
rect 83568 402914 83596 405742
rect 83384 402886 83596 402914
rect 83384 398834 83412 402886
rect 83292 398806 83412 398834
rect 83292 394618 83320 398806
rect 83292 394590 83412 394618
rect 83016 393638 83228 393666
rect 83016 393394 83044 393638
rect 83016 393366 83136 393394
rect 83108 388634 83136 393366
rect 83108 388606 83320 388634
rect 83292 386322 83320 388606
rect 83384 386424 83412 394590
rect 83384 386396 83596 386424
rect 82924 386306 83320 386322
rect 82912 386300 83320 386306
rect 82964 386294 83320 386300
rect 82912 386242 82964 386248
rect 83568 386186 83596 386396
rect 82924 386158 83596 386186
rect 82924 374898 82952 386158
rect 82924 374870 83412 374898
rect 82820 374808 82872 374814
rect 82872 374756 83044 374762
rect 82820 374750 83044 374756
rect 82832 374734 83044 374750
rect 83016 374626 83044 374734
rect 83016 374598 83136 374626
rect 83108 367146 83136 374598
rect 83384 369866 83412 374870
rect 83384 369838 83596 369866
rect 83108 367118 83320 367146
rect 83292 366874 83320 367118
rect 83108 366846 83320 366874
rect 83108 346338 83136 366846
rect 83568 360754 83596 369838
rect 83384 360726 83596 360754
rect 83384 348106 83412 360726
rect 83384 348078 83596 348106
rect 83108 346310 83228 346338
rect 83200 342530 83228 346310
rect 82924 342514 83228 342530
rect 82912 342508 83228 342514
rect 82964 342502 83228 342508
rect 82912 342450 82964 342456
rect 83568 342394 83596 348078
rect 82924 342366 83596 342394
rect 82924 336954 82952 342366
rect 83660 342258 83688 421926
rect 83108 342230 83688 342258
rect 83108 341578 83136 342230
rect 83108 341550 83412 341578
rect 83384 337906 83412 341550
rect 83200 337878 83412 337906
rect 83200 337090 83228 337878
rect 83200 337062 83596 337090
rect 82924 336926 83504 336954
rect 82912 336864 82964 336870
rect 82964 336812 83044 336818
rect 82912 336806 83044 336812
rect 82924 336790 83044 336806
rect 83016 328522 83044 336790
rect 83476 333282 83504 336926
rect 83384 333254 83504 333282
rect 83016 328494 83320 328522
rect 83292 323762 83320 328494
rect 82924 323734 83320 323762
rect 82924 318850 82952 323734
rect 83384 323626 83412 333254
rect 83568 331514 83596 337062
rect 83476 331486 83596 331514
rect 83476 328930 83504 331486
rect 83476 328902 83688 328930
rect 83660 328386 83688 328902
rect 83292 323598 83412 323626
rect 83568 328358 83688 328386
rect 83568 323626 83596 328358
rect 83568 323598 83688 323626
rect 83292 321314 83320 323598
rect 83292 321286 83504 321314
rect 82820 318844 82872 318850
rect 82820 318786 82872 318792
rect 82912 318844 82964 318850
rect 82912 318786 82964 318792
rect 82832 309210 82860 318786
rect 83476 318730 83504 321286
rect 83384 318702 83504 318730
rect 83384 318186 83412 318702
rect 83660 318458 83688 323598
rect 83568 318430 83688 318458
rect 83384 318158 83504 318186
rect 83476 313970 83504 318158
rect 83384 313942 83504 313970
rect 83568 313970 83596 318430
rect 83568 313942 83688 313970
rect 83384 312066 83412 313942
rect 83384 312038 83504 312066
rect 82832 309182 83320 309210
rect 83292 302410 83320 309182
rect 83016 302382 83320 302410
rect 82912 299532 82964 299538
rect 83016 299520 83044 302382
rect 83476 302002 83504 312038
rect 83384 301974 83504 302002
rect 83384 301866 83412 301974
rect 82964 299492 83044 299520
rect 83292 301838 83412 301866
rect 82912 299474 82964 299480
rect 83292 299418 83320 301838
rect 82924 299390 83320 299418
rect 82924 294778 82952 299390
rect 82912 294772 82964 294778
rect 82912 294714 82964 294720
rect 82912 294636 82964 294642
rect 82912 294578 82964 294584
rect 82924 294386 82952 294578
rect 82924 294358 83504 294386
rect 82912 294296 82964 294302
rect 82912 294238 82964 294244
rect 82924 292482 82952 294238
rect 82924 292454 83136 292482
rect 83108 273986 83136 292454
rect 82832 273958 83136 273986
rect 82832 272354 82860 273958
rect 83476 273850 83504 294358
rect 82924 273834 83504 273850
rect 82912 273828 83504 273834
rect 82964 273822 83504 273828
rect 82912 273770 82964 273776
rect 82832 272326 83228 272354
rect 83200 260930 83228 272326
rect 83660 270042 83688 313942
rect 83384 270014 83688 270042
rect 83384 265690 83412 270014
rect 83384 265662 83504 265690
rect 83200 260902 83412 260930
rect 82924 259486 82952 259517
rect 82912 259480 82964 259486
rect 82832 259428 82912 259434
rect 82832 259422 82964 259428
rect 82832 259418 82952 259422
rect 82820 259412 82952 259418
rect 82872 259406 82952 259412
rect 82820 259354 82872 259360
rect 82912 259208 82964 259214
rect 82912 259150 82964 259156
rect 82924 246106 82952 259150
rect 83384 253042 83412 260902
rect 83476 254674 83504 265662
rect 83476 254646 83688 254674
rect 83384 253014 83504 253042
rect 83476 249778 83504 253014
rect 83292 249750 83504 249778
rect 83292 248554 83320 249750
rect 83292 248526 83504 248554
rect 82924 246078 83228 246106
rect 83200 232098 83228 246078
rect 83476 236722 83504 248526
rect 83476 236694 83596 236722
rect 83200 232070 83320 232098
rect 83292 231962 83320 232070
rect 83292 231934 83504 231962
rect 83476 219586 83504 231934
rect 82924 219570 83504 219586
rect 82912 219564 83504 219570
rect 82964 219558 83504 219564
rect 82912 219506 82964 219512
rect 83568 219450 83596 236694
rect 82924 219422 83596 219450
rect 82924 219026 82952 219422
rect 82912 219020 82964 219026
rect 82912 218962 82964 218968
rect 83660 217546 83688 254646
rect 82924 217518 83688 217546
rect 82924 210730 82952 217518
rect 83004 217456 83056 217462
rect 83056 217404 83688 217410
rect 83004 217398 83688 217404
rect 83016 217382 83688 217398
rect 83660 210746 83688 217382
rect 82912 210724 82964 210730
rect 82912 210666 82964 210672
rect 83108 210718 83688 210746
rect 83108 210610 83136 210718
rect 82924 210582 83136 210610
rect 82924 209982 82952 210582
rect 82912 209976 82964 209982
rect 82912 209918 82964 209924
rect 82912 209840 82964 209846
rect 82912 209782 82964 209788
rect 82924 208026 82952 209782
rect 82924 207998 83688 208026
rect 82924 207738 83136 207754
rect 82912 207732 83136 207738
rect 82964 207726 83136 207732
rect 82912 207674 82964 207680
rect 82912 207528 82964 207534
rect 82912 207470 82964 207476
rect 82924 195294 82952 207470
rect 83108 207074 83136 207726
rect 83108 207046 83320 207074
rect 82912 195288 82964 195294
rect 82912 195230 82964 195236
rect 83292 193066 83320 207046
rect 83292 193038 83596 193066
rect 83568 187218 83596 193038
rect 82832 187190 83596 187218
rect 82832 182866 82860 187190
rect 83660 186946 83688 207998
rect 82924 186918 83688 186946
rect 82924 182986 82952 186918
rect 82912 182980 82964 182986
rect 82912 182922 82964 182928
rect 82832 182838 83044 182866
rect 82912 182776 82964 182782
rect 82912 182718 82964 182724
rect 82268 178152 82320 178158
rect 82268 178094 82320 178100
rect 82634 175400 82690 175409
rect 82690 175358 82860 175386
rect 82634 175335 82690 175344
rect 82832 172530 82860 175358
rect 82924 173534 82952 182718
rect 83016 179058 83044 182838
rect 83016 179030 83136 179058
rect 83108 173754 83136 179030
rect 83108 173726 83228 173754
rect 82912 173528 82964 173534
rect 83200 173482 83228 173726
rect 82912 173470 82964 173476
rect 83108 173454 83228 173482
rect 82912 173392 82964 173398
rect 83108 173346 83136 173454
rect 82964 173340 83136 173346
rect 82912 173334 83136 173340
rect 82924 173318 83136 173334
rect 82832 172502 83044 172530
rect 83016 172394 83044 172502
rect 82832 172366 83044 172394
rect 82832 158710 82860 172366
rect 82912 172304 82964 172310
rect 82964 172252 83044 172258
rect 82912 172246 83044 172252
rect 82924 172230 83044 172246
rect 83016 171850 83044 172230
rect 83016 171822 83688 171850
rect 82820 158704 82872 158710
rect 82820 158646 82872 158652
rect 83660 158556 83688 171822
rect 82832 158528 83688 158556
rect 82832 157894 82860 158528
rect 82912 158432 82964 158438
rect 82964 158380 83412 158386
rect 82912 158374 83412 158380
rect 82924 158358 83412 158374
rect 82912 158024 82964 158030
rect 82912 157966 82964 157972
rect 83384 157978 83412 158358
rect 82820 157888 82872 157894
rect 82820 157830 82872 157836
rect 82728 157412 82780 157418
rect 82728 157354 82780 157360
rect 82082 155207 82138 155216
rect 82176 155236 82228 155242
rect 82176 155178 82228 155184
rect 82740 149138 82768 157354
rect 82924 155224 82952 157966
rect 83384 157950 83688 157978
rect 82924 155196 83596 155224
rect 83568 149138 83596 155196
rect 82740 149110 83044 149138
rect 83016 148322 83044 149110
rect 83476 149110 83596 149138
rect 83476 148730 83504 149110
rect 82924 148306 83044 148322
rect 82912 148300 83044 148306
rect 82964 148294 83044 148300
rect 83200 148702 83504 148730
rect 82912 148242 82964 148248
rect 83200 148186 83228 148702
rect 82924 148158 83228 148186
rect 82924 145246 82952 148158
rect 82912 145240 82964 145246
rect 82912 145182 82964 145188
rect 82924 145042 83504 145058
rect 82912 145036 83504 145042
rect 82964 145030 83504 145036
rect 82912 144978 82964 144984
rect 83476 144922 83504 145030
rect 83660 144922 83688 157950
rect 82820 144900 82872 144906
rect 83476 144894 83688 144922
rect 82820 144842 82872 144848
rect 82832 140282 82860 144842
rect 82912 144832 82964 144838
rect 82912 144774 82964 144780
rect 82924 144106 82952 144774
rect 82924 144078 83136 144106
rect 83108 143970 83136 144078
rect 83108 143942 83320 143970
rect 82912 143744 82964 143750
rect 82964 143692 83136 143698
rect 82912 143686 83136 143692
rect 82924 143670 83136 143686
rect 82912 143608 82964 143614
rect 82964 143556 83044 143562
rect 82912 143550 83044 143556
rect 82924 143534 83044 143550
rect 82820 140276 82872 140282
rect 82820 140218 82872 140224
rect 83016 140162 83044 143534
rect 82832 140134 83044 140162
rect 82542 138816 82598 138825
rect 82542 138751 82598 138760
rect 82556 132530 82584 138751
rect 82832 137306 82860 140134
rect 82912 140072 82964 140078
rect 83108 140060 83136 143670
rect 83292 143562 83320 143942
rect 83292 143534 83412 143562
rect 82964 140032 83136 140060
rect 82912 140014 82964 140020
rect 83384 138666 83412 143534
rect 83384 138638 83688 138666
rect 82740 137278 82860 137306
rect 82634 135008 82690 135017
rect 82634 134943 82690 134952
rect 82648 134774 82676 134943
rect 82636 134768 82688 134774
rect 82636 134710 82688 134716
rect 82544 132524 82596 132530
rect 82544 132466 82596 132472
rect 82174 120592 82230 120601
rect 82174 120527 82230 120536
rect 81900 120080 81952 120086
rect 81900 120022 81952 120028
rect 81990 117056 82046 117065
rect 81990 116991 82046 117000
rect 82004 101930 82032 116991
rect 81992 101924 82044 101930
rect 81992 101866 82044 101872
rect 82188 101318 82216 120527
rect 82636 106752 82688 106758
rect 82634 106720 82636 106729
rect 82688 106720 82690 106729
rect 82634 106655 82690 106664
rect 82740 102814 82768 137278
rect 82820 137216 82872 137222
rect 82820 137158 82872 137164
rect 82832 132546 82860 137158
rect 82912 134768 82964 134774
rect 82964 134716 83412 134722
rect 82912 134710 83412 134716
rect 82924 134694 83412 134710
rect 82924 132790 83320 132818
rect 82924 132666 82952 132790
rect 82912 132660 82964 132666
rect 82912 132602 82964 132608
rect 82832 132518 83044 132546
rect 83016 129146 83044 132518
rect 82832 129118 83044 129146
rect 82832 123978 82860 129118
rect 83292 128602 83320 132790
rect 83384 132512 83412 134694
rect 83384 132484 83504 132512
rect 83476 128602 83504 132484
rect 83292 128574 83412 128602
rect 83476 128574 83596 128602
rect 83384 124386 83412 128574
rect 83200 124358 83412 124386
rect 83200 124250 83228 124358
rect 82924 124234 83228 124250
rect 82912 124228 83228 124234
rect 82964 124222 83228 124228
rect 82912 124170 82964 124176
rect 82924 124098 83320 124114
rect 82912 124092 83320 124098
rect 82964 124086 83320 124092
rect 82912 124034 82964 124040
rect 83292 123978 83320 124086
rect 83568 123978 83596 128574
rect 82832 123950 83228 123978
rect 83292 123950 83596 123978
rect 83200 123026 83228 123950
rect 83108 122998 83228 123026
rect 82912 118720 82964 118726
rect 82912 118662 82964 118668
rect 82924 115258 82952 118662
rect 82912 115252 82964 115258
rect 82912 115194 82964 115200
rect 83108 115138 83136 122998
rect 83108 115110 83320 115138
rect 83292 111466 83320 115110
rect 83292 111438 83412 111466
rect 83384 111058 83412 111438
rect 82912 111036 82964 111042
rect 83384 111030 83504 111058
rect 82912 110978 82964 110984
rect 82924 110922 82952 110978
rect 82924 110894 83136 110922
rect 82912 106752 82964 106758
rect 82964 106700 83044 106706
rect 82912 106694 83044 106700
rect 82924 106678 83044 106694
rect 83016 104854 83044 106678
rect 83004 104848 83056 104854
rect 83004 104790 83056 104796
rect 82912 104780 82964 104786
rect 82912 104722 82964 104728
rect 82728 102808 82780 102814
rect 82728 102750 82780 102756
rect 82176 101312 82228 101318
rect 82176 101254 82228 101260
rect 82556 100570 82584 102068
rect 82544 100564 82596 100570
rect 82544 100506 82596 100512
rect 82924 99634 82952 104722
rect 83108 102474 83136 110894
rect 83476 105346 83504 111030
rect 83660 106978 83688 138638
rect 501524 137873 501552 555970
rect 501708 554878 501736 574058
rect 501696 554872 501748 554878
rect 501696 554814 501748 554820
rect 501604 554804 501656 554810
rect 501604 554746 501656 554752
rect 501616 536858 501644 554746
rect 501604 536852 501656 536858
rect 501604 536794 501656 536800
rect 501696 536716 501748 536722
rect 501696 536658 501748 536664
rect 501708 524498 501736 536658
rect 502352 535401 502380 697546
rect 502432 667956 502484 667962
rect 502432 667898 502484 667904
rect 502338 535392 502394 535401
rect 502338 535327 502394 535336
rect 501786 526416 501842 526425
rect 501786 526351 501842 526360
rect 501616 524470 501736 524498
rect 501616 524362 501644 524470
rect 501616 524334 501736 524362
rect 501708 520266 501736 524334
rect 501800 522889 501828 526351
rect 501878 524784 501934 524793
rect 501878 524719 501934 524728
rect 501786 522880 501842 522889
rect 501786 522815 501842 522824
rect 501892 522345 501920 524719
rect 501878 522336 501934 522345
rect 501878 522271 501934 522280
rect 501696 520260 501748 520266
rect 501696 520202 501748 520208
rect 501604 510672 501656 510678
rect 501604 510614 501656 510620
rect 501616 507822 501644 510614
rect 501604 507816 501656 507822
rect 501604 507758 501656 507764
rect 502062 507784 502118 507793
rect 502062 507719 502118 507728
rect 502076 498409 502104 507719
rect 502062 498400 502118 498409
rect 502062 498335 502118 498344
rect 501696 498228 501748 498234
rect 501696 498170 501748 498176
rect 501708 480282 501736 498170
rect 501970 481536 502026 481545
rect 501970 481471 502026 481480
rect 501604 480276 501656 480282
rect 501604 480218 501656 480224
rect 501696 480276 501748 480282
rect 501696 480218 501748 480224
rect 501616 467838 501644 480218
rect 501984 472025 502012 481471
rect 501970 472016 502026 472025
rect 501970 471951 502026 471960
rect 502062 471880 502118 471889
rect 502062 471815 502118 471824
rect 501604 467832 501656 467838
rect 501604 467774 501656 467780
rect 501696 467832 501748 467838
rect 501696 467774 501748 467780
rect 501708 449954 501736 467774
rect 502076 462641 502104 471815
rect 502062 462632 502118 462641
rect 502062 462567 502118 462576
rect 501970 458960 502026 458969
rect 501970 458895 502026 458904
rect 501984 452713 502012 458895
rect 501970 452704 502026 452713
rect 501970 452639 502026 452648
rect 502338 451344 502394 451353
rect 502338 451279 502394 451288
rect 501604 449948 501656 449954
rect 501604 449890 501656 449896
rect 501696 449948 501748 449954
rect 501696 449890 501748 449896
rect 501616 448526 501644 449890
rect 501604 448520 501656 448526
rect 501604 448462 501656 448468
rect 501696 448520 501748 448526
rect 501696 448462 501748 448468
rect 501708 430681 501736 448462
rect 502062 442912 502118 442921
rect 502062 442847 502118 442856
rect 502076 433401 502104 442847
rect 502062 433392 502118 433401
rect 502062 433327 502118 433336
rect 501694 430672 501750 430681
rect 501694 430607 501750 430616
rect 501878 430536 501934 430545
rect 501878 430471 501934 430480
rect 501892 420968 501920 430471
rect 502062 428496 502118 428505
rect 502062 428431 502118 428440
rect 502076 423706 502104 428431
rect 501972 423700 502024 423706
rect 501972 423642 502024 423648
rect 502064 423700 502116 423706
rect 502064 423642 502116 423648
rect 501800 420940 501920 420968
rect 501800 411330 501828 420940
rect 501984 415449 502012 423642
rect 501970 415440 502026 415449
rect 501970 415375 502026 415384
rect 502062 413944 502118 413953
rect 502062 413879 502118 413888
rect 501604 411324 501656 411330
rect 501604 411266 501656 411272
rect 501788 411324 501840 411330
rect 501788 411266 501840 411272
rect 501616 405226 501644 411266
rect 501616 405198 501828 405226
rect 501800 391950 501828 405198
rect 502076 404569 502104 413879
rect 502062 404560 502118 404569
rect 502062 404495 502118 404504
rect 502062 394632 502118 394641
rect 502062 394567 502118 394576
rect 501696 391944 501748 391950
rect 501696 391886 501748 391892
rect 501788 391944 501840 391950
rect 501788 391886 501840 391892
rect 501708 376718 501736 391886
rect 502076 385257 502104 394567
rect 502062 385248 502118 385257
rect 502062 385183 502118 385192
rect 501696 376712 501748 376718
rect 501696 376654 501748 376660
rect 501788 376712 501840 376718
rect 501788 376654 501840 376660
rect 501800 358834 501828 376654
rect 502062 360904 502118 360913
rect 502062 360839 502118 360848
rect 501696 358828 501748 358834
rect 501696 358770 501748 358776
rect 501788 358828 501840 358834
rect 501788 358770 501840 358776
rect 501708 357406 501736 358770
rect 501604 357400 501656 357406
rect 501604 357342 501656 357348
rect 501696 357400 501748 357406
rect 501696 357342 501748 357348
rect 501616 339454 501644 357342
rect 502076 356153 502104 360839
rect 502062 356144 502118 356153
rect 502062 356079 502118 356088
rect 502246 354648 502302 354657
rect 502246 354583 502302 354592
rect 502260 345273 502288 354583
rect 502246 345264 502302 345273
rect 502246 345199 502302 345208
rect 501604 339448 501656 339454
rect 501604 339390 501656 339396
rect 501696 339448 501748 339454
rect 501696 339390 501748 339396
rect 501708 327593 501736 339390
rect 502062 335336 502118 335345
rect 502062 335271 502118 335280
rect 501694 327584 501750 327593
rect 501694 327519 501750 327528
rect 502076 325825 502104 335271
rect 502062 325816 502118 325825
rect 502062 325751 502118 325760
rect 501602 321464 501658 321473
rect 501602 321399 501658 321408
rect 501616 312089 501644 321399
rect 501602 312080 501658 312089
rect 501602 312015 501658 312024
rect 501602 308272 501658 308281
rect 501602 308207 501658 308216
rect 501510 137864 501566 137873
rect 501510 137799 501566 137808
rect 501510 136640 501566 136649
rect 501510 136575 501566 136584
rect 83292 105318 83504 105346
rect 83568 106950 83688 106978
rect 83292 104394 83320 105318
rect 83568 105074 83596 106950
rect 83476 105046 83596 105074
rect 83476 104768 83504 105046
rect 83476 104740 83688 104768
rect 83660 104394 83688 104740
rect 83292 104366 83504 104394
rect 83096 102468 83148 102474
rect 83096 102410 83148 102416
rect 83372 102332 83424 102338
rect 83372 102274 83424 102280
rect 82924 99606 83136 99634
rect 81900 97436 81952 97442
rect 81900 97378 81952 97384
rect 81808 22772 81860 22778
rect 81808 22714 81860 22720
rect 81912 3398 81940 97378
rect 83108 94586 83136 99606
rect 83384 95946 83412 102274
rect 83372 95940 83424 95946
rect 83372 95882 83424 95888
rect 83476 94722 83504 104366
rect 83568 104366 83688 104394
rect 83568 100094 83596 104366
rect 133892 102734 134012 102762
rect 133892 102649 133920 102734
rect 108946 102640 109002 102649
rect 109130 102640 109186 102649
rect 109002 102598 109130 102626
rect 108946 102575 109002 102584
rect 109130 102575 109186 102584
rect 118422 102640 118478 102649
rect 118606 102640 118662 102649
rect 118478 102598 118606 102626
rect 118422 102575 118478 102584
rect 118606 102575 118662 102584
rect 125506 102640 125562 102649
rect 125506 102575 125562 102584
rect 133694 102640 133750 102649
rect 133694 102575 133750 102584
rect 133878 102640 133934 102649
rect 133878 102575 133934 102584
rect 125520 102542 125548 102575
rect 133708 102542 133736 102575
rect 125508 102536 125560 102542
rect 84014 102504 84070 102513
rect 83648 102468 83700 102474
rect 125508 102478 125560 102484
rect 133696 102536 133748 102542
rect 133984 102513 134012 102734
rect 201500 102740 201552 102746
rect 201500 102682 201552 102688
rect 176750 102640 176806 102649
rect 173992 102604 174044 102610
rect 173992 102546 174044 102552
rect 176672 102598 176750 102626
rect 133696 102478 133748 102484
rect 133970 102504 134026 102513
rect 84014 102439 84070 102448
rect 149072 102474 149178 102490
rect 133970 102439 134026 102448
rect 149060 102468 149178 102474
rect 83648 102410 83700 102416
rect 83660 101862 83688 102410
rect 83648 101856 83700 101862
rect 83648 101798 83700 101804
rect 83556 100088 83608 100094
rect 83556 100030 83608 100036
rect 83464 94716 83516 94722
rect 83464 94658 83516 94664
rect 83096 94580 83148 94586
rect 83096 94522 83148 94528
rect 83464 94580 83516 94586
rect 83464 94522 83516 94528
rect 83280 89412 83332 89418
rect 83280 89354 83332 89360
rect 83292 84946 83320 89354
rect 83476 85082 83504 94522
rect 83476 85054 83688 85082
rect 83292 84918 83596 84946
rect 83568 77330 83596 84918
rect 83476 77302 83596 77330
rect 83476 67674 83504 77302
rect 83660 70514 83688 85054
rect 84028 72486 84056 102439
rect 149112 102462 149178 102468
rect 149060 102410 149112 102416
rect 84844 102400 84896 102406
rect 84844 102342 84896 102348
rect 84106 75168 84162 75177
rect 84106 75103 84162 75112
rect 84016 72480 84068 72486
rect 84016 72422 84068 72428
rect 83648 70508 83700 70514
rect 83648 70450 83700 70456
rect 83648 70372 83700 70378
rect 83648 70314 83700 70320
rect 83384 67646 83504 67674
rect 83384 66230 83412 67646
rect 83372 66224 83424 66230
rect 83372 66166 83424 66172
rect 83556 57860 83608 57866
rect 83556 57802 83608 57808
rect 83568 51082 83596 57802
rect 83660 57254 83688 70314
rect 83648 57248 83700 57254
rect 83648 57190 83700 57196
rect 83384 51054 83596 51082
rect 83384 46306 83412 51054
rect 83372 46300 83424 46306
rect 83372 46242 83424 46248
rect 84120 3482 84148 75103
rect 84856 4078 84884 102342
rect 151570 102190 151768 102218
rect 88338 102096 88394 102105
rect 84962 102054 85528 102082
rect 84936 100564 84988 100570
rect 84936 100506 84988 100512
rect 84948 87650 84976 100506
rect 84936 87644 84988 87650
rect 84936 87586 84988 87592
rect 85500 76634 85528 102054
rect 85578 101960 85634 101969
rect 85578 101895 85634 101904
rect 85592 101454 85620 101895
rect 85580 101448 85632 101454
rect 85580 101390 85632 101396
rect 85580 101312 85632 101318
rect 85580 101254 85632 101260
rect 85488 76628 85540 76634
rect 85488 76570 85540 76576
rect 85488 18624 85540 18630
rect 85488 18566 85540 18572
rect 84844 4072 84896 4078
rect 84844 4014 84896 4020
rect 83844 3454 84148 3482
rect 81900 3392 81952 3398
rect 81900 3334 81952 3340
rect 82636 3392 82688 3398
rect 82636 3334 82688 3340
rect 82648 480 82676 3334
rect 83844 480 83872 3454
rect 85500 3058 85528 18566
rect 85592 3482 85620 101254
rect 87340 100473 87368 102068
rect 88338 102031 88394 102040
rect 88352 100910 88380 102031
rect 88524 101720 88576 101726
rect 88524 101662 88576 101668
rect 88340 100904 88392 100910
rect 88340 100846 88392 100852
rect 88536 100722 88564 101662
rect 88352 100694 88564 100722
rect 87326 100464 87382 100473
rect 87326 100399 87382 100408
rect 88248 64184 88300 64190
rect 88248 64126 88300 64132
rect 85592 3454 86172 3482
rect 84936 3052 84988 3058
rect 84936 2994 84988 3000
rect 85488 3052 85540 3058
rect 85488 2994 85540 3000
rect 84948 480 84976 2994
rect 86144 480 86172 3454
rect 88260 3398 88288 64126
rect 87328 3392 87380 3398
rect 87328 3334 87380 3340
rect 88248 3392 88300 3398
rect 88352 3380 88380 100694
rect 89916 100162 89944 102068
rect 91112 102054 92322 102082
rect 94898 102054 95188 102082
rect 97290 102054 97948 102082
rect 89994 101688 90050 101697
rect 89994 101623 90050 101632
rect 89904 100156 89956 100162
rect 89904 100098 89956 100104
rect 90008 89706 90036 101623
rect 91008 100156 91060 100162
rect 91008 100098 91060 100104
rect 89916 89678 90036 89706
rect 89916 82142 89944 89678
rect 89904 82136 89956 82142
rect 89904 82078 89956 82084
rect 90088 82136 90140 82142
rect 90088 82078 90140 82084
rect 90100 77353 90128 82078
rect 89902 77344 89958 77353
rect 89824 77302 89902 77330
rect 89824 77194 89852 77302
rect 89902 77279 89958 77288
rect 90086 77344 90142 77353
rect 90086 77279 90142 77288
rect 89824 77166 89944 77194
rect 89916 70446 89944 77166
rect 89904 70440 89956 70446
rect 89904 70382 89956 70388
rect 89812 70236 89864 70242
rect 89812 70178 89864 70184
rect 89824 60790 89852 70178
rect 89812 60784 89864 60790
rect 89812 60726 89864 60732
rect 89996 60716 90048 60722
rect 89996 60658 90048 60664
rect 90008 57934 90036 60658
rect 89996 57928 90048 57934
rect 89996 57870 90048 57876
rect 89904 48340 89956 48346
rect 89904 48282 89956 48288
rect 89916 41426 89944 48282
rect 90916 47592 90968 47598
rect 90916 47534 90968 47540
rect 89824 41410 89944 41426
rect 89812 41404 89944 41410
rect 89864 41398 89944 41404
rect 89996 41404 90048 41410
rect 89812 41346 89864 41352
rect 89996 41346 90048 41352
rect 90008 31822 90036 41346
rect 89996 31816 90048 31822
rect 89996 31758 90048 31764
rect 89904 29096 89956 29102
rect 89824 29044 89904 29050
rect 89824 29038 89956 29044
rect 89824 29022 89944 29038
rect 89824 27606 89852 29022
rect 89812 27600 89864 27606
rect 89812 27542 89864 27548
rect 89996 21956 90048 21962
rect 89996 21898 90048 21904
rect 89720 3392 89772 3398
rect 88352 3352 88564 3380
rect 88248 3334 88300 3340
rect 87340 480 87368 3334
rect 88536 480 88564 3352
rect 89720 3334 89772 3340
rect 89732 480 89760 3334
rect 90008 3262 90036 21898
rect 90928 3398 90956 47534
rect 91020 17270 91048 100098
rect 91112 25566 91140 102054
rect 93952 101788 94004 101794
rect 93952 101730 94004 101736
rect 93768 71052 93820 71058
rect 93768 70994 93820 71000
rect 91100 25560 91152 25566
rect 91100 25502 91152 25508
rect 91008 17264 91060 17270
rect 91008 17206 91060 17212
rect 92388 14952 92440 14958
rect 92388 14894 92440 14900
rect 90916 3392 90968 3398
rect 92400 3380 92428 14894
rect 93780 3398 93808 70994
rect 93964 3398 93992 101730
rect 95160 21418 95188 102054
rect 96528 68332 96580 68338
rect 96528 68274 96580 68280
rect 95148 21412 95200 21418
rect 95148 21354 95200 21360
rect 96540 3398 96568 68274
rect 97920 60042 97948 102054
rect 99668 100162 99696 102068
rect 99656 100156 99708 100162
rect 99656 100098 99708 100104
rect 100668 100156 100720 100162
rect 100668 100098 100720 100104
rect 99472 100088 99524 100094
rect 99472 100030 99524 100036
rect 99288 61396 99340 61402
rect 99288 61338 99340 61344
rect 97908 60036 97960 60042
rect 97908 59978 97960 59984
rect 99194 26888 99250 26897
rect 99194 26823 99250 26832
rect 97908 25764 97960 25770
rect 97908 25706 97960 25712
rect 97920 3398 97948 25706
rect 99208 3482 99236 26823
rect 99300 3618 99328 61338
rect 99300 3590 99420 3618
rect 99208 3454 99328 3482
rect 90916 3334 90968 3340
rect 92124 3352 92428 3380
rect 93308 3392 93360 3398
rect 89996 3256 90048 3262
rect 89996 3198 90048 3204
rect 90916 3256 90968 3262
rect 90916 3198 90968 3204
rect 90928 480 90956 3198
rect 92124 480 92152 3352
rect 93308 3334 93360 3340
rect 93768 3392 93820 3398
rect 93768 3334 93820 3340
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 94504 3392 94556 3398
rect 94504 3334 94556 3340
rect 95700 3392 95752 3398
rect 95700 3334 95752 3340
rect 96528 3392 96580 3398
rect 96528 3334 96580 3340
rect 96896 3392 96948 3398
rect 96896 3334 96948 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 98092 3392 98144 3398
rect 98092 3334 98144 3340
rect 93320 480 93348 3334
rect 94516 480 94544 3334
rect 95712 480 95740 3334
rect 96908 480 96936 3334
rect 98104 480 98132 3334
rect 99300 480 99328 3454
rect 99392 3398 99420 3590
rect 99380 3392 99432 3398
rect 99380 3334 99432 3340
rect 99484 610 99512 100030
rect 100680 25634 100708 100098
rect 102244 99890 102272 102068
rect 104650 102054 104848 102082
rect 107226 102054 107516 102082
rect 109618 102054 110368 102082
rect 103612 101652 103664 101658
rect 103612 101594 103664 101600
rect 102232 99884 102284 99890
rect 102232 99826 102284 99832
rect 103428 99884 103480 99890
rect 103428 99826 103480 99832
rect 102048 84856 102100 84862
rect 102048 84798 102100 84804
rect 100668 25628 100720 25634
rect 100668 25570 100720 25576
rect 102060 3398 102088 84798
rect 103440 44946 103468 99826
rect 103428 44940 103480 44946
rect 103428 44882 103480 44888
rect 103428 28416 103480 28422
rect 103428 28358 103480 28364
rect 103440 3398 103468 28358
rect 103624 3482 103652 101594
rect 104820 40730 104848 102054
rect 106464 101924 106516 101930
rect 106464 101866 106516 101872
rect 106188 65544 106240 65550
rect 106188 65486 106240 65492
rect 104808 40724 104860 40730
rect 104808 40666 104860 40672
rect 103624 3454 104020 3482
rect 101588 3392 101640 3398
rect 101588 3334 101640 3340
rect 102048 3392 102100 3398
rect 102048 3334 102100 3340
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 99472 604 99524 610
rect 99472 546 99524 552
rect 100484 604 100536 610
rect 100484 546 100536 552
rect 100496 480 100524 546
rect 101600 480 101628 3334
rect 102796 480 102824 3334
rect 103992 480 104020 3454
rect 106200 3398 106228 65486
rect 105176 3392 105228 3398
rect 105176 3334 105228 3340
rect 106188 3392 106240 3398
rect 106188 3334 106240 3340
rect 106372 3392 106424 3398
rect 106476 3380 106504 101866
rect 107488 61538 107516 102054
rect 107660 101856 107712 101862
rect 107660 101798 107712 101804
rect 107568 73976 107620 73982
rect 107568 73918 107620 73924
rect 107476 61532 107528 61538
rect 107476 61474 107528 61480
rect 107580 3618 107608 73918
rect 107672 3754 107700 101798
rect 110236 43512 110288 43518
rect 110236 43454 110288 43460
rect 107672 3726 108804 3754
rect 107580 3590 107700 3618
rect 107672 3398 107700 3590
rect 107660 3392 107712 3398
rect 106476 3352 107608 3380
rect 106372 3334 106424 3340
rect 105188 480 105216 3334
rect 106384 480 106412 3334
rect 107580 480 107608 3352
rect 107660 3334 107712 3340
rect 108776 480 108804 3726
rect 110248 3482 110276 43454
rect 110340 25566 110368 102054
rect 112180 100230 112208 102068
rect 114572 100230 114600 102068
rect 116978 102054 117268 102082
rect 119554 102054 120028 102082
rect 116122 101552 116178 101561
rect 116122 101487 116178 101496
rect 112168 100224 112220 100230
rect 112168 100166 112220 100172
rect 114560 100224 114612 100230
rect 114560 100166 114612 100172
rect 115848 100224 115900 100230
rect 115848 100166 115900 100172
rect 110420 100020 110472 100026
rect 110420 99962 110472 99968
rect 110328 25560 110380 25566
rect 110328 25502 110380 25508
rect 109972 3454 110276 3482
rect 110432 3482 110460 99962
rect 115754 50280 115810 50289
rect 115754 50215 115810 50224
rect 113548 9376 113600 9382
rect 113548 9318 113600 9324
rect 112352 4820 112404 4826
rect 112352 4762 112404 4768
rect 110432 3454 111196 3482
rect 109972 480 110000 3454
rect 111168 480 111196 3454
rect 112364 480 112392 4762
rect 113560 480 113588 9318
rect 115768 3398 115796 50215
rect 115860 16046 115888 100166
rect 115848 16040 115900 16046
rect 115848 15982 115900 15988
rect 114744 3392 114796 3398
rect 114744 3334 114796 3340
rect 115756 3392 115808 3398
rect 115756 3334 115808 3340
rect 114756 480 114784 3334
rect 116136 626 116164 101487
rect 117240 18766 117268 102054
rect 117320 101584 117372 101590
rect 117320 101526 117372 101532
rect 117228 18760 117280 18766
rect 117228 18702 117280 18708
rect 117136 7608 117188 7614
rect 117136 7550 117188 7556
rect 115952 598 116164 626
rect 115952 480 115980 598
rect 117148 480 117176 7550
rect 117332 3398 117360 101526
rect 117964 100156 118016 100162
rect 117964 100098 118016 100104
rect 117976 19990 118004 100098
rect 120000 75206 120028 102054
rect 121932 99754 121960 102068
rect 124508 100609 124536 102068
rect 124494 100600 124550 100609
rect 124494 100535 124550 100544
rect 126900 100230 126928 102068
rect 128360 101516 128412 101522
rect 128360 101458 128412 101464
rect 124864 100224 124916 100230
rect 124864 100166 124916 100172
rect 126888 100224 126940 100230
rect 126888 100166 126940 100172
rect 121920 99748 121972 99754
rect 121920 99690 121972 99696
rect 122748 99748 122800 99754
rect 122748 99690 122800 99696
rect 120078 98968 120134 98977
rect 120078 98903 120134 98912
rect 119988 75200 120040 75206
rect 119988 75142 120040 75148
rect 119988 66904 120040 66910
rect 119988 66846 120040 66852
rect 117964 19984 118016 19990
rect 117964 19926 118016 19932
rect 120000 3398 120028 66846
rect 117320 3392 117372 3398
rect 117320 3334 117372 3340
rect 118240 3392 118292 3398
rect 118240 3334 118292 3340
rect 119436 3392 119488 3398
rect 119436 3334 119488 3340
rect 119988 3392 120040 3398
rect 119988 3334 120040 3340
rect 118252 480 118280 3334
rect 119448 480 119476 3334
rect 120092 610 120120 98903
rect 122760 19990 122788 99690
rect 122840 93288 122892 93294
rect 122840 93230 122892 93236
rect 122748 19984 122800 19990
rect 122748 19926 122800 19932
rect 121828 9648 121880 9654
rect 121828 9590 121880 9596
rect 120080 604 120132 610
rect 120080 546 120132 552
rect 120632 604 120684 610
rect 120632 546 120684 552
rect 120644 480 120672 546
rect 121840 480 121868 9590
rect 122852 3482 122880 93230
rect 124876 13122 124904 100166
rect 128268 68468 128320 68474
rect 128268 68410 128320 68416
rect 125508 17332 125560 17338
rect 125508 17274 125560 17280
rect 124864 13116 124916 13122
rect 124864 13058 124916 13064
rect 125416 6656 125468 6662
rect 125416 6598 125468 6604
rect 122852 3454 123064 3482
rect 123036 480 123064 3454
rect 124220 3392 124272 3398
rect 124220 3334 124272 3340
rect 124232 480 124260 3334
rect 125428 480 125456 6598
rect 125520 3398 125548 17274
rect 126888 13116 126940 13122
rect 126888 13058 126940 13064
rect 126900 3482 126928 13058
rect 126624 3454 126928 3482
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 126624 480 126652 3454
rect 128280 3398 128308 68410
rect 127808 3392 127860 3398
rect 127808 3334 127860 3340
rect 128268 3392 128320 3398
rect 128268 3334 128320 3340
rect 127820 480 127848 3334
rect 128372 610 128400 101458
rect 129476 97986 129504 102068
rect 131210 101416 131266 101425
rect 131210 101351 131266 101360
rect 129738 98696 129794 98705
rect 129738 98631 129794 98640
rect 129464 97980 129516 97986
rect 129464 97922 129516 97928
rect 129752 3398 129780 98631
rect 131224 3482 131252 101351
rect 131868 100298 131896 102068
rect 133892 102054 134274 102082
rect 131856 100292 131908 100298
rect 131856 100234 131908 100240
rect 131764 100020 131816 100026
rect 131764 99962 131816 99968
rect 131776 55894 131804 99962
rect 132592 99272 132644 99278
rect 132592 99214 132644 99220
rect 131764 55888 131816 55894
rect 131764 55830 131816 55836
rect 131224 3454 131436 3482
rect 129740 3392 129792 3398
rect 129740 3334 129792 3340
rect 130200 3392 130252 3398
rect 130200 3334 130252 3340
rect 128360 604 128412 610
rect 128360 546 128412 552
rect 129004 604 129056 610
rect 129004 546 129056 552
rect 129016 480 129044 546
rect 130212 480 130240 3334
rect 131408 480 131436 3454
rect 132604 480 132632 99214
rect 133892 73982 133920 102054
rect 136836 100298 136864 102068
rect 136824 100292 136876 100298
rect 136824 100234 136876 100240
rect 137928 100292 137980 100298
rect 137928 100234 137980 100240
rect 135166 79384 135222 79393
rect 135166 79319 135222 79328
rect 133880 73976 133932 73982
rect 133880 73918 133932 73924
rect 133696 4208 133748 4214
rect 133696 4150 133748 4156
rect 133708 2825 133736 4150
rect 133788 4140 133840 4146
rect 133788 4082 133840 4088
rect 133694 2816 133750 2825
rect 133694 2751 133750 2760
rect 133800 480 133828 4082
rect 135180 3380 135208 79319
rect 136548 55888 136600 55894
rect 136548 55830 136600 55836
rect 135258 5808 135314 5817
rect 135258 5743 135260 5752
rect 135312 5743 135314 5752
rect 135260 5714 135312 5720
rect 136560 3398 136588 55830
rect 137940 28354 137968 100234
rect 139228 100026 139256 102068
rect 141804 100745 141832 102068
rect 144210 102054 144868 102082
rect 141790 100736 141846 100745
rect 141790 100671 141846 100680
rect 142804 100088 142856 100094
rect 142804 100030 142856 100036
rect 139216 100020 139268 100026
rect 139216 99962 139268 99968
rect 142160 99204 142212 99210
rect 142160 99146 142212 99152
rect 138020 87644 138072 87650
rect 138020 87586 138072 87592
rect 138032 87009 138060 87586
rect 138018 87000 138074 87009
rect 138018 86935 138074 86944
rect 140778 87000 140834 87009
rect 140778 86935 140834 86944
rect 140792 77217 140820 86935
rect 140502 77208 140558 77217
rect 140502 77143 140558 77152
rect 140778 77208 140834 77217
rect 140778 77143 140834 77152
rect 140516 67697 140544 77143
rect 140502 67688 140558 67697
rect 140502 67623 140558 67632
rect 140778 67688 140834 67697
rect 140778 67623 140834 67632
rect 140792 67590 140820 67623
rect 140780 67584 140832 67590
rect 140780 67526 140832 67532
rect 140872 67584 140924 67590
rect 140872 67526 140924 67532
rect 140884 58018 140912 67526
rect 140792 57990 140912 58018
rect 140792 57934 140820 57990
rect 140688 57928 140740 57934
rect 140688 57870 140740 57876
rect 140780 57928 140832 57934
rect 140780 57870 140832 57876
rect 140700 56574 140728 57870
rect 140688 56568 140740 56574
rect 140688 56510 140740 56516
rect 140780 46980 140832 46986
rect 140780 46922 140832 46928
rect 140792 45558 140820 46922
rect 140780 45552 140832 45558
rect 140780 45494 140832 45500
rect 140686 44840 140742 44849
rect 140686 44775 140742 44784
rect 137928 28348 137980 28354
rect 137928 28290 137980 28296
rect 136640 18760 136692 18766
rect 136640 18702 136692 18708
rect 136652 3482 136680 18702
rect 138480 6656 138532 6662
rect 138480 6598 138532 6604
rect 136652 3454 137324 3482
rect 134904 3352 135208 3380
rect 136088 3392 136140 3398
rect 134904 480 134932 3352
rect 136088 3334 136140 3340
rect 136548 3392 136600 3398
rect 136548 3334 136600 3340
rect 136100 480 136128 3334
rect 137296 480 137324 3454
rect 138492 480 138520 6598
rect 140700 2922 140728 44775
rect 140872 35964 140924 35970
rect 140872 35906 140924 35912
rect 140884 29322 140912 35906
rect 140884 29294 141004 29322
rect 140976 28914 141004 29294
rect 140792 28886 141004 28914
rect 140792 27554 140820 28886
rect 140792 27526 140912 27554
rect 140884 22710 140912 27526
rect 140872 22704 140924 22710
rect 140872 22646 140924 22652
rect 142068 12436 142120 12442
rect 142068 12378 142120 12384
rect 140780 9716 140832 9722
rect 140780 9658 140832 9664
rect 140792 4842 140820 9658
rect 140792 4814 140912 4842
rect 139676 2916 139728 2922
rect 139676 2858 139728 2864
rect 140688 2916 140740 2922
rect 140688 2858 140740 2864
rect 139688 480 139716 2858
rect 140884 480 140912 4814
rect 142080 480 142108 12378
rect 142172 4078 142200 99146
rect 142816 22846 142844 100030
rect 144644 58812 144696 58818
rect 144644 58754 144696 58760
rect 144656 58018 144684 58754
rect 144656 57990 144776 58018
rect 144748 57934 144776 57990
rect 144736 57928 144788 57934
rect 144736 57870 144788 57876
rect 144736 48340 144788 48346
rect 144736 48282 144788 48288
rect 144748 38622 144776 48282
rect 144736 38616 144788 38622
rect 144736 38558 144788 38564
rect 144736 29028 144788 29034
rect 144736 28970 144788 28976
rect 142804 22840 142856 22846
rect 142804 22782 142856 22788
rect 144748 19310 144776 28970
rect 144840 28286 144868 102054
rect 146300 99068 146352 99074
rect 146300 99010 146352 99016
rect 146208 93152 146260 93158
rect 146208 93094 146260 93100
rect 144828 28280 144880 28286
rect 144828 28222 144880 28228
rect 144736 19304 144788 19310
rect 144736 19246 144788 19252
rect 144736 9716 144788 9722
rect 144736 9658 144788 9664
rect 142160 4072 142212 4078
rect 142160 4014 142212 4020
rect 143264 4072 143316 4078
rect 143264 4014 143316 4020
rect 143276 480 143304 4014
rect 144748 2854 144776 9658
rect 144828 5772 144880 5778
rect 144828 5714 144880 5720
rect 144840 5658 144868 5714
rect 145010 5672 145066 5681
rect 144840 5630 145010 5658
rect 145010 5607 145066 5616
rect 146220 4078 146248 93094
rect 146312 4078 146340 99010
rect 146772 97986 146800 102068
rect 149704 100020 149756 100026
rect 149704 99962 149756 99968
rect 149060 99136 149112 99142
rect 149060 99078 149112 99084
rect 146760 97980 146812 97986
rect 146760 97922 146812 97928
rect 148966 36544 149022 36553
rect 148966 36479 149022 36488
rect 145656 4072 145708 4078
rect 145656 4014 145708 4020
rect 146208 4072 146260 4078
rect 146208 4014 146260 4020
rect 146300 4072 146352 4078
rect 146300 4014 146352 4020
rect 146852 4072 146904 4078
rect 146852 4014 146904 4020
rect 144736 2848 144788 2854
rect 144736 2790 144788 2796
rect 144460 2780 144512 2786
rect 144460 2722 144512 2728
rect 144472 480 144500 2722
rect 145668 480 145696 4014
rect 146864 480 146892 4014
rect 148980 3398 149008 36479
rect 149072 3482 149100 99078
rect 149716 7614 149744 99962
rect 151740 96642 151768 102190
rect 151648 96614 151768 96642
rect 153212 102054 154146 102082
rect 156538 102054 157288 102082
rect 151648 87038 151676 96614
rect 151728 95940 151780 95946
rect 151728 95882 151780 95888
rect 151544 87032 151596 87038
rect 151544 86974 151596 86980
rect 151636 87032 151688 87038
rect 151636 86974 151688 86980
rect 151556 81122 151584 86974
rect 151544 81116 151596 81122
rect 151544 81058 151596 81064
rect 151544 77376 151596 77382
rect 151464 77324 151544 77330
rect 151464 77318 151596 77324
rect 151464 77302 151584 77318
rect 151464 77178 151492 77302
rect 151452 77172 151504 77178
rect 151452 77114 151504 77120
rect 151544 67652 151596 67658
rect 151544 67594 151596 67600
rect 151556 60858 151584 67594
rect 151544 60852 151596 60858
rect 151544 60794 151596 60800
rect 151452 60716 151504 60722
rect 151452 60658 151504 60664
rect 151464 51066 151492 60658
rect 151452 51060 151504 51066
rect 151452 51002 151504 51008
rect 151636 51060 151688 51066
rect 151636 51002 151688 51008
rect 151648 48278 151676 51002
rect 151636 48272 151688 48278
rect 151636 48214 151688 48220
rect 151544 38684 151596 38690
rect 151544 38626 151596 38632
rect 151556 31770 151584 38626
rect 151464 31742 151584 31770
rect 151464 26926 151492 31742
rect 151452 26920 151504 26926
rect 151452 26862 151504 26868
rect 149704 7608 149756 7614
rect 149704 7550 149756 7556
rect 150440 4004 150492 4010
rect 150440 3946 150492 3952
rect 149072 3454 149284 3482
rect 148048 3392 148100 3398
rect 148048 3334 148100 3340
rect 148968 3392 149020 3398
rect 148968 3334 149020 3340
rect 148060 480 148088 3334
rect 149256 480 149284 3454
rect 150452 480 150480 3946
rect 151740 3482 151768 95882
rect 153108 49020 153160 49026
rect 153108 48962 153160 48968
rect 153120 3482 153148 48962
rect 153212 26994 153240 102054
rect 155960 84924 156012 84930
rect 155960 84866 156012 84872
rect 155868 46232 155920 46238
rect 155868 46174 155920 46180
rect 153200 26988 153252 26994
rect 153200 26930 153252 26936
rect 153936 6860 153988 6866
rect 153936 6802 153988 6808
rect 151556 3454 151768 3482
rect 152752 3454 153148 3482
rect 151556 480 151584 3454
rect 152752 480 152780 3454
rect 153948 480 153976 6802
rect 155880 3330 155908 46174
rect 155972 3482 156000 84866
rect 157260 78062 157288 102054
rect 159100 100162 159128 102068
rect 159088 100156 159140 100162
rect 159088 100098 159140 100104
rect 161492 97889 161520 102068
rect 164068 100366 164096 102068
rect 166460 100842 166488 102068
rect 166448 100836 166500 100842
rect 166448 100778 166500 100784
rect 164056 100360 164108 100366
rect 164056 100302 164108 100308
rect 167000 99000 167052 99006
rect 167000 98942 167052 98948
rect 161478 97880 161534 97889
rect 161478 97815 161534 97824
rect 164146 95840 164202 95849
rect 164146 95775 164202 95784
rect 157248 78056 157300 78062
rect 157248 77998 157300 78004
rect 161388 38072 161440 38078
rect 161388 38014 161440 38020
rect 158628 14748 158680 14754
rect 158628 14690 158680 14696
rect 158640 4078 158668 14690
rect 159916 6792 159968 6798
rect 159916 6734 159968 6740
rect 157524 4072 157576 4078
rect 157524 4014 157576 4020
rect 158628 4072 158680 4078
rect 158628 4014 158680 4020
rect 155972 3454 156368 3482
rect 155132 3324 155184 3330
rect 155132 3266 155184 3272
rect 155868 3324 155920 3330
rect 155868 3266 155920 3272
rect 155144 480 155172 3266
rect 156340 480 156368 3454
rect 157536 480 157564 4014
rect 158720 3392 158772 3398
rect 158720 3334 158772 3340
rect 158732 480 158760 3334
rect 159928 480 159956 6734
rect 161400 2854 161428 38014
rect 162766 5944 162822 5953
rect 162766 5879 162822 5888
rect 162780 5545 162808 5879
rect 162766 5536 162822 5545
rect 163042 5536 163098 5545
rect 162766 5471 162822 5480
rect 162964 5494 163042 5522
rect 162964 5409 162992 5494
rect 163042 5471 163098 5480
rect 162950 5400 163006 5409
rect 162950 5335 163006 5344
rect 162308 3936 162360 3942
rect 162308 3878 162360 3884
rect 161112 2848 161164 2854
rect 161112 2790 161164 2796
rect 161388 2848 161440 2854
rect 161388 2790 161440 2796
rect 161124 480 161152 2790
rect 162320 480 162348 3878
rect 164160 3058 164188 95775
rect 165528 62824 165580 62830
rect 165528 62766 165580 62772
rect 165540 3058 165568 62766
rect 167012 4078 167040 98942
rect 168852 96626 168880 102068
rect 171428 100745 171456 102068
rect 173728 102054 173834 102082
rect 171414 100736 171470 100745
rect 171414 100671 171470 100680
rect 168840 96620 168892 96626
rect 168840 96562 168892 96568
rect 171140 73908 171192 73914
rect 171140 73850 171192 73856
rect 169760 19984 169812 19990
rect 169760 19926 169812 19932
rect 169772 12442 169800 19926
rect 169760 12436 169812 12442
rect 169760 12378 169812 12384
rect 170588 12436 170640 12442
rect 170588 12378 170640 12384
rect 167000 4072 167052 4078
rect 167000 4014 167052 4020
rect 168196 4072 168248 4078
rect 168196 4014 168248 4020
rect 169390 4040 169446 4049
rect 165896 3868 165948 3874
rect 165896 3810 165948 3816
rect 163504 3052 163556 3058
rect 163504 2994 163556 3000
rect 164148 3052 164200 3058
rect 164148 2994 164200 3000
rect 164700 3052 164752 3058
rect 164700 2994 164752 3000
rect 165528 3052 165580 3058
rect 165528 2994 165580 3000
rect 163516 480 163544 2994
rect 164712 480 164740 2994
rect 165908 480 165936 3810
rect 167092 3800 167144 3806
rect 167092 3742 167144 3748
rect 167104 480 167132 3742
rect 168208 480 168236 4014
rect 169390 3975 169446 3984
rect 169404 480 169432 3975
rect 170600 480 170628 12378
rect 171152 610 171180 73850
rect 173728 19990 173756 102054
rect 173808 93356 173860 93362
rect 173808 93298 173860 93304
rect 173716 19984 173768 19990
rect 173716 19926 173768 19932
rect 173820 3126 173848 93298
rect 172980 3120 173032 3126
rect 172980 3062 173032 3068
rect 173808 3120 173860 3126
rect 173808 3062 173860 3068
rect 171140 604 171192 610
rect 171140 546 171192 552
rect 171784 604 171836 610
rect 171784 546 171836 552
rect 171796 480 171824 546
rect 172992 480 173020 3062
rect 174004 626 174032 102546
rect 176396 100434 176424 102068
rect 176566 101416 176622 101425
rect 176566 101351 176622 101360
rect 176384 100428 176436 100434
rect 176384 100370 176436 100376
rect 176476 87644 176528 87650
rect 176476 87586 176528 87592
rect 175372 3324 175424 3330
rect 175372 3266 175424 3272
rect 174004 598 174216 626
rect 174188 480 174216 598
rect 175384 480 175412 3266
rect 176488 3074 176516 87586
rect 176580 3330 176608 101351
rect 176672 99362 176700 102598
rect 176750 102575 176806 102584
rect 176672 99334 176792 99362
rect 176764 96626 176792 99334
rect 178788 97850 178816 102068
rect 183756 99346 183784 102068
rect 186148 100502 186176 102068
rect 188448 102054 188738 102082
rect 187792 101856 187844 101862
rect 187792 101798 187844 101804
rect 186136 100496 186188 100502
rect 186136 100438 186188 100444
rect 186964 100156 187016 100162
rect 186964 100098 187016 100104
rect 183744 99340 183796 99346
rect 183744 99282 183796 99288
rect 184848 99340 184900 99346
rect 184848 99282 184900 99288
rect 179420 98864 179472 98870
rect 179420 98806 179472 98812
rect 178776 97844 178828 97850
rect 178776 97786 178828 97792
rect 176752 96620 176804 96626
rect 176752 96562 176804 96568
rect 176752 89684 176804 89690
rect 176752 89626 176804 89632
rect 176764 86986 176792 89626
rect 176672 86970 176792 86986
rect 176660 86964 176804 86970
rect 176712 86958 176752 86964
rect 176660 86906 176712 86912
rect 176752 86906 176804 86912
rect 176764 79914 176792 86906
rect 176764 79886 176884 79914
rect 176856 77178 176884 79886
rect 176844 77172 176896 77178
rect 176844 77114 176896 77120
rect 176752 67652 176804 67658
rect 176752 67594 176804 67600
rect 176764 60738 176792 67594
rect 176764 60710 176884 60738
rect 176856 57934 176884 60710
rect 176844 57928 176896 57934
rect 176844 57870 176896 57876
rect 176752 48340 176804 48346
rect 176752 48282 176804 48288
rect 176764 41426 176792 48282
rect 176764 41398 176884 41426
rect 176856 38622 176884 41398
rect 176844 38616 176896 38622
rect 176844 38558 176896 38564
rect 176752 31748 176804 31754
rect 176752 31690 176804 31696
rect 176764 22114 176792 31690
rect 176764 22086 176884 22114
rect 176856 19310 176884 22086
rect 176844 19304 176896 19310
rect 176844 19246 176896 19252
rect 176936 9716 176988 9722
rect 176936 9658 176988 9664
rect 176948 4078 176976 9658
rect 178960 7608 179012 7614
rect 178960 7550 179012 7556
rect 176936 4072 176988 4078
rect 176936 4014 176988 4020
rect 177764 4072 177816 4078
rect 177764 4014 177816 4020
rect 176568 3324 176620 3330
rect 176568 3266 176620 3272
rect 176488 3046 176608 3074
rect 176580 480 176608 3046
rect 177776 480 177804 4014
rect 178972 480 179000 7550
rect 179432 4078 179460 98806
rect 183468 93220 183520 93226
rect 183468 93162 183520 93168
rect 182088 32564 182140 32570
rect 182088 32506 182140 32512
rect 179420 4072 179472 4078
rect 179420 4014 179472 4020
rect 180156 4072 180208 4078
rect 180156 4014 180208 4020
rect 180168 480 180196 4014
rect 182100 2990 182128 32506
rect 182180 5704 182232 5710
rect 182178 5672 182180 5681
rect 182232 5672 182234 5681
rect 182178 5607 182234 5616
rect 183480 3330 183508 93162
rect 184860 76566 184888 99282
rect 186228 93288 186280 93294
rect 186228 93230 186280 93236
rect 184848 76560 184900 76566
rect 184848 76502 184900 76508
rect 184848 29708 184900 29714
rect 184848 29650 184900 29656
rect 183744 6724 183796 6730
rect 183744 6666 183796 6672
rect 182548 3324 182600 3330
rect 182548 3266 182600 3272
rect 183468 3324 183520 3330
rect 183468 3266 183520 3272
rect 181352 2984 181404 2990
rect 181352 2926 181404 2932
rect 182088 2984 182140 2990
rect 182088 2926 182140 2932
rect 181364 480 181392 2926
rect 182560 480 182588 3266
rect 183756 480 183784 6666
rect 184860 480 184888 29650
rect 186240 626 186268 93230
rect 186320 16040 186372 16046
rect 186320 15982 186372 15988
rect 186056 598 186268 626
rect 186332 610 186360 15982
rect 186976 14958 187004 100098
rect 187700 98048 187752 98054
rect 187700 97990 187752 97996
rect 187712 87650 187740 97990
rect 187700 87644 187752 87650
rect 187700 87586 187752 87592
rect 186964 14952 187016 14958
rect 186964 14894 187016 14900
rect 187804 3398 187832 101798
rect 188448 98054 188476 102054
rect 188436 98048 188488 98054
rect 188436 97990 188488 97996
rect 191116 96490 191144 102068
rect 193692 100881 193720 102068
rect 193678 100872 193734 100881
rect 193678 100807 193734 100816
rect 193220 98932 193272 98938
rect 193220 98874 193272 98880
rect 191104 96484 191156 96490
rect 191104 96426 191156 96432
rect 190366 46200 190422 46209
rect 190366 46135 190422 46144
rect 190380 3398 190408 46135
rect 193128 16040 193180 16046
rect 193128 15982 193180 15988
rect 190828 9580 190880 9586
rect 190828 9522 190880 9528
rect 187792 3392 187844 3398
rect 187792 3334 187844 3340
rect 188436 3392 188488 3398
rect 188436 3334 188488 3340
rect 189632 3392 189684 3398
rect 189632 3334 189684 3340
rect 190368 3392 190420 3398
rect 190368 3334 190420 3340
rect 186320 604 186372 610
rect 186056 480 186084 598
rect 186320 546 186372 552
rect 187240 604 187292 610
rect 187240 546 187292 552
rect 187252 480 187280 546
rect 188448 480 188476 3334
rect 189644 480 189672 3334
rect 190840 480 190868 9522
rect 193140 3398 193168 15982
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 192036 480 192064 3334
rect 193232 480 193260 98874
rect 195980 98796 196032 98802
rect 195980 98738 196032 98744
rect 195888 96008 195940 96014
rect 195888 95950 195940 95956
rect 194508 77988 194560 77994
rect 194508 77930 194560 77936
rect 194520 3482 194548 77930
rect 195900 3482 195928 95950
rect 194428 3454 194548 3482
rect 195624 3454 195928 3482
rect 194428 480 194456 3454
rect 195624 480 195652 3454
rect 195992 610 196020 98738
rect 196084 93362 196112 102068
rect 198660 100094 198688 102068
rect 200132 102054 201066 102082
rect 198740 101516 198792 101522
rect 198740 101458 198792 101464
rect 198648 100088 198700 100094
rect 198648 100030 198700 100036
rect 198752 96665 198780 101458
rect 198370 96656 198426 96665
rect 198370 96591 198426 96600
rect 198738 96656 198794 96665
rect 198738 96591 198794 96600
rect 196072 93356 196124 93362
rect 196072 93298 196124 93304
rect 198384 89706 198412 96591
rect 200028 93356 200080 93362
rect 200028 93298 200080 93304
rect 198384 89678 198596 89706
rect 198568 86970 198596 89678
rect 198556 86964 198608 86970
rect 198556 86906 198608 86912
rect 198464 77308 198516 77314
rect 198464 77250 198516 77256
rect 198476 77178 198504 77250
rect 198464 77172 198516 77178
rect 198464 77114 198516 77120
rect 198556 67652 198608 67658
rect 198556 67594 198608 67600
rect 198568 60858 198596 67594
rect 198556 60852 198608 60858
rect 198556 60794 198608 60800
rect 198464 60716 198516 60722
rect 198464 60658 198516 60664
rect 198476 57934 198504 60658
rect 198464 57928 198516 57934
rect 198464 57870 198516 57876
rect 198556 48340 198608 48346
rect 198556 48282 198608 48288
rect 198568 41478 198596 48282
rect 198556 41472 198608 41478
rect 198556 41414 198608 41420
rect 198464 41404 198516 41410
rect 198464 41346 198516 41352
rect 198476 38622 198504 41346
rect 198464 38616 198516 38622
rect 198464 38558 198516 38564
rect 198556 31680 198608 31686
rect 198556 31622 198608 31628
rect 198568 21978 198596 31622
rect 198568 21950 198688 21978
rect 198660 4078 198688 21950
rect 199934 5808 199990 5817
rect 199934 5743 199990 5752
rect 199948 5710 199976 5743
rect 199936 5704 199988 5710
rect 199936 5646 199988 5652
rect 200040 4078 200068 93298
rect 200132 47598 200160 102054
rect 201408 86420 201460 86426
rect 201408 86362 201460 86368
rect 200120 47592 200172 47598
rect 200120 47534 200172 47540
rect 198004 4072 198056 4078
rect 198004 4014 198056 4020
rect 198648 4072 198700 4078
rect 198648 4014 198700 4020
rect 199200 4072 199252 4078
rect 199200 4014 199252 4020
rect 200028 4072 200080 4078
rect 200028 4014 200080 4020
rect 195980 604 196032 610
rect 195980 546 196032 552
rect 196808 604 196860 610
rect 196808 546 196860 552
rect 196820 480 196848 546
rect 198016 480 198044 4014
rect 199212 480 199240 4014
rect 201420 3194 201448 86362
rect 201512 7546 201540 102682
rect 370504 102672 370556 102678
rect 307666 102640 307722 102649
rect 370504 102614 370556 102620
rect 416688 102672 416740 102678
rect 416688 102614 416740 102620
rect 307666 102575 307722 102584
rect 274546 102504 274602 102513
rect 274546 102439 274602 102448
rect 211002 102326 211200 102354
rect 203458 102054 204208 102082
rect 204076 29640 204128 29646
rect 204076 29582 204128 29588
rect 202788 16108 202840 16114
rect 202788 16050 202840 16056
rect 201500 7540 201552 7546
rect 201500 7482 201552 7488
rect 202696 7540 202748 7546
rect 202696 7482 202748 7488
rect 201592 5976 201644 5982
rect 201590 5944 201592 5953
rect 201644 5944 201646 5953
rect 201590 5879 201646 5888
rect 201500 4072 201552 4078
rect 201500 4014 201552 4020
rect 200396 3188 200448 3194
rect 200396 3130 200448 3136
rect 201408 3188 201460 3194
rect 201408 3130 201460 3136
rect 200408 480 200436 3130
rect 201512 480 201540 4014
rect 202708 480 202736 7482
rect 202800 4078 202828 16050
rect 202788 4072 202840 4078
rect 202788 4014 202840 4020
rect 204088 2854 204116 29582
rect 204180 14958 204208 102054
rect 206020 100298 206048 102068
rect 206008 100292 206060 100298
rect 206008 100234 206060 100240
rect 206928 100292 206980 100298
rect 206928 100234 206980 100240
rect 207664 100292 207716 100298
rect 207664 100234 207716 100240
rect 204260 75200 204312 75206
rect 204260 75142 204312 75148
rect 204168 14952 204220 14958
rect 204168 14894 204220 14900
rect 204272 12442 204300 75142
rect 204260 12436 204312 12442
rect 204260 12378 204312 12384
rect 205088 12436 205140 12442
rect 205088 12378 205140 12384
rect 204076 2848 204128 2854
rect 204076 2790 204128 2796
rect 203892 604 203944 610
rect 203892 546 203944 552
rect 203904 480 203932 546
rect 205100 480 205128 12378
rect 206284 9512 206336 9518
rect 206284 9454 206336 9460
rect 206296 480 206324 9454
rect 206940 4894 206968 100234
rect 207020 98660 207072 98666
rect 207020 98602 207072 98608
rect 206928 4888 206980 4894
rect 206928 4830 206980 4836
rect 207032 4078 207060 98602
rect 207676 29782 207704 100234
rect 208412 65550 208440 102068
rect 211172 96642 211200 102326
rect 212262 101552 212318 101561
rect 212262 101487 212318 101496
rect 212276 96694 212304 101487
rect 213380 100162 213408 102068
rect 215970 102054 216536 102082
rect 213368 100156 213420 100162
rect 213368 100098 213420 100104
rect 212540 97300 212592 97306
rect 212540 97242 212592 97248
rect 211080 96614 211200 96642
rect 212264 96688 212316 96694
rect 212264 96630 212316 96636
rect 212356 96688 212408 96694
rect 212408 96636 212488 96642
rect 212356 96630 212488 96636
rect 212368 96614 212488 96630
rect 209686 87680 209742 87689
rect 209686 87615 209742 87624
rect 208400 65544 208452 65550
rect 208400 65486 208452 65492
rect 207664 29776 207716 29782
rect 207664 29718 207716 29724
rect 209700 4078 209728 87615
rect 210884 83564 210936 83570
rect 210884 83506 210936 83512
rect 210896 4078 210924 83506
rect 211080 82142 211108 96614
rect 212460 96506 212488 96614
rect 212368 96478 212488 96506
rect 212368 91746 212396 96478
rect 212368 91718 212488 91746
rect 211068 82136 211120 82142
rect 211068 82078 211120 82084
rect 210976 65544 211028 65550
rect 210976 65486 211028 65492
rect 210988 48346 211016 65486
rect 212460 57934 212488 91718
rect 212448 57928 212500 57934
rect 212448 57870 212500 57876
rect 210976 48340 211028 48346
rect 210976 48282 211028 48288
rect 212448 48340 212500 48346
rect 212448 48282 212500 48288
rect 210976 46980 211028 46986
rect 210976 46922 211028 46928
rect 210988 46866 211016 46922
rect 210988 46838 211108 46866
rect 211080 37330 211108 46838
rect 210976 37324 211028 37330
rect 210976 37266 211028 37272
rect 211068 37324 211120 37330
rect 211068 37266 211120 37272
rect 210988 27606 211016 37266
rect 210976 27600 211028 27606
rect 210976 27542 211028 27548
rect 212460 19310 212488 48282
rect 211160 19304 211212 19310
rect 211160 19246 211212 19252
rect 212448 19304 212500 19310
rect 212448 19246 212500 19252
rect 211068 5976 211120 5982
rect 211066 5944 211068 5953
rect 211120 5944 211122 5953
rect 211066 5879 211122 5888
rect 211172 4876 211200 19246
rect 212552 12442 212580 97242
rect 213918 86320 213974 86329
rect 213918 86255 213974 86264
rect 213932 12442 213960 86255
rect 216508 24206 216536 102054
rect 218348 100502 218376 102068
rect 220648 102054 220754 102082
rect 223330 102054 223528 102082
rect 225722 102054 226288 102082
rect 228298 102054 229048 102082
rect 218336 100496 218388 100502
rect 218336 100438 218388 100444
rect 219348 100496 219400 100502
rect 219348 100438 219400 100444
rect 218060 98728 218112 98734
rect 218060 98670 218112 98676
rect 216588 98660 216640 98666
rect 216588 98602 216640 98608
rect 216496 24200 216548 24206
rect 216496 24142 216548 24148
rect 212540 12436 212592 12442
rect 212540 12378 212592 12384
rect 213460 12436 213512 12442
rect 213460 12378 213512 12384
rect 213920 12436 213972 12442
rect 213920 12378 213972 12384
rect 214656 12436 214708 12442
rect 214656 12378 214708 12384
rect 212448 9716 212500 9722
rect 212448 9658 212500 9664
rect 211080 4848 211200 4876
rect 207020 4072 207072 4078
rect 207020 4014 207072 4020
rect 207480 4072 207532 4078
rect 207480 4014 207532 4020
rect 208676 4072 208728 4078
rect 208676 4014 208728 4020
rect 209688 4072 209740 4078
rect 209688 4014 209740 4020
rect 209872 4072 209924 4078
rect 209872 4014 209924 4020
rect 210884 4072 210936 4078
rect 210884 4014 210936 4020
rect 207492 480 207520 4014
rect 208688 480 208716 4014
rect 209884 480 209912 4014
rect 211080 480 211108 4848
rect 212460 2854 212488 9658
rect 212448 2848 212500 2854
rect 212448 2790 212500 2796
rect 212264 2780 212316 2786
rect 212264 2722 212316 2728
rect 212276 480 212304 2722
rect 213472 480 213500 12378
rect 214668 480 214696 12378
rect 216600 3194 216628 98602
rect 217968 93424 218020 93430
rect 217968 93366 218020 93372
rect 217980 4078 218008 93366
rect 218072 4078 218100 98670
rect 219256 58676 219308 58682
rect 219256 58618 219308 58624
rect 217048 4072 217100 4078
rect 217048 4014 217100 4020
rect 217968 4072 218020 4078
rect 217968 4014 218020 4020
rect 218060 4072 218112 4078
rect 218060 4014 218112 4020
rect 215852 3188 215904 3194
rect 215852 3130 215904 3136
rect 216588 3188 216640 3194
rect 216588 3130 216640 3136
rect 215864 480 215892 3130
rect 217060 480 217088 4014
rect 219268 3262 219296 58618
rect 219360 32502 219388 100438
rect 220648 55962 220676 102054
rect 220728 93492 220780 93498
rect 220728 93434 220780 93440
rect 220636 55956 220688 55962
rect 220636 55898 220688 55904
rect 219348 32496 219400 32502
rect 219348 32438 219400 32444
rect 220634 6080 220690 6089
rect 220634 6015 220690 6024
rect 220648 5409 220676 6015
rect 220634 5400 220690 5409
rect 220634 5335 220690 5344
rect 219348 4072 219400 4078
rect 219348 4014 219400 4020
rect 218152 3256 218204 3262
rect 218152 3198 218204 3204
rect 219256 3256 219308 3262
rect 219256 3198 219308 3204
rect 218164 480 218192 3198
rect 219360 480 219388 4014
rect 220740 610 220768 93434
rect 222108 61668 222160 61674
rect 222108 61610 222160 61616
rect 222120 626 222148 61610
rect 223500 44878 223528 102054
rect 225604 100088 225656 100094
rect 225604 100030 225656 100036
rect 223488 44872 223540 44878
rect 223488 44814 223540 44820
rect 223580 32428 223632 32434
rect 223580 32370 223632 32376
rect 222936 3664 222988 3670
rect 222936 3606 222988 3612
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 221752 598 222148 626
rect 220556 480 220584 546
rect 221752 480 221780 598
rect 222948 480 222976 3606
rect 223592 610 223620 32370
rect 225616 6594 225644 100030
rect 226260 71126 226288 102054
rect 227628 98728 227680 98734
rect 227628 98670 227680 98676
rect 226248 71120 226300 71126
rect 226248 71062 226300 71068
rect 225604 6588 225656 6594
rect 225604 6530 225656 6536
rect 225328 4888 225380 4894
rect 225328 4830 225380 4836
rect 223580 604 223632 610
rect 223580 546 223632 552
rect 224132 604 224184 610
rect 224132 546 224184 552
rect 224144 480 224172 546
rect 225340 480 225368 4830
rect 227640 3398 227668 98670
rect 228916 80708 228968 80714
rect 228916 80650 228968 80656
rect 228824 38004 228876 38010
rect 228824 37946 228876 37952
rect 227720 3664 227772 3670
rect 227720 3606 227772 3612
rect 226524 3392 226576 3398
rect 226524 3334 226576 3340
rect 227628 3392 227680 3398
rect 227628 3334 227680 3340
rect 226536 480 226564 3334
rect 227732 480 227760 3606
rect 228836 3482 228864 37946
rect 228928 3670 228956 80650
rect 229020 6594 229048 102054
rect 230676 100502 230704 102068
rect 230664 100496 230716 100502
rect 230664 100438 230716 100444
rect 231768 100496 231820 100502
rect 231768 100438 231820 100444
rect 230480 78056 230532 78062
rect 230480 77998 230532 78004
rect 229100 12368 229152 12374
rect 229100 12310 229152 12316
rect 229008 6588 229060 6594
rect 229008 6530 229060 6536
rect 228916 3664 228968 3670
rect 228916 3606 228968 3612
rect 229112 3482 229140 12310
rect 230492 3482 230520 77998
rect 231780 17406 231808 100438
rect 233148 75200 233200 75206
rect 233148 75142 233200 75148
rect 231768 17400 231820 17406
rect 231768 17342 231820 17348
rect 228836 3454 228956 3482
rect 229112 3454 230152 3482
rect 230492 3454 231348 3482
rect 228928 480 228956 3454
rect 230124 480 230152 3454
rect 231320 480 231348 3454
rect 233160 3398 233188 75142
rect 233252 15978 233280 102068
rect 235658 102054 235948 102082
rect 234620 50380 234672 50386
rect 234620 50322 234672 50328
rect 233332 24200 233384 24206
rect 233332 24142 233384 24148
rect 233240 15972 233292 15978
rect 233240 15914 233292 15920
rect 232504 3392 232556 3398
rect 232504 3334 232556 3340
rect 233148 3392 233200 3398
rect 233148 3334 233200 3340
rect 233344 3346 233372 24142
rect 234632 3346 234660 50322
rect 235920 42158 235948 102054
rect 237392 102054 238050 102082
rect 237286 98696 237342 98705
rect 237286 98631 237342 98640
rect 235908 42152 235960 42158
rect 235908 42094 235960 42100
rect 237196 31068 237248 31074
rect 237196 31010 237248 31016
rect 237208 3670 237236 31010
rect 236000 3664 236052 3670
rect 236000 3606 236052 3612
rect 237196 3664 237248 3670
rect 237196 3606 237248 3612
rect 232516 480 232544 3334
rect 233344 3318 233740 3346
rect 234632 3318 234844 3346
rect 233712 480 233740 3318
rect 234816 480 234844 3318
rect 236012 480 236040 3606
rect 237300 3482 237328 98631
rect 237392 4826 237420 102054
rect 240612 100094 240640 102068
rect 245580 100842 245608 102068
rect 247986 102054 248276 102082
rect 250562 102054 251036 102082
rect 245568 100836 245620 100842
rect 245568 100778 245620 100784
rect 240784 100224 240836 100230
rect 240784 100166 240836 100172
rect 240600 100088 240652 100094
rect 240600 100030 240652 100036
rect 240048 73976 240100 73982
rect 240048 73918 240100 73924
rect 237472 46300 237524 46306
rect 237472 46242 237524 46248
rect 237380 4820 237432 4826
rect 237380 4762 237432 4768
rect 237208 3454 237328 3482
rect 237484 3482 237512 46242
rect 237484 3454 238432 3482
rect 237208 480 237236 3454
rect 238404 480 238432 3454
rect 240060 3398 240088 73918
rect 240796 62898 240824 100166
rect 241428 98796 241480 98802
rect 241428 98738 241480 98744
rect 240784 62892 240836 62898
rect 240784 62834 240836 62840
rect 241440 3398 241468 98738
rect 242806 97200 242862 97209
rect 242806 97135 242862 97144
rect 239588 3392 239640 3398
rect 239588 3334 239640 3340
rect 240048 3392 240100 3398
rect 240048 3334 240100 3340
rect 240784 3392 240836 3398
rect 240784 3334 240836 3340
rect 241428 3392 241480 3398
rect 241428 3334 241480 3340
rect 239600 480 239628 3334
rect 240796 480 240824 3334
rect 242820 3330 242848 97135
rect 245568 78056 245620 78062
rect 245568 77998 245620 78004
rect 242900 76628 242952 76634
rect 242900 76570 242952 76576
rect 241980 3324 242032 3330
rect 241980 3266 242032 3272
rect 242808 3324 242860 3330
rect 242808 3266 242860 3272
rect 241992 480 242020 3266
rect 242912 626 242940 76570
rect 244372 9240 244424 9246
rect 244372 9182 244424 9188
rect 242912 598 243216 626
rect 243188 480 243216 598
rect 244384 480 244412 9182
rect 245580 480 245608 77998
rect 248248 33794 248276 102054
rect 249708 93560 249760 93566
rect 249708 93502 249760 93508
rect 248326 72448 248382 72457
rect 248326 72383 248382 72392
rect 248236 33788 248288 33794
rect 248236 33730 248288 33736
rect 246948 25696 247000 25702
rect 246948 25638 247000 25644
rect 246960 626 246988 25638
rect 246776 598 246988 626
rect 248340 610 248368 72383
rect 249720 3398 249748 93502
rect 251008 50386 251036 102054
rect 252572 102054 252954 102082
rect 251824 100088 251876 100094
rect 251824 100030 251876 100036
rect 251088 98864 251140 98870
rect 251088 98806 251140 98812
rect 250996 50380 251048 50386
rect 250996 50322 251048 50328
rect 251100 3398 251128 98806
rect 251836 25770 251864 100030
rect 252572 32570 252600 102054
rect 255332 100502 255360 102068
rect 256712 102054 257922 102082
rect 255320 100496 255372 100502
rect 255320 100438 255372 100444
rect 256608 100496 256660 100502
rect 256608 100438 256660 100444
rect 253848 86352 253900 86358
rect 253848 86294 253900 86300
rect 252560 32564 252612 32570
rect 252560 32506 252612 32512
rect 251824 25764 251876 25770
rect 251824 25706 251876 25712
rect 253754 9344 253810 9353
rect 253754 9279 253810 9288
rect 252652 3664 252704 3670
rect 252652 3606 252704 3612
rect 249156 3392 249208 3398
rect 249156 3334 249208 3340
rect 249708 3392 249760 3398
rect 249708 3334 249760 3340
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 251456 3392 251508 3398
rect 251456 3334 251508 3340
rect 247960 604 248012 610
rect 246776 480 246804 598
rect 247960 546 248012 552
rect 248328 604 248380 610
rect 248328 546 248380 552
rect 247972 480 248000 546
rect 249168 480 249196 3334
rect 250364 480 250392 3334
rect 251468 480 251496 3334
rect 252664 480 252692 3606
rect 253768 3482 253796 9279
rect 253860 3670 253888 86294
rect 256516 66972 256568 66978
rect 256516 66914 256568 66920
rect 253940 10464 253992 10470
rect 253940 10406 253992 10412
rect 253848 3664 253900 3670
rect 253848 3606 253900 3612
rect 253952 3482 253980 10406
rect 256528 3482 256556 66914
rect 256620 32434 256648 100438
rect 256608 32428 256660 32434
rect 256608 32370 256660 32376
rect 256712 6662 256740 102054
rect 260300 100026 260328 102068
rect 262890 102054 263548 102082
rect 261484 100156 261536 100162
rect 261484 100098 261536 100104
rect 260288 100020 260340 100026
rect 260288 99962 260340 99968
rect 261496 84862 261524 100098
rect 263414 86320 263470 86329
rect 263414 86255 263470 86264
rect 261484 84856 261536 84862
rect 261484 84798 261536 84804
rect 260748 61464 260800 61470
rect 260748 61406 260800 61412
rect 256700 6656 256752 6662
rect 256700 6598 256752 6604
rect 258632 6520 258684 6526
rect 258632 6462 258684 6468
rect 257436 3868 257488 3874
rect 257436 3810 257488 3816
rect 253768 3454 253888 3482
rect 253952 3454 255084 3482
rect 253860 480 253888 3454
rect 255056 480 255084 3454
rect 256252 3454 256556 3482
rect 256252 480 256280 3454
rect 257448 480 257476 3810
rect 258644 480 258672 6462
rect 259366 6080 259422 6089
rect 259366 6015 259422 6024
rect 259380 5681 259408 6015
rect 260760 5914 260788 61406
rect 260840 12300 260892 12306
rect 260840 12242 260892 12248
rect 259828 5908 259880 5914
rect 259828 5850 259880 5856
rect 260748 5908 260800 5914
rect 260748 5850 260800 5856
rect 259366 5672 259422 5681
rect 259366 5607 259422 5616
rect 259840 480 259868 5850
rect 260852 3482 260880 12242
rect 263322 3632 263378 3641
rect 263322 3567 263378 3576
rect 260852 3454 261064 3482
rect 261036 480 261064 3454
rect 262220 3392 262272 3398
rect 262220 3334 262272 3340
rect 262232 480 262260 3334
rect 263336 3210 263364 3567
rect 263428 3398 263456 86255
rect 263520 6526 263548 102054
rect 265268 99686 265296 102068
rect 267844 100502 267872 102068
rect 269132 102054 270250 102082
rect 272642 102054 273208 102082
rect 267832 100496 267884 100502
rect 267832 100438 267884 100444
rect 269028 100496 269080 100502
rect 269028 100438 269080 100444
rect 265256 99680 265308 99686
rect 265256 99622 265308 99628
rect 266268 99680 266320 99686
rect 266268 99622 266320 99628
rect 263600 78124 263652 78130
rect 263600 78066 263652 78072
rect 263508 6520 263560 6526
rect 263508 6462 263560 6468
rect 263612 3482 263640 78066
rect 266174 71224 266230 71233
rect 266174 71159 266230 71168
rect 266188 3482 266216 71159
rect 266280 26994 266308 99622
rect 266358 71360 266414 71369
rect 266358 71295 266414 71304
rect 266268 26988 266320 26994
rect 266268 26930 266320 26936
rect 263612 3454 264652 3482
rect 263416 3392 263468 3398
rect 263416 3334 263468 3340
rect 263336 3182 263456 3210
rect 263428 480 263456 3182
rect 264624 480 264652 3454
rect 265820 3454 266216 3482
rect 266372 3482 266400 71295
rect 267740 61600 267792 61606
rect 267740 61542 267792 61548
rect 267752 3482 267780 61542
rect 269040 22846 269068 100438
rect 269132 61674 269160 102054
rect 271788 79416 271840 79422
rect 271788 79358 271840 79364
rect 269120 61668 269172 61674
rect 269120 61610 269172 61616
rect 269028 22840 269080 22846
rect 269028 22782 269080 22788
rect 269120 12232 269172 12238
rect 269120 12174 269172 12180
rect 269132 3482 269160 12174
rect 270500 3732 270552 3738
rect 270500 3674 270552 3680
rect 266372 3454 267044 3482
rect 267752 3454 268148 3482
rect 269132 3454 269344 3482
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 268120 480 268148 3454
rect 269316 480 269344 3454
rect 270512 480 270540 3674
rect 271800 3482 271828 79358
rect 273180 9246 273208 102054
rect 273168 9240 273220 9246
rect 273168 9182 273220 9188
rect 273902 5808 273958 5817
rect 273902 5743 273958 5752
rect 273916 5545 273944 5743
rect 273902 5536 273958 5545
rect 273902 5471 273958 5480
rect 272892 4820 272944 4826
rect 272892 4762 272944 4768
rect 271708 3454 271828 3482
rect 271708 480 271736 3454
rect 272904 480 272932 4762
rect 274560 4078 274588 102439
rect 274652 102054 275218 102082
rect 274652 86426 274680 102054
rect 277596 100298 277624 102068
rect 280172 100502 280200 102068
rect 282578 102054 282868 102082
rect 280160 100496 280212 100502
rect 280160 100438 280212 100444
rect 281448 100496 281500 100502
rect 281448 100438 281500 100444
rect 277584 100292 277636 100298
rect 277584 100234 277636 100240
rect 280528 99340 280580 99346
rect 280528 99282 280580 99288
rect 280540 96642 280568 99282
rect 280540 96614 280660 96642
rect 275928 96076 275980 96082
rect 275928 96018 275980 96024
rect 274640 86420 274692 86426
rect 274640 86362 274692 86368
rect 275940 4078 275968 96018
rect 278688 91860 278740 91866
rect 278688 91802 278740 91808
rect 276480 12164 276532 12170
rect 276480 12106 276532 12112
rect 274088 4072 274140 4078
rect 274088 4014 274140 4020
rect 274548 4072 274600 4078
rect 274548 4014 274600 4020
rect 275284 4072 275336 4078
rect 275284 4014 275336 4020
rect 275928 4072 275980 4078
rect 275928 4014 275980 4020
rect 274100 480 274128 4014
rect 275296 480 275324 4014
rect 276492 480 276520 12106
rect 278700 3262 278728 91802
rect 280632 89706 280660 96614
rect 280540 89678 280660 89706
rect 280068 89004 280120 89010
rect 280068 88946 280120 88952
rect 279976 9444 280028 9450
rect 279976 9386 280028 9392
rect 278872 4072 278924 4078
rect 278872 4014 278924 4020
rect 277676 3256 277728 3262
rect 277676 3198 277728 3204
rect 278688 3256 278740 3262
rect 278688 3198 278740 3204
rect 277688 480 277716 3198
rect 278884 480 278912 4014
rect 279988 3890 280016 9386
rect 280080 4078 280108 88946
rect 280540 86970 280568 89678
rect 280528 86964 280580 86970
rect 280528 86906 280580 86912
rect 280436 77308 280488 77314
rect 280436 77250 280488 77256
rect 280448 77217 280476 77250
rect 280250 77208 280306 77217
rect 280250 77143 280306 77152
rect 280434 77208 280490 77217
rect 280434 77143 280490 77152
rect 280264 70446 280292 77143
rect 280252 70440 280304 70446
rect 280252 70382 280304 70388
rect 280344 70372 280396 70378
rect 280344 70314 280396 70320
rect 280356 60738 280384 70314
rect 280356 60710 280476 60738
rect 280448 57934 280476 60710
rect 280436 57928 280488 57934
rect 280436 57870 280488 57876
rect 280344 48340 280396 48346
rect 280344 48282 280396 48288
rect 280356 41426 280384 48282
rect 281460 46306 281488 100438
rect 281448 46300 281500 46306
rect 281448 46242 281500 46248
rect 280356 41398 280476 41426
rect 280448 38622 280476 41398
rect 280436 38616 280488 38622
rect 280436 38558 280488 38564
rect 280344 31748 280396 31754
rect 280344 31690 280396 31696
rect 280356 22114 280384 31690
rect 281540 24132 281592 24138
rect 281540 24074 281592 24080
rect 280356 22086 280476 22114
rect 280448 12458 280476 22086
rect 280264 12442 280476 12458
rect 281552 12442 281580 24074
rect 282840 20126 282868 102054
rect 285140 100706 285168 102068
rect 285128 100700 285180 100706
rect 285128 100642 285180 100648
rect 286324 100292 286376 100298
rect 286324 100234 286376 100240
rect 284208 98932 284260 98938
rect 284208 98874 284260 98880
rect 282828 20120 282880 20126
rect 282828 20062 282880 20068
rect 280252 12436 280476 12442
rect 280304 12430 280476 12436
rect 281172 12436 281224 12442
rect 280252 12378 280304 12384
rect 281172 12378 281224 12384
rect 281540 12436 281592 12442
rect 281540 12378 281592 12384
rect 282460 12436 282512 12442
rect 282460 12378 282512 12384
rect 280264 12347 280292 12378
rect 281184 12322 281212 12378
rect 281184 12294 281304 12322
rect 280068 4072 280120 4078
rect 280068 4014 280120 4020
rect 279988 3862 280108 3890
rect 280080 480 280108 3862
rect 281276 480 281304 12294
rect 282472 480 282500 12378
rect 282826 5808 282882 5817
rect 283010 5808 283066 5817
rect 282882 5766 283010 5794
rect 282826 5743 282882 5752
rect 283010 5743 283066 5752
rect 284220 3398 284248 98874
rect 284300 71120 284352 71126
rect 284300 71062 284352 71068
rect 284312 3482 284340 71062
rect 286336 9110 286364 100234
rect 287532 99414 287560 102068
rect 289832 102054 289938 102082
rect 287520 99408 287572 99414
rect 287520 99350 287572 99356
rect 288348 99408 288400 99414
rect 288348 99350 288400 99356
rect 287060 83632 287112 83638
rect 287060 83574 287112 83580
rect 286968 15972 287020 15978
rect 286968 15914 287020 15920
rect 286324 9104 286376 9110
rect 286324 9046 286376 9052
rect 284312 3454 284800 3482
rect 283656 3392 283708 3398
rect 283656 3334 283708 3340
rect 284208 3392 284260 3398
rect 284208 3334 284260 3340
rect 283668 480 283696 3334
rect 284772 480 284800 3454
rect 286980 3398 287008 15914
rect 287072 3398 287100 83574
rect 288360 15026 288388 99350
rect 289726 98968 289782 98977
rect 289726 98903 289782 98912
rect 288348 15020 288400 15026
rect 288348 14962 288400 14968
rect 287152 4888 287204 4894
rect 287152 4830 287204 4836
rect 285956 3392 286008 3398
rect 285956 3334 286008 3340
rect 286968 3392 287020 3398
rect 286968 3334 287020 3340
rect 287060 3392 287112 3398
rect 287060 3334 287112 3340
rect 285968 480 285996 3334
rect 287164 480 287192 4830
rect 289740 3482 289768 98903
rect 289832 68474 289860 102054
rect 292500 100706 292528 102068
rect 293972 102054 294906 102082
rect 297482 102054 297956 102082
rect 292488 100700 292540 100706
rect 292488 100642 292540 100648
rect 293868 87644 293920 87650
rect 293868 87586 293920 87592
rect 289820 68468 289872 68474
rect 289820 68410 289872 68416
rect 290740 9308 290792 9314
rect 290740 9250 290792 9256
rect 289556 3454 289768 3482
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 288360 480 288388 3334
rect 289556 480 289584 3454
rect 290752 480 290780 9250
rect 291936 4956 291988 4962
rect 291936 4898 291988 4904
rect 291948 480 291976 4898
rect 293880 3398 293908 87586
rect 293972 13122 294000 102054
rect 294052 32496 294104 32502
rect 294052 32438 294104 32444
rect 293960 13116 294012 13122
rect 293960 13058 294012 13064
rect 294064 3482 294092 32438
rect 297824 29776 297876 29782
rect 297824 29718 297876 29724
rect 295522 7576 295578 7585
rect 295522 7511 295578 7520
rect 294064 3454 294368 3482
rect 293132 3392 293184 3398
rect 293132 3334 293184 3340
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 293144 480 293172 3334
rect 294340 480 294368 3454
rect 295536 480 295564 7511
rect 297836 3482 297864 29718
rect 297928 21486 297956 102054
rect 299492 102054 299874 102082
rect 302252 102054 302450 102082
rect 303632 102054 304842 102082
rect 307234 102054 307616 102082
rect 298008 90432 298060 90438
rect 298008 90374 298060 90380
rect 297916 21480 297968 21486
rect 297916 21422 297968 21428
rect 297836 3454 297956 3482
rect 296720 3392 296772 3398
rect 296720 3334 296772 3340
rect 296732 480 296760 3334
rect 297928 480 297956 3454
rect 298020 3398 298048 90374
rect 299492 7682 299520 102054
rect 302148 100020 302200 100026
rect 302148 99962 302200 99968
rect 299480 7676 299532 7682
rect 299480 7618 299532 7624
rect 300308 3800 300360 3806
rect 300308 3742 300360 3748
rect 299110 3496 299166 3505
rect 299110 3431 299166 3440
rect 298008 3392 298060 3398
rect 298008 3334 298060 3340
rect 299124 480 299152 3431
rect 300320 480 300348 3742
rect 302160 3398 302188 99962
rect 302252 3482 302280 102054
rect 303632 66978 303660 102054
rect 306288 99000 306340 99006
rect 306288 98942 306340 98948
rect 304906 97336 304962 97345
rect 304906 97271 304962 97280
rect 303620 66972 303672 66978
rect 303620 66914 303672 66920
rect 302252 3454 302648 3482
rect 301412 3392 301464 3398
rect 301412 3334 301464 3340
rect 302148 3392 302200 3398
rect 302148 3334 302200 3340
rect 301424 480 301452 3334
rect 302620 480 302648 3454
rect 304920 3398 304948 97271
rect 305000 89072 305052 89078
rect 305000 89014 305052 89020
rect 305012 3398 305040 89014
rect 303804 3392 303856 3398
rect 303804 3334 303856 3340
rect 304908 3392 304960 3398
rect 304908 3334 304960 3340
rect 305000 3392 305052 3398
rect 305000 3334 305052 3340
rect 306196 3392 306248 3398
rect 306196 3334 306248 3340
rect 303816 480 303844 3334
rect 305000 3256 305052 3262
rect 305000 3198 305052 3204
rect 305012 480 305040 3198
rect 306208 480 306236 3334
rect 306300 3262 306328 98942
rect 307588 39370 307616 102054
rect 307576 39364 307628 39370
rect 307576 39306 307628 39312
rect 307680 3482 307708 102575
rect 309244 102054 309810 102082
rect 311912 102054 312202 102082
rect 309138 94480 309194 94489
rect 309138 94415 309194 94424
rect 308588 9172 308640 9178
rect 308588 9114 308640 9120
rect 307404 3454 307708 3482
rect 306288 3256 306340 3262
rect 306288 3198 306340 3204
rect 307404 480 307432 3454
rect 308600 480 308628 9114
rect 309152 3482 309180 94415
rect 309244 75206 309272 102054
rect 309232 75200 309284 75206
rect 309232 75142 309284 75148
rect 311912 31074 311940 102054
rect 314764 100298 314792 102068
rect 314752 100292 314804 100298
rect 314752 100234 314804 100240
rect 317156 99414 317184 102068
rect 319746 102054 320128 102082
rect 315304 99408 315356 99414
rect 315304 99350 315356 99356
rect 317144 99408 317196 99414
rect 317144 99350 317196 99356
rect 314568 84856 314620 84862
rect 314568 84798 314620 84804
rect 311992 61532 312044 61538
rect 311992 61474 312044 61480
rect 311900 31068 311952 31074
rect 311900 31010 311952 31016
rect 310520 15020 310572 15026
rect 310520 14962 310572 14968
rect 310532 3482 310560 14962
rect 312004 3482 312032 61474
rect 313372 6520 313424 6526
rect 313372 6462 313424 6468
rect 309152 3454 309824 3482
rect 310532 3454 311020 3482
rect 312004 3454 312216 3482
rect 309796 480 309824 3454
rect 310992 480 311020 3454
rect 312188 480 312216 3454
rect 313384 480 313412 6462
rect 314580 480 314608 84798
rect 315316 3602 315344 99350
rect 319994 95976 320050 95985
rect 319994 95911 320050 95920
rect 315948 65612 316000 65618
rect 315948 65554 316000 65560
rect 315304 3596 315356 3602
rect 315304 3538 315356 3544
rect 315960 3482 315988 65554
rect 317326 51776 317382 51785
rect 317326 51711 317382 51720
rect 317340 3482 317368 51711
rect 318064 6452 318116 6458
rect 318064 6394 318116 6400
rect 315776 3454 315988 3482
rect 316972 3454 317368 3482
rect 315776 480 315804 3454
rect 316972 480 317000 3454
rect 318076 480 318104 6394
rect 320008 3058 320036 95911
rect 320100 5166 320128 102054
rect 322124 100638 322152 102068
rect 324226 101824 324282 101833
rect 324226 101759 324282 101768
rect 322846 101688 322902 101697
rect 322846 101623 322902 101632
rect 322112 100632 322164 100638
rect 322112 100574 322164 100580
rect 320180 68400 320232 68406
rect 320180 68342 320232 68348
rect 320088 5160 320140 5166
rect 320088 5102 320140 5108
rect 320192 3482 320220 68342
rect 322860 3602 322888 101623
rect 323584 99408 323636 99414
rect 323584 99350 323636 99356
rect 323596 58750 323624 99350
rect 323584 58744 323636 58750
rect 323584 58686 323636 58692
rect 321652 3596 321704 3602
rect 321652 3538 321704 3544
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 322940 3596 322992 3602
rect 322940 3538 322992 3544
rect 320192 3454 320496 3482
rect 319260 3052 319312 3058
rect 319260 2994 319312 3000
rect 319996 3052 320048 3058
rect 319996 2994 320048 3000
rect 319272 480 319300 2994
rect 320468 480 320496 3454
rect 321664 480 321692 3538
rect 322952 3482 322980 3538
rect 324240 3482 324268 101759
rect 324516 99414 324544 102068
rect 327092 100638 327120 102068
rect 327080 100632 327132 100638
rect 327080 100574 327132 100580
rect 329484 100570 329512 102068
rect 329472 100564 329524 100570
rect 329472 100506 329524 100512
rect 327724 100292 327776 100298
rect 327724 100234 327776 100240
rect 324504 99408 324556 99414
rect 324504 99350 324556 99356
rect 326988 96144 327040 96150
rect 326988 96086 327040 96092
rect 325238 6352 325294 6361
rect 325238 6287 325294 6296
rect 322860 3454 322980 3482
rect 324056 3454 324268 3482
rect 322860 480 322888 3454
rect 324056 480 324084 3454
rect 325252 480 325280 6287
rect 327000 3398 327028 96086
rect 327736 15910 327764 100234
rect 334452 99414 334480 102068
rect 336752 102054 337042 102082
rect 338132 102054 339434 102082
rect 334440 99408 334492 99414
rect 334440 99350 334492 99356
rect 335268 99408 335320 99414
rect 335268 99350 335320 99356
rect 331128 99068 331180 99074
rect 331128 99010 331180 99016
rect 329748 97300 329800 97306
rect 329748 97242 329800 97248
rect 327724 15904 327776 15910
rect 327724 15846 327776 15852
rect 327632 5024 327684 5030
rect 327632 4966 327684 4972
rect 326436 3392 326488 3398
rect 326436 3334 326488 3340
rect 326988 3392 327040 3398
rect 326988 3334 327040 3340
rect 326448 480 326476 3334
rect 327644 480 327672 4966
rect 329760 3194 329788 97242
rect 330850 5808 330906 5817
rect 330906 5766 330984 5794
rect 330850 5743 330906 5752
rect 330956 5681 330984 5766
rect 330942 5672 330998 5681
rect 330942 5607 330998 5616
rect 331140 3398 331168 99010
rect 331218 98832 331274 98841
rect 331218 98767 331274 98776
rect 331232 7682 331260 98767
rect 332508 73908 332560 73914
rect 332508 73850 332560 73856
rect 331220 7676 331272 7682
rect 331220 7618 331272 7624
rect 332416 7676 332468 7682
rect 332416 7618 332468 7624
rect 331220 4072 331272 4078
rect 331220 4014 331272 4020
rect 330024 3392 330076 3398
rect 330024 3334 330076 3340
rect 331128 3392 331180 3398
rect 331128 3334 331180 3340
rect 328828 3188 328880 3194
rect 328828 3130 328880 3136
rect 329748 3188 329800 3194
rect 329748 3130 329800 3136
rect 328840 480 328868 3130
rect 330036 480 330064 3334
rect 331232 480 331260 4014
rect 332428 480 332456 7618
rect 332520 4078 332548 73850
rect 333888 60172 333940 60178
rect 333888 60114 333940 60120
rect 333900 57934 333928 60114
rect 333888 57928 333940 57934
rect 333888 57870 333940 57876
rect 333888 48340 333940 48346
rect 333888 48282 333940 48288
rect 333900 19310 333928 48282
rect 335280 46306 335308 99350
rect 335360 90364 335412 90370
rect 335360 90306 335412 90312
rect 333980 46300 334032 46306
rect 333980 46242 334032 46248
rect 335268 46300 335320 46306
rect 335268 46242 335320 46248
rect 333992 19310 334020 46242
rect 333888 19304 333940 19310
rect 333888 19246 333940 19252
rect 333980 19304 334032 19310
rect 333980 19246 334032 19252
rect 334808 19304 334860 19310
rect 334808 19246 334860 19252
rect 333888 9716 333940 9722
rect 333888 9658 333940 9664
rect 332508 4072 332560 4078
rect 332508 4014 332560 4020
rect 333900 2854 333928 9658
rect 334820 3176 334848 19246
rect 335372 12442 335400 90306
rect 335360 12436 335412 12442
rect 335360 12378 335412 12384
rect 335912 12436 335964 12442
rect 335912 12378 335964 12384
rect 334728 3148 334848 3176
rect 333888 2848 333940 2854
rect 333888 2790 333940 2796
rect 333612 2780 333664 2786
rect 333612 2722 333664 2728
rect 333624 480 333652 2722
rect 334728 480 334756 3148
rect 335924 480 335952 12378
rect 336752 9382 336780 102054
rect 338132 73846 338160 102054
rect 341812 100298 341840 102068
rect 344402 102054 344876 102082
rect 341800 100292 341852 100298
rect 341800 100234 341852 100240
rect 342260 86284 342312 86290
rect 342260 86226 342312 86232
rect 338120 73840 338172 73846
rect 338120 73782 338172 73788
rect 342168 72548 342220 72554
rect 342168 72490 342220 72496
rect 338028 69760 338080 69766
rect 338028 69702 338080 69708
rect 336740 9376 336792 9382
rect 336740 9318 336792 9324
rect 338040 4078 338068 69702
rect 340786 57216 340842 57225
rect 340786 57151 340842 57160
rect 338212 20052 338264 20058
rect 338212 19994 338264 20000
rect 338224 19394 338252 19994
rect 338132 19366 338252 19394
rect 338132 19310 338160 19366
rect 338120 19304 338172 19310
rect 338120 19246 338172 19252
rect 338304 9716 338356 9722
rect 338304 9658 338356 9664
rect 337108 4072 337160 4078
rect 337108 4014 337160 4020
rect 338028 4072 338080 4078
rect 338028 4014 338080 4020
rect 337120 480 337148 4014
rect 338316 480 338344 9658
rect 340696 9036 340748 9042
rect 340696 8978 340748 8984
rect 339500 3324 339552 3330
rect 339500 3266 339552 3272
rect 339512 480 339540 3266
rect 340708 480 340736 8978
rect 340800 3330 340828 57151
rect 342180 3482 342208 72490
rect 341904 3454 342208 3482
rect 342272 3482 342300 86226
rect 344848 57322 344876 102054
rect 344926 98832 344982 98841
rect 344926 98767 344982 98776
rect 344836 57316 344888 57322
rect 344836 57258 344888 57264
rect 342272 3454 343128 3482
rect 340788 3324 340840 3330
rect 340788 3266 340840 3272
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344940 3398 344968 98767
rect 346780 97918 346808 102068
rect 350552 102054 351762 102082
rect 354338 102054 354536 102082
rect 346768 97912 346820 97918
rect 346768 97854 346820 97860
rect 349068 96212 349120 96218
rect 349068 96154 349120 96160
rect 348976 68400 349028 68406
rect 348976 68342 349028 68348
rect 345020 13864 345072 13870
rect 345020 13806 345072 13812
rect 345032 3482 345060 13806
rect 346674 9344 346730 9353
rect 346674 9279 346730 9288
rect 345032 3454 345520 3482
rect 344284 3392 344336 3398
rect 344284 3334 344336 3340
rect 344928 3392 344980 3398
rect 344928 3334 344980 3340
rect 344296 480 344324 3334
rect 345492 480 345520 3454
rect 346688 480 346716 9279
rect 347872 3052 347924 3058
rect 347872 2994 347924 3000
rect 347884 480 347912 2994
rect 348988 1578 349016 68342
rect 349080 3058 349108 96154
rect 350552 10402 350580 102054
rect 354508 56030 354536 102054
rect 356716 100230 356744 102068
rect 359108 100570 359136 102068
rect 361592 102054 361698 102082
rect 364090 102054 364288 102082
rect 359096 100564 359148 100570
rect 359096 100506 359148 100512
rect 360108 100564 360160 100570
rect 360108 100506 360160 100512
rect 356704 100224 356756 100230
rect 356704 100166 356756 100172
rect 354588 99136 354640 99142
rect 354588 99078 354640 99084
rect 350632 56024 350684 56030
rect 350632 55966 350684 55972
rect 354496 56024 354548 56030
rect 354496 55966 354548 55972
rect 350644 12442 350672 55966
rect 353300 32496 353352 32502
rect 353300 32438 353352 32444
rect 353312 27266 353340 32438
rect 351184 27260 351236 27266
rect 351184 27202 351236 27208
rect 353300 27260 353352 27266
rect 353300 27202 353352 27208
rect 351196 13870 351224 27202
rect 351920 14952 351972 14958
rect 351920 14894 351972 14900
rect 351184 13864 351236 13870
rect 351184 13806 351236 13812
rect 351932 12442 351960 14894
rect 350632 12436 350684 12442
rect 350632 12378 350684 12384
rect 351368 12436 351420 12442
rect 351368 12378 351420 12384
rect 351920 12436 351972 12442
rect 351920 12378 351972 12384
rect 352564 12436 352616 12442
rect 352564 12378 352616 12384
rect 350540 10396 350592 10402
rect 350540 10338 350592 10344
rect 350446 5672 350502 5681
rect 350630 5672 350686 5681
rect 350502 5630 350630 5658
rect 350446 5607 350502 5616
rect 350630 5607 350686 5616
rect 350264 5092 350316 5098
rect 350264 5034 350316 5040
rect 349068 3052 349120 3058
rect 349068 2994 349120 3000
rect 348988 1550 349108 1578
rect 349080 480 349108 1550
rect 350276 480 350304 5034
rect 351380 480 351408 12378
rect 352576 480 352604 12378
rect 354600 3194 354628 99078
rect 355968 97368 356020 97374
rect 355968 97310 356020 97316
rect 355980 3194 356008 97310
rect 356520 96688 356572 96694
rect 356520 96630 356572 96636
rect 356532 89758 356560 96630
rect 357346 96112 357402 96121
rect 357346 96047 357402 96056
rect 356520 89752 356572 89758
rect 356520 89694 356572 89700
rect 356612 89616 356664 89622
rect 356612 89558 356664 89564
rect 356624 80102 356652 89558
rect 356612 80096 356664 80102
rect 356612 80038 356664 80044
rect 356704 79960 356756 79966
rect 356704 79902 356756 79908
rect 356716 77178 356744 79902
rect 356704 77172 356756 77178
rect 356704 77114 356756 77120
rect 356796 70304 356848 70310
rect 356796 70246 356848 70252
rect 356808 60738 356836 70246
rect 356624 60710 356836 60738
rect 356624 57934 356652 60710
rect 356612 57928 356664 57934
rect 356612 57870 356664 57876
rect 357256 50448 357308 50454
rect 357256 50390 357308 50396
rect 356704 48340 356756 48346
rect 356704 48282 356756 48288
rect 356716 41426 356744 48282
rect 356716 41398 356928 41426
rect 356900 38078 356928 41398
rect 356888 38072 356940 38078
rect 356888 38014 356940 38020
rect 356152 4072 356204 4078
rect 356152 4014 356204 4020
rect 353760 3188 353812 3194
rect 353760 3130 353812 3136
rect 354588 3188 354640 3194
rect 354588 3130 354640 3136
rect 354956 3188 355008 3194
rect 354956 3130 355008 3136
rect 355968 3188 356020 3194
rect 355968 3130 356020 3136
rect 353772 480 353800 3130
rect 354968 480 354996 3130
rect 356164 480 356192 4014
rect 357268 1578 357296 50390
rect 357360 4078 357388 96047
rect 360120 65686 360148 100506
rect 360200 76560 360252 76566
rect 360200 76502 360252 76508
rect 360108 65680 360160 65686
rect 360108 65622 360160 65628
rect 358820 42084 358872 42090
rect 358820 42026 358872 42032
rect 358544 8968 358596 8974
rect 358544 8910 358596 8916
rect 357348 4072 357400 4078
rect 357348 4014 357400 4020
rect 357268 1550 357388 1578
rect 357360 480 357388 1550
rect 358556 480 358584 8910
rect 358832 610 358860 42026
rect 360212 3482 360240 76502
rect 360844 39432 360896 39438
rect 360844 39374 360896 39380
rect 360856 32502 360884 39374
rect 360844 32496 360896 32502
rect 360844 32438 360896 32444
rect 360212 3454 360976 3482
rect 358820 604 358872 610
rect 358820 546 358872 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 359752 480 359780 546
rect 360948 480 360976 3454
rect 361592 3398 361620 102054
rect 364156 71120 364208 71126
rect 364156 71062 364208 71068
rect 364168 3398 364196 71062
rect 364260 18766 364288 102054
rect 365732 102054 366666 102082
rect 368492 102054 369058 102082
rect 365628 97436 365680 97442
rect 365628 97378 365680 97384
rect 364248 18760 364300 18766
rect 364248 18702 364300 18708
rect 365640 3398 365668 97378
rect 365732 71058 365760 102054
rect 367008 94580 367060 94586
rect 367008 94522 367060 94528
rect 365720 71052 365772 71058
rect 365720 70994 365772 71000
rect 365720 17400 365772 17406
rect 365720 17342 365772 17348
rect 365732 3398 365760 17342
rect 361580 3392 361632 3398
rect 361580 3334 361632 3340
rect 362132 3392 362184 3398
rect 362132 3334 362184 3340
rect 363328 3392 363380 3398
rect 363328 3334 363380 3340
rect 364156 3392 364208 3398
rect 364156 3334 364208 3340
rect 364524 3392 364576 3398
rect 364524 3334 364576 3340
rect 365628 3392 365680 3398
rect 365628 3334 365680 3340
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 366916 3392 366968 3398
rect 366916 3334 366968 3340
rect 362144 480 362172 3334
rect 363340 480 363368 3334
rect 364536 480 364564 3334
rect 365720 3256 365772 3262
rect 365720 3198 365772 3204
rect 365732 480 365760 3198
rect 366928 480 366956 3334
rect 367020 3262 367048 94522
rect 367100 40792 367152 40798
rect 367100 40734 367152 40740
rect 367112 3482 367140 40734
rect 368492 16114 368520 102054
rect 370516 39438 370544 102614
rect 371252 102054 371634 102082
rect 370596 100224 370648 100230
rect 370596 100166 370648 100172
rect 370608 60110 370636 100166
rect 371252 71126 371280 102054
rect 374012 99414 374040 102068
rect 376404 100298 376432 102068
rect 378244 102054 378994 102082
rect 376392 100292 376444 100298
rect 376392 100234 376444 100240
rect 374000 99408 374052 99414
rect 374000 99350 374052 99356
rect 375288 99408 375340 99414
rect 375288 99350 375340 99356
rect 371240 71120 371292 71126
rect 371240 71062 371292 71068
rect 375196 71052 375248 71058
rect 375196 70994 375248 71000
rect 371148 66972 371200 66978
rect 371148 66914 371200 66920
rect 370596 60104 370648 60110
rect 370596 60046 370648 60052
rect 370504 39432 370556 39438
rect 370504 39374 370556 39380
rect 368480 16108 368532 16114
rect 368480 16050 368532 16056
rect 369214 9072 369270 9081
rect 369214 9007 369270 9016
rect 367112 3454 368060 3482
rect 367008 3256 367060 3262
rect 367008 3198 367060 3204
rect 368032 480 368060 3454
rect 369228 480 369256 9007
rect 371160 3398 371188 66914
rect 371240 14884 371292 14890
rect 371240 14826 371292 14832
rect 371252 3482 371280 14826
rect 372620 12096 372672 12102
rect 372620 12038 372672 12044
rect 372632 3482 372660 12038
rect 371252 3454 371648 3482
rect 372632 3454 372844 3482
rect 370412 3392 370464 3398
rect 370412 3334 370464 3340
rect 371148 3392 371200 3398
rect 371148 3334 371200 3340
rect 370424 480 370452 3334
rect 371620 480 371648 3454
rect 372816 480 372844 3454
rect 375208 3398 375236 70994
rect 375300 14890 375328 99350
rect 378140 79348 378192 79354
rect 378140 79290 378192 79296
rect 376760 57248 376812 57254
rect 376760 57190 376812 57196
rect 375288 14884 375340 14890
rect 375288 14826 375340 14832
rect 376392 9036 376444 9042
rect 376392 8978 376444 8984
rect 375286 5808 375342 5817
rect 375286 5743 375342 5752
rect 375300 5545 375328 5743
rect 375286 5536 375342 5545
rect 375286 5471 375342 5480
rect 375288 3868 375340 3874
rect 375288 3810 375340 3816
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 374012 480 374040 3334
rect 375300 1986 375328 3810
rect 375208 1958 375328 1986
rect 375208 480 375236 1958
rect 376404 480 376432 8978
rect 376772 610 376800 57190
rect 378152 3482 378180 79290
rect 378244 66978 378272 102054
rect 381372 99414 381400 102068
rect 383948 99414 383976 102068
rect 385052 102054 386354 102082
rect 381360 99408 381412 99414
rect 381360 99350 381412 99356
rect 382188 99408 382240 99414
rect 382188 99350 382240 99356
rect 383936 99408 383988 99414
rect 383936 99350 383988 99356
rect 384948 99408 385000 99414
rect 384948 99350 385000 99356
rect 378232 66972 378284 66978
rect 378232 66914 378284 66920
rect 380808 57248 380860 57254
rect 380808 57190 380860 57196
rect 378692 5092 378744 5098
rect 378692 5034 378744 5040
rect 378704 3806 378732 5034
rect 378692 3800 378744 3806
rect 378692 3742 378744 3748
rect 378152 3454 378824 3482
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 377600 480 377628 546
rect 378796 480 378824 3454
rect 380820 3398 380848 57190
rect 382200 49162 382228 99350
rect 384960 51746 384988 99350
rect 385052 73982 385080 102054
rect 388916 100502 388944 102068
rect 391322 102054 391888 102082
rect 388904 100496 388956 100502
rect 388904 100438 388956 100444
rect 389088 96280 389140 96286
rect 389088 96222 389140 96228
rect 386328 93628 386380 93634
rect 386328 93570 386380 93576
rect 385040 73976 385092 73982
rect 385040 73918 385092 73924
rect 382280 51740 382332 51746
rect 382280 51682 382332 51688
rect 384948 51740 385000 51746
rect 384948 51682 385000 51688
rect 382188 49156 382240 49162
rect 382188 49098 382240 49104
rect 381174 3496 381230 3505
rect 381174 3431 381230 3440
rect 379980 3392 380032 3398
rect 379980 3334 380032 3340
rect 380808 3392 380860 3398
rect 380808 3334 380860 3340
rect 379992 480 380020 3334
rect 381188 480 381216 3431
rect 382292 3398 382320 51682
rect 384948 16108 385000 16114
rect 384948 16050 385000 16056
rect 382372 8968 382424 8974
rect 382372 8910 382424 8916
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 8910
rect 384960 3482 384988 16050
rect 384684 3454 384988 3482
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 384684 480 384712 3454
rect 386340 3398 386368 93570
rect 386418 11792 386474 11801
rect 386418 11727 386474 11736
rect 386432 3482 386460 11727
rect 386432 3454 387104 3482
rect 385868 3392 385920 3398
rect 385868 3334 385920 3340
rect 386328 3392 386380 3398
rect 386328 3334 386380 3340
rect 385880 480 385908 3334
rect 387076 480 387104 3454
rect 389100 3398 389128 96222
rect 389178 53136 389234 53145
rect 389178 53071 389234 53080
rect 391756 53100 391808 53106
rect 389192 19310 389220 53071
rect 391756 53042 391808 53048
rect 391768 19310 391796 53042
rect 391860 40798 391888 102054
rect 393700 100162 393728 102068
rect 396184 102054 396290 102082
rect 397472 102054 398682 102082
rect 393688 100156 393740 100162
rect 393688 100098 393740 100104
rect 393228 94648 393280 94654
rect 393228 94590 393280 94596
rect 391848 40792 391900 40798
rect 391848 40734 391900 40740
rect 389180 19304 389232 19310
rect 389180 19246 389232 19252
rect 391756 19304 391808 19310
rect 391756 19246 391808 19252
rect 389456 9716 389508 9722
rect 389456 9658 389508 9664
rect 391848 9716 391900 9722
rect 391848 9658 391900 9664
rect 388260 3392 388312 3398
rect 388260 3334 388312 3340
rect 389088 3392 389140 3398
rect 389088 3334 389140 3340
rect 388272 480 388300 3334
rect 389468 480 389496 9658
rect 390650 9208 390706 9217
rect 390650 9143 390706 9152
rect 390664 480 390692 9143
rect 391860 480 391888 9658
rect 393240 2854 393268 94590
rect 396080 82136 396132 82142
rect 396080 82078 396132 82084
rect 393320 50380 393372 50386
rect 393320 50322 393372 50328
rect 393228 2848 393280 2854
rect 393228 2790 393280 2796
rect 393332 610 393360 50322
rect 395434 9072 395490 9081
rect 395434 9007 395490 9016
rect 394606 6080 394662 6089
rect 394606 6015 394662 6024
rect 394620 5681 394648 6015
rect 394606 5672 394662 5681
rect 394606 5607 394662 5616
rect 393044 604 393096 610
rect 393044 546 393096 552
rect 393320 604 393372 610
rect 393320 546 393372 552
rect 394240 604 394292 610
rect 394240 546 394292 552
rect 393056 480 393084 546
rect 394252 480 394280 546
rect 395448 480 395476 9007
rect 396092 610 396120 82078
rect 396184 58818 396212 102054
rect 396172 58812 396224 58818
rect 396172 58754 396224 58760
rect 397472 16046 397500 102054
rect 401244 100434 401272 102068
rect 401232 100428 401284 100434
rect 401232 100370 401284 100376
rect 403636 100366 403664 102068
rect 403624 100360 403676 100366
rect 403624 100302 403676 100308
rect 406212 100094 406240 102068
rect 408604 100230 408632 102068
rect 410996 100570 411024 102068
rect 410984 100564 411036 100570
rect 410984 100506 411036 100512
rect 408592 100224 408644 100230
rect 408592 100166 408644 100172
rect 406200 100088 406252 100094
rect 406200 100030 406252 100036
rect 406382 99104 406438 99113
rect 406382 99039 406438 99048
rect 398748 96348 398800 96354
rect 398748 96290 398800 96296
rect 397460 16040 397512 16046
rect 397460 15982 397512 15988
rect 398760 4078 398788 96290
rect 400126 50416 400182 50425
rect 400126 50351 400182 50360
rect 400140 4078 400168 50351
rect 404360 49088 404412 49094
rect 404360 49030 404412 49036
rect 401600 26988 401652 26994
rect 401600 26930 401652 26936
rect 400220 22840 400272 22846
rect 400220 22782 400272 22788
rect 397828 4072 397880 4078
rect 397828 4014 397880 4020
rect 398748 4072 398800 4078
rect 398748 4014 398800 4020
rect 399024 4072 399076 4078
rect 399024 4014 399076 4020
rect 400128 4072 400180 4078
rect 400128 4014 400180 4020
rect 396080 604 396132 610
rect 396080 546 396132 552
rect 396632 604 396684 610
rect 396632 546 396684 552
rect 396644 480 396672 546
rect 397840 480 397868 4014
rect 399036 480 399064 4014
rect 400232 480 400260 22782
rect 401324 3800 401376 3806
rect 401324 3742 401376 3748
rect 401336 480 401364 3742
rect 401612 610 401640 26930
rect 404372 12442 404400 49030
rect 404360 12436 404412 12442
rect 404360 12378 404412 12384
rect 404912 12436 404964 12442
rect 404912 12378 404964 12384
rect 403714 6488 403770 6497
rect 403714 6423 403770 6432
rect 401600 604 401652 610
rect 401600 546 401652 552
rect 402520 604 402572 610
rect 402520 546 402572 552
rect 402532 480 402560 546
rect 403728 480 403756 6423
rect 404924 480 404952 12378
rect 406108 6656 406160 6662
rect 406108 6598 406160 6604
rect 406120 480 406148 6598
rect 406396 3874 406424 99039
rect 413572 96558 413600 102068
rect 415412 102054 415978 102082
rect 413560 96552 413612 96558
rect 413560 96494 413612 96500
rect 411168 87032 411220 87038
rect 411168 86974 411220 86980
rect 411180 77178 411208 86974
rect 411168 77172 411220 77178
rect 411168 77114 411220 77120
rect 411168 67652 411220 67658
rect 411168 67594 411220 67600
rect 411180 57934 411208 67594
rect 411168 57928 411220 57934
rect 411168 57870 411220 57876
rect 415412 50454 415440 102054
rect 415400 50448 415452 50454
rect 415400 50390 415452 50396
rect 411168 48340 411220 48346
rect 411168 48282 411220 48288
rect 409878 35184 409934 35193
rect 409878 35119 409934 35128
rect 409788 31068 409840 31074
rect 409788 31010 409840 31016
rect 408500 25628 408552 25634
rect 408500 25570 408552 25576
rect 408512 7682 408540 25570
rect 408500 7676 408552 7682
rect 408500 7618 408552 7624
rect 409696 7676 409748 7682
rect 409696 7618 409748 7624
rect 407302 6352 407358 6361
rect 407302 6287 407358 6296
rect 406384 3868 406436 3874
rect 406384 3810 406436 3816
rect 407316 480 407344 6287
rect 408500 4072 408552 4078
rect 408500 4014 408552 4020
rect 408512 480 408540 4014
rect 409708 480 409736 7618
rect 409800 4078 409828 31010
rect 409892 29209 409920 35119
rect 409878 29200 409934 29209
rect 409878 29135 409934 29144
rect 411180 28966 411208 48282
rect 414018 29064 414074 29073
rect 414018 28999 414074 29008
rect 411168 28960 411220 28966
rect 411168 28902 411220 28908
rect 411352 28960 411404 28966
rect 411352 28902 411404 28908
rect 411364 19417 411392 28902
rect 411166 19408 411222 19417
rect 411166 19343 411222 19352
rect 411350 19408 411406 19417
rect 411350 19343 411406 19352
rect 411180 19310 411208 19343
rect 414032 19310 414060 28999
rect 411168 19304 411220 19310
rect 411168 19246 411220 19252
rect 414020 19304 414072 19310
rect 414020 19246 414072 19252
rect 414480 19304 414532 19310
rect 414480 19246 414532 19252
rect 412548 15904 412600 15910
rect 412548 15846 412600 15852
rect 411168 9784 411220 9790
rect 411168 9726 411220 9732
rect 411180 9654 411208 9726
rect 411168 9648 411220 9654
rect 411168 9590 411220 9596
rect 412560 4078 412588 15846
rect 412640 14816 412692 14822
rect 412640 14758 412692 14764
rect 412652 12442 412680 14758
rect 412640 12436 412692 12442
rect 412640 12378 412692 12384
rect 413284 12436 413336 12442
rect 413284 12378 413336 12384
rect 409788 4072 409840 4078
rect 409788 4014 409840 4020
rect 412088 4072 412140 4078
rect 412088 4014 412140 4020
rect 412548 4072 412600 4078
rect 412548 4014 412600 4020
rect 410892 604 410944 610
rect 410892 546 410944 552
rect 410904 480 410932 546
rect 412100 480 412128 4014
rect 413296 480 413324 12378
rect 414492 480 414520 19246
rect 415398 6624 415454 6633
rect 415398 6559 415454 6568
rect 415412 6089 415440 6559
rect 415398 6080 415454 6089
rect 415398 6015 415454 6024
rect 416700 3126 416728 102614
rect 483018 102232 483074 102241
rect 483018 102167 483074 102176
rect 418172 102054 418554 102082
rect 418172 71058 418200 102054
rect 419448 100904 419500 100910
rect 419448 100846 419500 100852
rect 419460 100298 419488 100846
rect 419448 100292 419500 100298
rect 419448 100234 419500 100240
rect 419448 99204 419500 99210
rect 419448 99146 419500 99152
rect 418160 71052 418212 71058
rect 418160 70994 418212 71000
rect 416780 14680 416832 14686
rect 416780 14622 416832 14628
rect 416792 7682 416820 14622
rect 416780 7676 416832 7682
rect 416780 7618 416832 7624
rect 417976 7676 418028 7682
rect 417976 7618 418028 7624
rect 416872 6588 416924 6594
rect 416872 6530 416924 6536
rect 415676 3120 415728 3126
rect 415676 3062 415728 3068
rect 416688 3120 416740 3126
rect 416688 3062 416740 3068
rect 415688 480 415716 3062
rect 416884 480 416912 6530
rect 417988 480 418016 7618
rect 419460 3482 419488 99146
rect 419540 56024 419592 56030
rect 419540 55966 419592 55972
rect 419184 3454 419488 3482
rect 419552 3482 419580 55966
rect 420932 28422 420960 102068
rect 423416 102054 423522 102082
rect 425914 102054 426388 102082
rect 423416 96665 423444 102054
rect 423402 96656 423458 96665
rect 423402 96591 423458 96600
rect 423586 96656 423642 96665
rect 423586 96591 423642 96600
rect 422206 82104 422262 82113
rect 422206 82039 422262 82048
rect 420920 28416 420972 28422
rect 420920 28358 420972 28364
rect 419552 3454 420408 3482
rect 419184 480 419212 3454
rect 420380 480 420408 3454
rect 422220 3398 422248 82039
rect 423600 28422 423628 96591
rect 425060 44940 425112 44946
rect 425060 44882 425112 44888
rect 423588 28416 423640 28422
rect 423588 28358 423640 28364
rect 424966 6624 425022 6633
rect 424966 6559 425022 6568
rect 423956 6520 424008 6526
rect 423956 6462 424008 6468
rect 422760 6452 422812 6458
rect 422760 6394 422812 6400
rect 421564 3392 421616 3398
rect 421564 3334 421616 3340
rect 422208 3392 422260 3398
rect 422208 3334 422260 3340
rect 421576 480 421604 3334
rect 422772 480 422800 6394
rect 423968 480 423996 6462
rect 424980 6089 425008 6559
rect 424966 6080 425022 6089
rect 424966 6015 425022 6024
rect 425072 3398 425100 44882
rect 426360 13122 426388 102054
rect 427832 102054 428306 102082
rect 430592 102054 430882 102082
rect 431972 102054 433274 102082
rect 434732 102054 435850 102082
rect 437492 102054 438242 102082
rect 426438 66872 426494 66881
rect 426438 66807 426494 66816
rect 426348 13116 426400 13122
rect 426348 13058 426400 13064
rect 425150 6624 425206 6633
rect 425150 6559 425206 6568
rect 425060 3392 425112 3398
rect 425060 3334 425112 3340
rect 425164 480 425192 6559
rect 426348 3392 426400 3398
rect 426348 3334 426400 3340
rect 426452 3346 426480 66807
rect 427832 15910 427860 102054
rect 429200 46300 429252 46306
rect 429200 46242 429252 46248
rect 427820 15904 427872 15910
rect 427820 15846 427872 15852
rect 427820 14612 427872 14618
rect 427820 14554 427872 14560
rect 427832 3346 427860 14554
rect 429212 3346 429240 46242
rect 430592 29782 430620 102054
rect 431972 57254 432000 102054
rect 433248 93764 433300 93770
rect 433248 93706 433300 93712
rect 431960 57248 432012 57254
rect 431960 57190 432012 57196
rect 430580 29776 430632 29782
rect 430580 29718 430632 29724
rect 433260 6050 433288 93706
rect 433340 65680 433392 65686
rect 433340 65622 433392 65628
rect 432328 6044 432380 6050
rect 432328 5986 432380 5992
rect 433248 6044 433300 6050
rect 433248 5986 433300 5992
rect 431132 3868 431184 3874
rect 431132 3810 431184 3816
rect 426360 480 426388 3334
rect 426452 3318 427584 3346
rect 427832 3318 428780 3346
rect 429212 3318 429976 3346
rect 427556 480 427584 3318
rect 428752 480 428780 3318
rect 429948 480 429976 3318
rect 431144 480 431172 3810
rect 432340 480 432368 5986
rect 433352 3398 433380 65622
rect 433430 47560 433486 47569
rect 433430 47495 433486 47504
rect 433444 3482 433472 47495
rect 434732 6662 434760 102054
rect 436008 91928 436060 91934
rect 436008 91870 436060 91876
rect 434720 6656 434772 6662
rect 434720 6598 434772 6604
rect 433444 3454 433564 3482
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433536 480 433564 3454
rect 434628 3392 434680 3398
rect 436020 3346 436048 91870
rect 436100 37936 436152 37942
rect 436100 37878 436152 37884
rect 434628 3334 434680 3340
rect 434640 480 434668 3334
rect 435836 3318 436048 3346
rect 436112 3346 436140 37878
rect 437492 10334 437520 102054
rect 439504 101584 439556 101590
rect 439504 101526 439556 101532
rect 437570 71088 437626 71097
rect 437570 71023 437626 71032
rect 437480 10328 437532 10334
rect 437480 10270 437532 10276
rect 437584 3346 437612 71023
rect 438122 5808 438178 5817
rect 438122 5743 438124 5752
rect 438176 5743 438178 5752
rect 438124 5714 438176 5720
rect 439516 3874 439544 101526
rect 440804 100298 440832 102068
rect 443012 102054 443210 102082
rect 445496 102054 445602 102082
rect 448178 102054 448468 102082
rect 450570 102054 451228 102082
rect 440792 100292 440844 100298
rect 440792 100234 440844 100240
rect 440148 96416 440200 96422
rect 440148 96358 440200 96364
rect 439504 3868 439556 3874
rect 439504 3810 439556 3816
rect 440160 3398 440188 96358
rect 441620 40792 441672 40798
rect 441620 40734 441672 40740
rect 440240 28416 440292 28422
rect 440240 28358 440292 28364
rect 439412 3392 439464 3398
rect 436112 3318 437060 3346
rect 437584 3318 438256 3346
rect 439412 3334 439464 3340
rect 440148 3392 440200 3398
rect 440148 3334 440200 3340
rect 440252 3346 440280 28358
rect 441632 3346 441660 40734
rect 443012 7614 443040 102054
rect 445496 96665 445524 102054
rect 445482 96656 445538 96665
rect 445482 96591 445538 96600
rect 445666 96656 445722 96665
rect 445666 96591 445722 96600
rect 444380 91792 444432 91798
rect 444380 91734 444432 91740
rect 444196 9104 444248 9110
rect 444196 9046 444248 9052
rect 443000 7608 443052 7614
rect 443000 7550 443052 7556
rect 442906 5808 442962 5817
rect 442906 5743 442908 5752
rect 442960 5743 442962 5752
rect 442908 5714 442960 5720
rect 443000 3868 443052 3874
rect 443000 3810 443052 3816
rect 435836 480 435864 3318
rect 437032 480 437060 3318
rect 438228 480 438256 3318
rect 439424 480 439452 3334
rect 440252 3318 440648 3346
rect 441632 3318 441844 3346
rect 440620 480 440648 3318
rect 441816 480 441844 3318
rect 443012 480 443040 3810
rect 444208 480 444236 9046
rect 444392 3346 444420 91734
rect 445680 67538 445708 96591
rect 445760 69692 445812 69698
rect 445760 69634 445812 69640
rect 445588 67510 445708 67538
rect 445588 58002 445616 67510
rect 445576 57996 445628 58002
rect 445576 57938 445628 57944
rect 445668 57996 445720 58002
rect 445668 57938 445720 57944
rect 445680 48226 445708 57938
rect 445588 48198 445708 48226
rect 445588 38690 445616 48198
rect 445576 38684 445628 38690
rect 445576 38626 445628 38632
rect 445668 38684 445720 38690
rect 445668 38626 445720 38632
rect 445680 28914 445708 38626
rect 445588 28886 445708 28914
rect 445588 19378 445616 28886
rect 445576 19372 445628 19378
rect 445576 19314 445628 19320
rect 445668 19372 445720 19378
rect 445668 19314 445720 19320
rect 445680 9586 445708 19314
rect 445668 9580 445720 9586
rect 445668 9522 445720 9528
rect 444392 3318 445432 3346
rect 445404 480 445432 3318
rect 445772 2242 445800 69634
rect 448440 15910 448468 102054
rect 448518 86184 448574 86193
rect 448518 86119 448574 86128
rect 448428 15904 448480 15910
rect 448428 15846 448480 15852
rect 448532 12442 448560 86119
rect 451200 33862 451228 102054
rect 452672 102054 453146 102082
rect 451280 83496 451332 83502
rect 451280 83438 451332 83444
rect 451188 33856 451240 33862
rect 451188 33798 451240 33804
rect 449164 20052 449216 20058
rect 449164 19994 449216 20000
rect 448520 12436 448572 12442
rect 448520 12378 448572 12384
rect 448980 12436 449032 12442
rect 448980 12378 449032 12384
rect 447416 7676 447468 7682
rect 447416 7618 447468 7624
rect 447046 5808 447102 5817
rect 447102 5766 447272 5794
rect 447046 5743 447102 5752
rect 447244 5681 447272 5766
rect 447230 5672 447286 5681
rect 447230 5607 447286 5616
rect 447428 4962 447456 7618
rect 447784 6588 447836 6594
rect 447784 6530 447836 6536
rect 447416 4956 447468 4962
rect 447416 4898 447468 4904
rect 445760 2236 445812 2242
rect 445760 2178 445812 2184
rect 446588 2236 446640 2242
rect 446588 2178 446640 2184
rect 446600 480 446628 2178
rect 447796 480 447824 6530
rect 448992 480 449020 12378
rect 449176 7682 449204 19994
rect 450544 17400 450596 17406
rect 450544 17342 450596 17348
rect 449164 7676 449216 7682
rect 449164 7618 449216 7624
rect 450556 4894 450584 17342
rect 451292 7614 451320 83438
rect 452568 22228 452620 22234
rect 452568 22170 452620 22176
rect 452580 20058 452608 22170
rect 452568 20052 452620 20058
rect 452568 19994 452620 20000
rect 452672 17338 452700 102054
rect 453948 101652 454000 101658
rect 453948 101594 454000 101600
rect 452660 17332 452712 17338
rect 452660 17274 452712 17280
rect 451280 7608 451332 7614
rect 451280 7550 451332 7556
rect 452476 7608 452528 7614
rect 452476 7550 452528 7556
rect 450544 4888 450596 4894
rect 450544 4830 450596 4836
rect 451370 3768 451426 3777
rect 451370 3703 451426 3712
rect 450174 3632 450230 3641
rect 450174 3567 450230 3576
rect 450188 480 450216 3567
rect 451384 1850 451412 3703
rect 451292 1822 451412 1850
rect 451292 480 451320 1822
rect 452488 480 452516 7550
rect 453960 2854 453988 101594
rect 455524 100298 455552 102068
rect 456812 102054 458114 102082
rect 459572 102054 460506 102082
rect 462332 102054 462898 102082
rect 465092 102054 465474 102082
rect 455512 100292 455564 100298
rect 455512 100234 455564 100240
rect 456708 100292 456760 100298
rect 456708 100234 456760 100240
rect 456616 96552 456668 96558
rect 456616 96494 456668 96500
rect 454038 90536 454094 90545
rect 454038 90471 454094 90480
rect 454052 12442 454080 90471
rect 456064 44056 456116 44062
rect 456064 43998 456116 44004
rect 456076 22234 456104 43998
rect 456064 22228 456116 22234
rect 456064 22170 456116 22176
rect 455420 22160 455472 22166
rect 455420 22102 455472 22108
rect 455432 20754 455460 22102
rect 455340 20726 455460 20754
rect 455340 17406 455368 20726
rect 455328 17400 455380 17406
rect 455328 17342 455380 17348
rect 454040 12436 454092 12442
rect 454040 12378 454092 12384
rect 454868 12436 454920 12442
rect 454868 12378 454920 12384
rect 453672 2848 453724 2854
rect 453672 2790 453724 2796
rect 453948 2848 454000 2854
rect 453948 2790 454000 2796
rect 453684 480 453712 2790
rect 454880 480 454908 12378
rect 456628 4078 456656 96494
rect 456720 4962 456748 100234
rect 456812 60178 456840 102054
rect 456800 60172 456852 60178
rect 456800 60114 456852 60120
rect 458178 59936 458234 59945
rect 458178 59871 458234 59880
rect 457444 30252 457496 30258
rect 457444 30194 457496 30200
rect 457456 22166 457484 30194
rect 457444 22160 457496 22166
rect 457444 22102 457496 22108
rect 456800 19984 456852 19990
rect 456800 19926 456852 19932
rect 456708 4956 456760 4962
rect 456708 4898 456760 4904
rect 456064 4072 456116 4078
rect 456064 4014 456116 4020
rect 456616 4072 456668 4078
rect 456616 4014 456668 4020
rect 456076 480 456104 4014
rect 456812 3346 456840 19926
rect 457444 11008 457496 11014
rect 457444 10950 457496 10956
rect 457456 5030 457484 10950
rect 457444 5024 457496 5030
rect 457444 4966 457496 4972
rect 458192 3346 458220 59871
rect 458272 34536 458324 34542
rect 458272 34478 458324 34484
rect 458284 30258 458312 34478
rect 458272 30252 458324 30258
rect 458272 30194 458324 30200
rect 459572 16114 459600 102054
rect 461584 49700 461636 49706
rect 461584 49642 461636 49648
rect 461596 44198 461624 49642
rect 461584 44192 461636 44198
rect 461584 44134 461636 44140
rect 460204 41472 460256 41478
rect 460204 41414 460256 41420
rect 459560 16108 459612 16114
rect 459560 16050 459612 16056
rect 459560 14544 459612 14550
rect 459560 14486 459612 14492
rect 459572 3398 459600 14486
rect 459652 6656 459704 6662
rect 459652 6598 459704 6604
rect 459560 3392 459612 3398
rect 456812 3318 457300 3346
rect 458192 3318 458496 3346
rect 459560 3334 459612 3340
rect 457272 480 457300 3318
rect 458468 480 458496 3318
rect 459664 480 459692 6598
rect 460216 4826 460244 41414
rect 461584 39908 461636 39914
rect 461584 39850 461636 39856
rect 461596 34542 461624 39850
rect 461584 34536 461636 34542
rect 461584 34478 461636 34484
rect 460940 32428 460992 32434
rect 460940 32370 460992 32376
rect 460204 4820 460256 4826
rect 460204 4762 460256 4768
rect 460952 3482 460980 32370
rect 462332 25702 462360 102054
rect 463608 97504 463660 97510
rect 463608 97446 463660 97452
rect 462412 57860 462464 57866
rect 462412 57802 462464 57808
rect 462424 49706 462452 57802
rect 462412 49700 462464 49706
rect 462412 49642 462464 49648
rect 462688 43580 462740 43586
rect 462688 43522 462740 43528
rect 462700 41478 462728 43522
rect 462688 41472 462740 41478
rect 462688 41414 462740 41420
rect 462964 34536 463016 34542
rect 462964 34478 463016 34484
rect 462320 25696 462372 25702
rect 462320 25638 462372 25644
rect 462976 11014 463004 34478
rect 462964 11008 463016 11014
rect 462964 10950 463016 10956
rect 462320 8900 462372 8906
rect 462320 8842 462372 8848
rect 462332 8242 462360 8842
rect 462240 8214 462360 8242
rect 462240 5098 462268 8214
rect 462228 5092 462280 5098
rect 462228 5034 462280 5040
rect 463620 3482 463648 97446
rect 464344 53848 464396 53854
rect 464344 53790 464396 53796
rect 464356 43586 464384 53790
rect 464344 43580 464396 43586
rect 464344 43522 464396 43528
rect 463792 42832 463844 42838
rect 463792 42774 463844 42780
rect 463804 39914 463832 42774
rect 463792 39908 463844 39914
rect 463792 39850 463844 39856
rect 465092 11966 465120 102054
rect 467852 100774 467880 102068
rect 469232 102054 470442 102082
rect 472834 102054 473308 102082
rect 467840 100768 467892 100774
rect 467840 100710 467892 100716
rect 469128 99340 469180 99346
rect 469128 99282 469180 99288
rect 468944 69080 468996 69086
rect 468944 69022 468996 69028
rect 467104 67516 467156 67522
rect 467104 67458 467156 67464
rect 465172 62144 465224 62150
rect 465172 62086 465224 62092
rect 465184 57866 465212 62086
rect 465172 57860 465224 57866
rect 465172 57802 465224 57808
rect 465816 47932 465868 47938
rect 465816 47874 465868 47880
rect 465828 42838 465856 47874
rect 465816 42832 465868 42838
rect 465816 42774 465868 42780
rect 465724 40112 465776 40118
rect 465724 40054 465776 40060
rect 465736 34542 465764 40054
rect 465724 34536 465776 34542
rect 465724 34478 465776 34484
rect 467116 23526 467144 67458
rect 468956 67250 468984 69022
rect 467196 67244 467248 67250
rect 467196 67186 467248 67192
rect 468944 67244 468996 67250
rect 468944 67186 468996 67192
rect 467208 62150 467236 67186
rect 467196 62144 467248 62150
rect 467196 62086 467248 62092
rect 467748 60104 467800 60110
rect 467748 60046 467800 60052
rect 465724 23520 465776 23526
rect 465724 23462 465776 23468
rect 467104 23520 467156 23526
rect 467104 23462 467156 23468
rect 465080 11960 465132 11966
rect 465080 11902 465132 11908
rect 465736 8906 465764 23462
rect 465724 8900 465776 8906
rect 465724 8842 465776 8848
rect 467760 4078 467788 60046
rect 467840 57792 467892 57798
rect 467840 57734 467892 57740
rect 467852 53854 467880 57734
rect 467840 53848 467892 53854
rect 467840 53790 467892 53796
rect 467840 52488 467892 52494
rect 467840 52430 467892 52436
rect 467852 47938 467880 52430
rect 467840 47932 467892 47938
rect 467840 47874 467892 47880
rect 468482 5944 468538 5953
rect 468482 5879 468538 5888
rect 468496 5545 468524 5879
rect 468482 5536 468538 5545
rect 468482 5471 468538 5480
rect 467932 4956 467984 4962
rect 467932 4898 467984 4904
rect 466828 4072 466880 4078
rect 466828 4014 466880 4020
rect 467748 4072 467800 4078
rect 467748 4014 467800 4020
rect 464434 3904 464490 3913
rect 464434 3839 464490 3848
rect 460952 3454 462084 3482
rect 460848 3392 460900 3398
rect 460848 3334 460900 3340
rect 460860 480 460888 3334
rect 462056 480 462084 3454
rect 463252 3454 463648 3482
rect 463252 480 463280 3454
rect 464448 480 464476 3839
rect 465630 2816 465686 2825
rect 465630 2751 465686 2760
rect 465644 480 465672 2751
rect 466840 480 466868 4014
rect 467944 480 467972 4898
rect 469140 480 469168 99282
rect 469232 31074 469260 102054
rect 473280 86290 473308 102054
rect 475396 100298 475424 102068
rect 475384 100292 475436 100298
rect 475384 100234 475436 100240
rect 477788 99958 477816 102068
rect 480076 101856 480128 101862
rect 480076 101798 480128 101804
rect 478788 100088 478840 100094
rect 478788 100030 478840 100036
rect 477776 99952 477828 99958
rect 477776 99894 477828 99900
rect 478696 99952 478748 99958
rect 478696 99894 478748 99900
rect 473268 86284 473320 86290
rect 473268 86226 473320 86232
rect 477500 85604 477552 85610
rect 477500 85546 477552 85552
rect 476120 84176 476172 84182
rect 476120 84118 476172 84124
rect 476132 80102 476160 84118
rect 477512 81546 477540 85546
rect 477420 81518 477540 81546
rect 474648 80096 474700 80102
rect 474648 80038 474700 80044
rect 476120 80096 476172 80102
rect 476120 80038 476172 80044
rect 473268 79348 473320 79354
rect 473268 79290 473320 79296
rect 471244 78124 471296 78130
rect 471244 78066 471296 78072
rect 470600 76764 470652 76770
rect 470600 76706 470652 76712
rect 470612 73250 470640 76706
rect 470520 73222 470640 73250
rect 469312 72004 469364 72010
rect 469312 71946 469364 71952
rect 469324 67522 469352 71946
rect 469864 69284 469916 69290
rect 469864 69226 469916 69232
rect 469312 67516 469364 67522
rect 469312 67458 469364 67464
rect 469876 57798 469904 69226
rect 470520 69086 470548 73222
rect 471256 72010 471284 78066
rect 473280 76770 473308 79290
rect 474660 78130 474688 80038
rect 477420 79354 477448 81518
rect 477408 79348 477460 79354
rect 477408 79290 477460 79296
rect 474648 78124 474700 78130
rect 474648 78066 474700 78072
rect 475384 77580 475436 77586
rect 475384 77522 475436 77528
rect 473268 76764 473320 76770
rect 473268 76706 473320 76712
rect 471244 72004 471296 72010
rect 471244 71946 471296 71952
rect 475396 70650 475424 77522
rect 472440 70644 472492 70650
rect 472440 70586 472492 70592
rect 475384 70644 475436 70650
rect 475384 70586 475436 70592
rect 472452 69290 472480 70586
rect 472440 69284 472492 69290
rect 472440 69226 472492 69232
rect 470508 69080 470560 69086
rect 470508 69022 470560 69028
rect 476764 62688 476816 62694
rect 476764 62630 476816 62636
rect 469864 57792 469916 57798
rect 469864 57734 469916 57740
rect 472900 53916 472952 53922
rect 472900 53858 472952 53864
rect 472912 52494 472940 53858
rect 476776 52494 476804 62630
rect 472900 52488 472952 52494
rect 472900 52430 472952 52436
rect 474004 52488 474056 52494
rect 474004 52430 474056 52436
rect 476764 52488 476816 52494
rect 476764 52430 476816 52436
rect 474016 42090 474044 52430
rect 476120 51740 476172 51746
rect 476120 51682 476172 51688
rect 469312 42084 469364 42090
rect 469312 42026 469364 42032
rect 474004 42084 474056 42090
rect 474004 42026 474056 42032
rect 469324 40118 469352 42026
rect 469312 40112 469364 40118
rect 469312 40054 469364 40060
rect 469220 31068 469272 31074
rect 469220 31010 469272 31016
rect 473360 21412 473412 21418
rect 473360 21354 473412 21360
rect 473372 12442 473400 21354
rect 473360 12436 473412 12442
rect 473360 12378 473412 12384
rect 473912 12436 473964 12442
rect 473912 12378 473964 12384
rect 472716 12028 472768 12034
rect 472716 11970 472768 11976
rect 471518 6760 471574 6769
rect 471518 6695 471574 6704
rect 470324 4004 470376 4010
rect 470324 3946 470376 3952
rect 470336 480 470364 3946
rect 471532 480 471560 6695
rect 472728 480 472756 11970
rect 473924 480 473952 12378
rect 475108 6724 475160 6730
rect 475108 6666 475160 6672
rect 475120 480 475148 6666
rect 476132 3482 476160 51682
rect 478708 21418 478736 99894
rect 478696 21412 478748 21418
rect 478696 21354 478748 21360
rect 477500 3936 477552 3942
rect 477500 3878 477552 3884
rect 476132 3454 476344 3482
rect 476316 480 476344 3454
rect 477512 480 477540 3878
rect 478800 3482 478828 100030
rect 480088 96370 480116 101798
rect 480180 96529 480208 102068
rect 481652 102054 482770 102082
rect 480166 96520 480222 96529
rect 480166 96455 480222 96464
rect 480088 96342 480208 96370
rect 478880 81456 478932 81462
rect 478880 81398 478932 81404
rect 478892 77586 478920 81398
rect 478880 77580 478932 77586
rect 478880 77522 478932 77528
rect 478880 56024 478932 56030
rect 478880 55966 478932 55972
rect 478892 53922 478920 55966
rect 478880 53916 478932 53922
rect 478880 53858 478932 53864
rect 480180 3482 480208 96342
rect 480720 91112 480772 91118
rect 480720 91054 480772 91060
rect 480732 85610 480760 91054
rect 480720 85604 480772 85610
rect 480720 85546 480772 85552
rect 481088 82884 481140 82890
rect 481088 82826 481140 82832
rect 481100 81462 481128 82826
rect 481088 81456 481140 81462
rect 481088 81398 481140 81404
rect 481652 77994 481680 102054
rect 483032 97345 483060 102167
rect 492862 102096 492918 102105
rect 484412 102054 485162 102082
rect 487172 102054 487738 102082
rect 489932 102054 490130 102082
rect 484308 101720 484360 101726
rect 484308 101662 484360 101668
rect 483018 97336 483074 97345
rect 483018 97271 483074 97280
rect 484216 95056 484268 95062
rect 484216 94998 484268 95004
rect 481732 94988 481784 94994
rect 481732 94930 481784 94936
rect 481744 91118 481772 94930
rect 481732 91112 481784 91118
rect 481732 91054 481784 91060
rect 483020 91112 483072 91118
rect 483020 91054 483072 91060
rect 482284 88528 482336 88534
rect 482284 88470 482336 88476
rect 481640 77988 481692 77994
rect 481640 77930 481692 77936
rect 481638 77888 481694 77897
rect 481638 77823 481694 77832
rect 480904 75880 480956 75886
rect 480904 75822 480956 75828
rect 480916 62694 480944 75822
rect 480904 62688 480956 62694
rect 480904 62630 480956 62636
rect 481088 6724 481140 6730
rect 481088 6666 481140 6672
rect 478708 3454 478828 3482
rect 479904 3454 480208 3482
rect 478708 480 478736 3454
rect 479904 480 479932 3454
rect 481100 480 481128 6666
rect 481652 3346 481680 77823
rect 482296 75886 482324 88470
rect 483032 85626 483060 91054
rect 484228 88534 484256 94998
rect 484216 88528 484268 88534
rect 484216 88470 484268 88476
rect 483756 86964 483808 86970
rect 483756 86906 483808 86912
rect 482940 85598 483060 85626
rect 482940 84250 482968 85598
rect 482928 84244 482980 84250
rect 482928 84186 482980 84192
rect 483768 82890 483796 86906
rect 483756 82884 483808 82890
rect 483756 82826 483808 82832
rect 483664 78260 483716 78266
rect 483664 78202 483716 78208
rect 482284 75880 482336 75886
rect 482284 75822 482336 75828
rect 483676 60790 483704 78202
rect 482008 60784 482060 60790
rect 482008 60726 482060 60732
rect 483664 60784 483716 60790
rect 483664 60726 483716 60732
rect 482020 56030 482048 60726
rect 482008 56024 482060 56030
rect 482008 55966 482060 55972
rect 481824 5976 481876 5982
rect 481822 5944 481824 5953
rect 481876 5944 481878 5953
rect 481822 5879 481878 5888
rect 484320 3398 484348 101662
rect 484412 29714 484440 102054
rect 487068 101788 487120 101794
rect 487068 101730 487120 101736
rect 486976 99272 487028 99278
rect 486976 99214 487028 99220
rect 484490 96656 484546 96665
rect 484490 96591 484546 96600
rect 484504 94994 484532 96591
rect 484492 94988 484544 94994
rect 484492 94930 484544 94936
rect 484492 88664 484544 88670
rect 484492 88606 484544 88612
rect 484504 86970 484532 88606
rect 484492 86964 484544 86970
rect 484492 86906 484544 86912
rect 485504 82884 485556 82890
rect 485504 82826 485556 82832
rect 485516 78266 485544 82826
rect 485504 78260 485556 78266
rect 485504 78202 485556 78208
rect 484400 29708 484452 29714
rect 484400 29650 484452 29656
rect 484400 21412 484452 21418
rect 484400 21354 484452 21360
rect 483480 3392 483532 3398
rect 481652 3318 482324 3346
rect 483480 3334 483532 3340
rect 484308 3392 484360 3398
rect 484308 3334 484360 3340
rect 484412 3346 484440 21354
rect 486884 12436 486936 12442
rect 486884 12378 486936 12384
rect 485780 4072 485832 4078
rect 485780 4014 485832 4020
rect 482296 480 482324 3318
rect 483492 480 483520 3334
rect 484412 3318 484624 3346
rect 484596 480 484624 3318
rect 485792 480 485820 4014
rect 486896 3890 486924 12378
rect 486988 4078 487016 99214
rect 487080 12442 487108 101730
rect 487172 53106 487200 102054
rect 488448 101924 488500 101930
rect 488448 101866 488500 101872
rect 487804 97572 487856 97578
rect 487804 97514 487856 97520
rect 487816 95062 487844 97514
rect 487804 95056 487856 95062
rect 487804 94998 487856 95004
rect 487804 93900 487856 93906
rect 487804 93842 487856 93848
rect 487816 88670 487844 93842
rect 487804 88664 487856 88670
rect 487804 88606 487856 88612
rect 487252 86692 487304 86698
rect 487252 86634 487304 86640
rect 487264 82890 487292 86634
rect 487252 82884 487304 82890
rect 487252 82826 487304 82832
rect 487160 53100 487212 53106
rect 487160 53042 487212 53048
rect 488460 12510 488488 101866
rect 488630 96656 488686 96665
rect 488630 96591 488686 96600
rect 488540 91996 488592 92002
rect 488540 91938 488592 91944
rect 488552 86698 488580 91938
rect 488644 91118 488672 96591
rect 488632 91112 488684 91118
rect 488632 91054 488684 91060
rect 488540 86692 488592 86698
rect 488540 86634 488592 86640
rect 489932 72554 489960 102054
rect 491300 97640 491352 97646
rect 491300 97582 491352 97588
rect 491312 93906 491340 97582
rect 491300 93900 491352 93906
rect 491300 93842 491352 93848
rect 489920 72548 489972 72554
rect 489920 72490 489972 72496
rect 492692 46238 492720 102068
rect 495254 102096 495310 102105
rect 492862 102031 492918 102040
rect 494072 102054 495098 102082
rect 492876 96121 492904 102031
rect 492862 96112 492918 96121
rect 492862 96047 492918 96056
rect 492772 94716 492824 94722
rect 492772 94658 492824 94664
rect 492784 92002 492812 94658
rect 492772 91996 492824 92002
rect 492772 91938 492824 91944
rect 494072 60110 494100 102054
rect 495254 102031 495310 102040
rect 496832 102054 497490 102082
rect 494150 101960 494206 101969
rect 494150 101895 494206 101904
rect 494060 60104 494112 60110
rect 494060 60046 494112 60052
rect 492680 46232 492732 46238
rect 492680 46174 492732 46180
rect 492680 42152 492732 42158
rect 492680 42094 492732 42100
rect 491300 28348 491352 28354
rect 491300 28290 491352 28296
rect 488448 12504 488500 12510
rect 488448 12446 488500 12452
rect 487068 12436 487120 12442
rect 487068 12378 487120 12384
rect 488172 9716 488224 9722
rect 488172 9658 488224 9664
rect 486976 4072 487028 4078
rect 486976 4014 487028 4020
rect 486896 3862 487016 3890
rect 486988 480 487016 3862
rect 488184 480 488212 9658
rect 491208 5976 491260 5982
rect 491206 5944 491208 5953
rect 491260 5944 491262 5953
rect 491206 5879 491262 5888
rect 489366 4040 489422 4049
rect 489366 3975 489422 3984
rect 489380 480 489408 3975
rect 490562 3768 490618 3777
rect 490562 3703 490618 3712
rect 490576 480 490604 3703
rect 491312 626 491340 28290
rect 491312 598 491800 626
rect 492692 610 492720 42094
rect 494060 40724 494112 40730
rect 494060 40666 494112 40672
rect 494072 7614 494100 40666
rect 494060 7608 494112 7614
rect 494060 7550 494112 7556
rect 494164 4010 494192 101895
rect 495268 101454 495296 102031
rect 495256 101448 495308 101454
rect 495256 101390 495308 101396
rect 494704 99408 494756 99414
rect 494704 99350 494756 99356
rect 494716 11898 494744 99350
rect 496832 69766 496860 102054
rect 499488 101992 499540 101998
rect 499488 101934 499540 101940
rect 499118 100736 499174 100745
rect 499118 100671 499174 100680
rect 496820 69760 496872 69766
rect 496820 69702 496872 69708
rect 499132 67697 499160 100671
rect 499118 67688 499174 67697
rect 499118 67623 499174 67632
rect 499210 67008 499266 67017
rect 499210 66943 499266 66952
rect 499224 60081 499252 66943
rect 499210 60072 499266 60081
rect 499210 60007 499266 60016
rect 499210 55176 499266 55185
rect 499210 55111 499266 55120
rect 499224 45801 499252 55111
rect 499210 45792 499266 45801
rect 499210 45727 499266 45736
rect 496358 45520 496414 45529
rect 496358 45455 496414 45464
rect 499210 45520 499266 45529
rect 499210 45455 499266 45464
rect 496372 40769 496400 45455
rect 499224 40769 499252 45455
rect 496358 40760 496414 40769
rect 496358 40695 496414 40704
rect 499210 40760 499266 40769
rect 499210 40695 499266 40704
rect 495440 33788 495492 33794
rect 495440 33730 495492 33736
rect 494704 11892 494756 11898
rect 494704 11834 494756 11840
rect 495348 7608 495400 7614
rect 495348 7550 495400 7556
rect 494152 4004 494204 4010
rect 494152 3946 494204 3952
rect 494152 3324 494204 3330
rect 494152 3266 494204 3272
rect 491772 480 491800 598
rect 492680 604 492732 610
rect 492680 546 492732 552
rect 492956 604 493008 610
rect 492956 546 493008 552
rect 492968 480 492996 546
rect 494164 480 494192 3266
rect 495360 480 495388 7550
rect 495452 610 495480 33730
rect 498382 28792 498438 28801
rect 498382 28727 498438 28736
rect 498396 21185 498424 28727
rect 498382 21176 498438 21185
rect 498382 21111 498438 21120
rect 499500 4078 499528 101934
rect 500052 99414 500080 102068
rect 500868 101448 500920 101454
rect 500868 101390 500920 101396
rect 500040 99408 500092 99414
rect 500040 99350 500092 99356
rect 500498 87680 500554 87689
rect 500498 87615 500554 87624
rect 500512 82113 500540 87615
rect 500498 82104 500554 82113
rect 500498 82039 500554 82048
rect 500038 45520 500094 45529
rect 500038 45455 500094 45464
rect 500052 39273 500080 45455
rect 500038 39264 500094 39273
rect 500038 39199 500094 39208
rect 498936 4072 498988 4078
rect 498936 4014 498988 4020
rect 499488 4072 499540 4078
rect 499488 4014 499540 4020
rect 497740 4004 497792 4010
rect 497740 3946 497792 3952
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 3946
rect 498948 480 498976 4014
rect 500880 3942 500908 101390
rect 501524 38010 501552 136575
rect 501616 94586 501644 308207
rect 501786 279168 501842 279177
rect 501786 279103 501842 279112
rect 501694 271960 501750 271969
rect 501694 271895 501750 271904
rect 501604 94580 501656 94586
rect 501604 94522 501656 94528
rect 501708 73914 501736 271895
rect 501800 96354 501828 279103
rect 501970 228848 502026 228857
rect 501970 228783 502026 228792
rect 501984 220969 502012 228783
rect 501970 220960 502026 220969
rect 501970 220895 502026 220904
rect 501878 183968 501934 183977
rect 501878 183903 501934 183912
rect 501892 122777 501920 183903
rect 501970 126984 502026 126993
rect 501970 126919 502026 126928
rect 501878 122768 501934 122777
rect 501878 122703 501934 122712
rect 501878 121952 501934 121961
rect 501878 121887 501934 121896
rect 501788 96348 501840 96354
rect 501788 96290 501840 96296
rect 501892 78062 501920 121887
rect 501984 119377 502012 126919
rect 501970 119368 502026 119377
rect 501970 119303 502026 119312
rect 501880 78056 501932 78062
rect 501880 77998 501932 78004
rect 501696 73908 501748 73914
rect 501696 73850 501748 73856
rect 502352 61470 502380 451279
rect 502444 414905 502472 667898
rect 504824 607300 504876 607306
rect 504824 607242 504876 607248
rect 503904 605872 503956 605878
rect 503904 605814 503956 605820
rect 502984 604784 503036 604790
rect 502984 604726 503036 604732
rect 502430 414896 502486 414905
rect 502430 414831 502486 414840
rect 502522 411088 502578 411097
rect 502522 411023 502578 411032
rect 502430 312624 502486 312633
rect 502430 312559 502486 312568
rect 502340 61464 502392 61470
rect 502340 61406 502392 61412
rect 501512 38004 501564 38010
rect 501512 37946 501564 37952
rect 502340 18692 502392 18698
rect 502340 18634 502392 18640
rect 500960 13116 501012 13122
rect 500960 13058 501012 13064
rect 500132 3936 500184 3942
rect 500132 3878 500184 3884
rect 500868 3936 500920 3942
rect 500868 3878 500920 3884
rect 500144 480 500172 3878
rect 500972 610 501000 13058
rect 502352 12442 502380 18634
rect 502340 12436 502392 12442
rect 502340 12378 502392 12384
rect 502444 4690 502472 312559
rect 502536 101862 502564 411023
rect 502996 382974 503024 604726
rect 503812 604716 503864 604722
rect 503812 604658 503864 604664
rect 503720 604512 503772 604518
rect 503720 604454 503772 604460
rect 502984 382968 503036 382974
rect 502984 382910 503036 382916
rect 502614 352608 502670 352617
rect 502614 352543 502670 352552
rect 502524 101856 502576 101862
rect 502524 101798 502576 101804
rect 502628 68406 502656 352543
rect 502706 265024 502762 265033
rect 502706 264959 502762 264968
rect 502720 83570 502748 264959
rect 503626 254416 503682 254425
rect 503626 254351 503682 254360
rect 503640 253881 503668 254351
rect 503626 253872 503682 253881
rect 503626 253807 503682 253816
rect 502890 217696 502946 217705
rect 502890 217631 502946 217640
rect 502798 159216 502854 159225
rect 502798 159151 502854 159160
rect 502708 83564 502760 83570
rect 502708 83506 502760 83512
rect 502616 68400 502668 68406
rect 502616 68342 502668 68348
rect 502812 15978 502840 159151
rect 502904 99346 502932 217631
rect 503732 174049 503760 604454
rect 503824 181257 503852 604658
rect 503916 593881 503944 605814
rect 504836 601390 504864 607242
rect 505744 607232 505796 607238
rect 505744 607174 505796 607180
rect 504824 601384 504876 601390
rect 504824 601326 504876 601332
rect 503996 601316 504048 601322
rect 503996 601258 504048 601264
rect 504008 598330 504036 601258
rect 503996 598324 504048 598330
rect 503996 598266 504048 598272
rect 504364 596216 504416 596222
rect 504364 596158 504416 596164
rect 503902 593872 503958 593881
rect 503902 593807 503958 593816
rect 504376 592770 504404 596158
rect 504376 592742 504496 592770
rect 503904 586560 503956 586566
rect 503902 586528 503904 586537
rect 503956 586528 503958 586537
rect 503902 586463 503958 586472
rect 503902 582720 503958 582729
rect 503902 582655 503958 582664
rect 503916 582418 503944 582655
rect 503904 582412 503956 582418
rect 503904 582354 503956 582360
rect 504468 578270 504496 592742
rect 504364 578264 504416 578270
rect 504364 578206 504416 578212
rect 504456 578264 504508 578270
rect 504456 578206 504508 578212
rect 504376 572830 504404 578206
rect 504454 575648 504510 575657
rect 504454 575583 504510 575592
rect 504364 572824 504416 572830
rect 504364 572766 504416 572772
rect 504272 572688 504324 572694
rect 504272 572630 504324 572636
rect 503902 571840 503958 571849
rect 503902 571775 503958 571784
rect 503916 571402 503944 571775
rect 503904 571396 503956 571402
rect 503904 571338 503956 571344
rect 504284 569922 504312 572630
rect 504362 569936 504418 569945
rect 504284 569894 504362 569922
rect 504362 569871 504418 569880
rect 503902 568304 503958 568313
rect 503902 568239 503958 568248
rect 503916 567254 503944 568239
rect 503904 567248 503956 567254
rect 503904 567190 503956 567196
rect 503902 564496 503958 564505
rect 503902 564431 503904 564440
rect 503956 564431 503958 564440
rect 503904 564402 503956 564408
rect 504364 562964 504416 562970
rect 504364 562906 504416 562912
rect 503902 560960 503958 560969
rect 503902 560895 503958 560904
rect 503916 560318 503944 560895
rect 503904 560312 503956 560318
rect 503904 560254 503956 560260
rect 503904 554736 503956 554742
rect 503904 554678 503956 554684
rect 503916 553625 503944 554678
rect 503902 553616 503958 553625
rect 503902 553551 503958 553560
rect 503902 550080 503958 550089
rect 503902 550015 503958 550024
rect 503916 549302 503944 550015
rect 503904 549296 503956 549302
rect 503904 549238 503956 549244
rect 503902 546272 503958 546281
rect 503902 546207 503958 546216
rect 503916 545222 503944 546207
rect 503904 545216 503956 545222
rect 503904 545158 503956 545164
rect 504376 543810 504404 562906
rect 504468 547194 504496 575583
rect 504546 569936 504602 569945
rect 504546 569871 504602 569880
rect 504560 562970 504588 569871
rect 504548 562964 504600 562970
rect 504548 562906 504600 562912
rect 504456 547188 504508 547194
rect 504456 547130 504508 547136
rect 504376 543782 504496 543810
rect 503902 542736 503958 542745
rect 503902 542671 503958 542680
rect 503916 541686 503944 542671
rect 503904 541680 503956 541686
rect 503904 541622 503956 541628
rect 503902 538928 503958 538937
rect 503902 538863 503958 538872
rect 503916 538286 503944 538863
rect 503904 538280 503956 538286
rect 503904 538222 503956 538228
rect 504468 534206 504496 543782
rect 504456 534200 504508 534206
rect 504456 534142 504508 534148
rect 504376 531350 504404 531381
rect 504364 531344 504416 531350
rect 504416 531292 504496 531298
rect 504364 531286 504496 531292
rect 504376 531282 504496 531286
rect 504376 531276 504508 531282
rect 504376 531270 504456 531276
rect 504456 531218 504508 531224
rect 503902 524512 503958 524521
rect 503902 524447 503904 524456
rect 503956 524447 503958 524456
rect 503904 524418 503956 524424
rect 504456 524340 504508 524346
rect 504456 524282 504508 524288
rect 504468 521642 504496 524282
rect 504376 521614 504496 521642
rect 503902 520704 503958 520713
rect 503902 520639 503958 520648
rect 503916 520334 503944 520639
rect 503904 520328 503956 520334
rect 503904 520270 503956 520276
rect 504376 514826 504404 521614
rect 504364 514820 504416 514826
rect 504364 514762 504416 514768
rect 504364 512032 504416 512038
rect 504364 511974 504416 511980
rect 504376 505170 504404 511974
rect 504364 505164 504416 505170
rect 504364 505106 504416 505112
rect 504456 505028 504508 505034
rect 504456 504970 504508 504976
rect 504468 502330 504496 504970
rect 504376 502302 504496 502330
rect 503902 498944 503958 498953
rect 503902 498879 503958 498888
rect 503916 498234 503944 498879
rect 503904 498228 503956 498234
rect 503904 498170 503956 498176
rect 504376 497554 504404 502302
rect 504180 497548 504232 497554
rect 504180 497490 504232 497496
rect 504364 497548 504416 497554
rect 504364 497490 504416 497496
rect 503902 495136 503958 495145
rect 503902 495071 503958 495080
rect 503916 494086 503944 495071
rect 503904 494080 503956 494086
rect 503904 494022 503956 494028
rect 504192 492697 504220 497490
rect 504178 492688 504234 492697
rect 504178 492623 504234 492632
rect 504362 492688 504418 492697
rect 504362 492623 504418 492632
rect 503902 487792 503958 487801
rect 503902 487727 503958 487736
rect 503916 487218 503944 487727
rect 503904 487212 503956 487218
rect 503904 487154 503956 487160
rect 504376 485858 504404 492623
rect 504364 485852 504416 485858
rect 504364 485794 504416 485800
rect 504456 485716 504508 485722
rect 504456 485658 504508 485664
rect 503902 484256 503958 484265
rect 503902 484191 503958 484200
rect 503916 483070 503944 484191
rect 503904 483064 503956 483070
rect 503904 483006 503956 483012
rect 504468 483002 504496 485658
rect 504456 482996 504508 483002
rect 504456 482938 504508 482944
rect 504640 482996 504692 483002
rect 504640 482938 504692 482944
rect 503902 476912 503958 476921
rect 503902 476847 503958 476856
rect 503916 476134 503944 476847
rect 503904 476128 503956 476134
rect 503904 476070 503956 476076
rect 503904 473408 503956 473414
rect 503902 473376 503904 473385
rect 504652 473385 504680 482938
rect 503956 473376 503958 473385
rect 504454 473376 504510 473385
rect 503902 473311 503958 473320
rect 504376 473334 504454 473362
rect 503902 469568 503958 469577
rect 503902 469503 503958 469512
rect 503916 469266 503944 469503
rect 503904 469260 503956 469266
rect 503904 469202 503956 469208
rect 504376 466478 504404 473334
rect 504454 473311 504510 473320
rect 504638 473376 504694 473385
rect 504638 473311 504694 473320
rect 504364 466472 504416 466478
rect 504364 466414 504416 466420
rect 504456 466404 504508 466410
rect 504456 466346 504508 466352
rect 504468 463690 504496 466346
rect 504180 463684 504232 463690
rect 504180 463626 504232 463632
rect 504456 463684 504508 463690
rect 504456 463626 504508 463632
rect 503902 462224 503958 462233
rect 503902 462159 503958 462168
rect 503916 461582 503944 462159
rect 503904 461576 503956 461582
rect 503904 461518 503956 461524
rect 504192 454073 504220 463626
rect 504178 454064 504234 454073
rect 504178 453999 504234 454008
rect 504362 454064 504418 454073
rect 504362 453999 504418 454008
rect 503902 447808 503958 447817
rect 503902 447743 503958 447752
rect 503916 447166 503944 447743
rect 503904 447160 503956 447166
rect 503904 447102 503956 447108
rect 504376 446978 504404 453999
rect 504376 446950 504496 446978
rect 504468 444378 504496 446950
rect 504456 444372 504508 444378
rect 504456 444314 504508 444320
rect 503902 444000 503958 444009
rect 503902 443935 503958 443944
rect 503916 443018 503944 443935
rect 503904 443012 503956 443018
rect 503904 442954 503956 442960
rect 503902 440464 503958 440473
rect 503902 440399 503958 440408
rect 503916 440298 503944 440399
rect 503904 440292 503956 440298
rect 503904 440234 503956 440240
rect 503902 436656 503958 436665
rect 503902 436591 503958 436600
rect 503916 436150 503944 436591
rect 503904 436144 503956 436150
rect 503904 436086 503956 436092
rect 504364 434784 504416 434790
rect 504364 434726 504416 434732
rect 503902 433120 503958 433129
rect 503902 433055 503958 433064
rect 503916 432546 503944 433055
rect 503904 432540 503956 432546
rect 503904 432482 503956 432488
rect 503902 429312 503958 429321
rect 503902 429247 503958 429256
rect 503916 429214 503944 429247
rect 503904 429208 503956 429214
rect 503904 429150 503956 429156
rect 504376 427854 504404 434726
rect 504364 427848 504416 427854
rect 504364 427790 504416 427796
rect 504456 427780 504508 427786
rect 504456 427722 504508 427728
rect 503902 425776 503958 425785
rect 503902 425711 503958 425720
rect 503916 425134 503944 425711
rect 503904 425128 503956 425134
rect 503904 425070 503956 425076
rect 504468 425066 504496 427722
rect 504456 425060 504508 425066
rect 504456 425002 504508 425008
rect 503902 422240 503958 422249
rect 503902 422175 503958 422184
rect 503916 420986 503944 422175
rect 503904 420980 503956 420986
rect 503904 420922 503956 420928
rect 504364 415472 504416 415478
rect 504364 415414 504416 415420
rect 504376 408542 504404 415414
rect 504364 408536 504416 408542
rect 504364 408478 504416 408484
rect 504456 408400 504508 408406
rect 504456 408342 504508 408348
rect 503902 407552 503958 407561
rect 503902 407487 503958 407496
rect 503916 407182 503944 407487
rect 503904 407176 503956 407182
rect 503904 407118 503956 407124
rect 503902 403744 503958 403753
rect 503902 403679 503958 403688
rect 503916 403034 503944 403679
rect 503904 403028 503956 403034
rect 503904 402970 503956 402976
rect 504468 400926 504496 408342
rect 504456 400920 504508 400926
rect 504456 400862 504508 400868
rect 504640 400920 504692 400926
rect 504640 400862 504692 400868
rect 503902 400208 503958 400217
rect 503902 400143 503958 400152
rect 503916 398886 503944 400143
rect 503904 398880 503956 398886
rect 503904 398822 503956 398828
rect 504652 396137 504680 400862
rect 505098 396672 505154 396681
rect 505098 396607 505154 396616
rect 504454 396128 504510 396137
rect 504376 396086 504454 396114
rect 504376 393310 504404 396086
rect 504454 396063 504510 396072
rect 504638 396128 504694 396137
rect 504638 396063 504694 396072
rect 504364 393304 504416 393310
rect 504364 393246 504416 393252
rect 504456 393304 504508 393310
rect 504456 393246 504508 393252
rect 503902 389328 503958 389337
rect 503902 389263 503958 389272
rect 503916 389230 503944 389263
rect 503904 389224 503956 389230
rect 503904 389166 503956 389172
rect 503902 385520 503958 385529
rect 503902 385455 503958 385464
rect 503916 385082 503944 385455
rect 503904 385076 503956 385082
rect 503904 385018 503956 385024
rect 503902 381984 503958 381993
rect 503902 381919 503958 381928
rect 503916 380934 503944 381919
rect 503904 380928 503956 380934
rect 503904 380870 503956 380876
rect 503904 378208 503956 378214
rect 503902 378176 503904 378185
rect 503956 378176 503958 378185
rect 503902 378111 503958 378120
rect 503904 375352 503956 375358
rect 503904 375294 503956 375300
rect 503916 374649 503944 375294
rect 503902 374640 503958 374649
rect 503902 374575 503958 374584
rect 503902 371104 503958 371113
rect 503902 371039 503958 371048
rect 503810 181248 503866 181257
rect 503810 181183 503866 181192
rect 503810 177440 503866 177449
rect 503810 177375 503866 177384
rect 503718 174040 503774 174049
rect 503718 173975 503774 173984
rect 503720 170808 503772 170814
rect 503720 170750 503772 170756
rect 503732 170105 503760 170750
rect 503718 170096 503774 170105
rect 503718 170031 503774 170040
rect 503718 166560 503774 166569
rect 503718 166495 503774 166504
rect 503732 165646 503760 166495
rect 503720 165640 503772 165646
rect 503720 165582 503772 165588
rect 503718 151872 503774 151881
rect 503718 151807 503720 151816
rect 503772 151807 503774 151816
rect 503720 151778 503772 151784
rect 503718 148064 503774 148073
rect 503718 147999 503774 148008
rect 503074 133648 503130 133657
rect 503074 133583 503130 133592
rect 503088 133074 503116 133583
rect 503076 133068 503128 133074
rect 503076 133010 503128 133016
rect 503258 111616 503314 111625
rect 503258 111551 503314 111560
rect 503272 110498 503300 111551
rect 503260 110492 503312 110498
rect 503260 110434 503312 110440
rect 503350 108080 503406 108089
rect 503350 108015 503406 108024
rect 503364 107710 503392 108015
rect 503352 107704 503404 107710
rect 503352 107646 503404 107652
rect 502984 105528 503036 105534
rect 502984 105470 503036 105476
rect 502892 99340 502944 99346
rect 502892 99282 502944 99288
rect 502800 15972 502852 15978
rect 502800 15914 502852 15920
rect 502524 12436 502576 12442
rect 502524 12378 502576 12384
rect 502536 9654 502564 12378
rect 502524 9648 502576 9654
rect 502524 9590 502576 9596
rect 502432 4684 502484 4690
rect 502432 4626 502484 4632
rect 502996 3874 503024 105470
rect 503076 99340 503128 99346
rect 503076 99282 503128 99288
rect 503088 97646 503116 99282
rect 503076 97640 503128 97646
rect 503076 97582 503128 97588
rect 503732 14754 503760 147999
rect 503824 55894 503852 177375
rect 503916 107574 503944 371039
rect 503994 367296 504050 367305
rect 503994 367231 504050 367240
rect 504008 367130 504036 367231
rect 503996 367124 504048 367130
rect 503996 367066 504048 367072
rect 504468 367062 504496 393246
rect 504456 367056 504508 367062
rect 504456 366998 504508 367004
rect 504364 366988 504416 366994
rect 504364 366930 504416 366936
rect 503994 363760 504050 363769
rect 503994 363695 504050 363704
rect 504008 362982 504036 363695
rect 503996 362976 504048 362982
rect 503996 362918 504048 362924
rect 503994 359952 504050 359961
rect 503994 359887 504050 359896
rect 504008 151201 504036 359887
rect 504086 345536 504142 345545
rect 504086 345471 504142 345480
rect 504100 345098 504128 345471
rect 504088 345092 504140 345098
rect 504376 345080 504404 366930
rect 504376 345052 504496 345080
rect 504088 345034 504140 345040
rect 504086 341728 504142 341737
rect 504086 341663 504142 341672
rect 504100 340950 504128 341663
rect 504088 340944 504140 340950
rect 504088 340886 504140 340892
rect 504086 338192 504142 338201
rect 504086 338127 504088 338136
rect 504140 338127 504142 338136
rect 504088 338098 504140 338104
rect 504088 335300 504140 335306
rect 504088 335242 504140 335248
rect 504100 334393 504128 335242
rect 504086 334384 504142 334393
rect 504086 334319 504142 334328
rect 504468 325802 504496 345052
rect 504468 325774 504588 325802
rect 504560 325666 504588 325774
rect 504468 325638 504588 325666
rect 504086 323504 504142 323513
rect 504086 323439 504142 323448
rect 504100 322998 504128 323439
rect 504088 322992 504140 322998
rect 504088 322934 504140 322940
rect 504086 319968 504142 319977
rect 504086 319903 504142 319912
rect 504100 318850 504128 319903
rect 504088 318844 504140 318850
rect 504088 318786 504140 318792
rect 504086 316160 504142 316169
rect 504086 316095 504142 316104
rect 504100 316062 504128 316095
rect 504088 316056 504140 316062
rect 504088 315998 504140 316004
rect 504468 314702 504496 325638
rect 504364 314696 504416 314702
rect 504364 314638 504416 314644
rect 504456 314696 504508 314702
rect 504456 314638 504508 314644
rect 504376 307034 504404 314638
rect 504376 307006 504496 307034
rect 504088 306332 504140 306338
rect 504088 306274 504140 306280
rect 504100 305289 504128 306274
rect 504086 305280 504142 305289
rect 504086 305215 504142 305224
rect 504086 294400 504142 294409
rect 504086 294335 504142 294344
rect 504100 294030 504128 294335
rect 504088 294024 504140 294030
rect 504088 293966 504140 293972
rect 504468 293298 504496 307006
rect 504376 293270 504496 293298
rect 504086 290592 504142 290601
rect 504086 290527 504142 290536
rect 504100 289882 504128 290527
rect 504088 289876 504140 289882
rect 504088 289818 504140 289824
rect 504086 287056 504142 287065
rect 504086 286991 504142 287000
rect 504100 285734 504128 286991
rect 504088 285728 504140 285734
rect 504088 285670 504140 285676
rect 504178 283384 504234 283393
rect 504178 283319 504234 283328
rect 504086 283248 504142 283257
rect 504086 283183 504142 283192
rect 504100 282946 504128 283183
rect 504088 282940 504140 282946
rect 504088 282882 504140 282888
rect 504192 280401 504220 283319
rect 504178 280392 504234 280401
rect 504178 280327 504234 280336
rect 504086 275904 504142 275913
rect 504086 275839 504142 275848
rect 504100 274718 504128 275839
rect 504088 274712 504140 274718
rect 504088 274654 504140 274660
rect 504086 268832 504142 268841
rect 504086 268767 504142 268776
rect 504100 267782 504128 268767
rect 504088 267776 504140 267782
rect 504088 267718 504140 267724
rect 504086 261488 504142 261497
rect 504086 261423 504142 261432
rect 504100 260914 504128 261423
rect 504088 260908 504140 260914
rect 504088 260850 504140 260856
rect 504086 257680 504142 257689
rect 504086 257615 504142 257624
rect 504100 256766 504128 257615
rect 504088 256760 504140 256766
rect 504088 256702 504140 256708
rect 504086 250336 504142 250345
rect 504086 250271 504142 250280
rect 504100 249830 504128 250271
rect 504088 249824 504140 249830
rect 504088 249766 504140 249772
rect 504086 246800 504142 246809
rect 504086 246735 504142 246744
rect 504100 245682 504128 246735
rect 504088 245676 504140 245682
rect 504088 245618 504140 245624
rect 504086 243264 504142 243273
rect 504086 243199 504142 243208
rect 504100 242962 504128 243199
rect 504088 242956 504140 242962
rect 504088 242898 504140 242904
rect 504086 235920 504142 235929
rect 504086 235855 504142 235864
rect 504100 234666 504128 235855
rect 504088 234660 504140 234666
rect 504088 234602 504140 234608
rect 504086 232112 504142 232121
rect 504086 232047 504142 232056
rect 504100 231878 504128 232047
rect 504088 231872 504140 231878
rect 504088 231814 504140 231820
rect 504086 228576 504142 228585
rect 504086 228511 504142 228520
rect 504100 227798 504128 228511
rect 504088 227792 504140 227798
rect 504088 227734 504140 227740
rect 504086 224768 504142 224777
rect 504086 224703 504142 224712
rect 504100 223650 504128 224703
rect 504088 223644 504140 223650
rect 504088 223586 504140 223592
rect 504086 221232 504142 221241
rect 504086 221167 504142 221176
rect 504100 220930 504128 221167
rect 504088 220924 504140 220930
rect 504088 220866 504140 220872
rect 504086 213888 504142 213897
rect 504086 213823 504142 213832
rect 504100 212566 504128 213823
rect 504088 212560 504140 212566
rect 504088 212502 504140 212508
rect 504086 210352 504142 210361
rect 504086 210287 504142 210296
rect 504100 209846 504128 210287
rect 504088 209840 504140 209846
rect 504088 209782 504140 209788
rect 504086 203008 504142 203017
rect 504086 202943 504142 202952
rect 503994 151192 504050 151201
rect 503994 151127 504050 151136
rect 503994 118960 504050 118969
rect 503994 118895 504050 118904
rect 503904 107568 503956 107574
rect 503904 107510 503956 107516
rect 504008 98870 504036 118895
rect 503996 98864 504048 98870
rect 503996 98806 504048 98812
rect 504100 65550 504128 202943
rect 504178 195664 504234 195673
rect 504178 195599 504234 195608
rect 504192 194614 504220 195599
rect 504180 194608 504232 194614
rect 504180 194550 504232 194556
rect 504270 194440 504326 194449
rect 504270 194375 504326 194384
rect 504178 188320 504234 188329
rect 504178 188255 504234 188264
rect 504192 187746 504220 188255
rect 504180 187740 504232 187746
rect 504180 187682 504232 187688
rect 504284 186402 504312 194375
rect 504376 193866 504404 293270
rect 504364 193860 504416 193866
rect 504364 193802 504416 193808
rect 504192 186374 504312 186402
rect 504192 185201 504220 186374
rect 504270 186280 504326 186289
rect 504270 186215 504326 186224
rect 504284 185337 504312 186215
rect 504270 185328 504326 185337
rect 504270 185263 504326 185272
rect 504178 185192 504234 185201
rect 504178 185127 504234 185136
rect 504270 184784 504326 184793
rect 504270 184719 504326 184728
rect 504178 176624 504234 176633
rect 504178 176559 504234 176568
rect 504192 175409 504220 176559
rect 504178 175400 504234 175409
rect 504178 175335 504234 175344
rect 504178 173632 504234 173641
rect 504178 173567 504234 173576
rect 504192 68338 504220 173567
rect 504284 86358 504312 184719
rect 504362 175128 504418 175137
rect 504362 175063 504418 175072
rect 504376 165889 504404 175063
rect 504362 165880 504418 165889
rect 504362 165815 504418 165824
rect 504454 162752 504510 162761
rect 504454 162687 504510 162696
rect 504364 107568 504416 107574
rect 504364 107510 504416 107516
rect 504376 101590 504404 107510
rect 504468 105534 504496 162687
rect 504546 144528 504602 144537
rect 504546 144463 504602 144472
rect 504560 143614 504588 144463
rect 504548 143608 504600 143614
rect 504548 143550 504600 143556
rect 504546 140992 504602 141001
rect 504546 140927 504602 140936
rect 504560 140826 504588 140927
rect 504548 140820 504600 140826
rect 504548 140762 504600 140768
rect 504546 126304 504602 126313
rect 504546 126239 504602 126248
rect 504560 125662 504588 126239
rect 504548 125656 504600 125662
rect 504548 125598 504600 125604
rect 504456 105528 504508 105534
rect 504456 105470 504508 105476
rect 504546 104272 504602 104281
rect 504546 104207 504602 104216
rect 504560 103562 504588 104207
rect 504548 103556 504600 103562
rect 504548 103498 504600 103504
rect 504364 101584 504416 101590
rect 504364 101526 504416 101532
rect 505112 91866 505140 396607
rect 505190 392864 505246 392873
rect 505190 392799 505246 392808
rect 505204 93498 505232 392799
rect 505282 356416 505338 356425
rect 505282 356351 505338 356360
rect 505192 93492 505244 93498
rect 505192 93434 505244 93440
rect 505100 91860 505152 91866
rect 505100 91802 505152 91808
rect 504272 86352 504324 86358
rect 504272 86294 504324 86300
rect 504180 68332 504232 68338
rect 504180 68274 504232 68280
rect 505296 65618 505324 356351
rect 505756 355366 505784 607174
rect 508504 606144 508556 606150
rect 508504 606086 508556 606092
rect 507216 603152 507268 603158
rect 507216 603094 507268 603100
rect 507124 601724 507176 601730
rect 507124 601666 507176 601672
rect 506480 524476 506532 524482
rect 506480 524418 506532 524424
rect 505744 355360 505796 355366
rect 505744 355302 505796 355308
rect 505374 330848 505430 330857
rect 505374 330783 505430 330792
rect 505388 97510 505416 330783
rect 505466 301472 505522 301481
rect 505466 301407 505522 301416
rect 505376 97504 505428 97510
rect 505376 97446 505428 97452
rect 505480 80714 505508 301407
rect 505558 254144 505614 254153
rect 505558 254079 505614 254088
rect 505572 94654 505600 254079
rect 505650 180976 505706 180985
rect 505650 180911 505706 180920
rect 505664 101658 505692 180911
rect 505742 129840 505798 129849
rect 505742 129775 505798 129784
rect 505652 101652 505704 101658
rect 505652 101594 505704 101600
rect 505756 100094 505784 129775
rect 505744 100088 505796 100094
rect 505744 100030 505796 100036
rect 505560 94648 505612 94654
rect 505560 94590 505612 94596
rect 505468 80708 505520 80714
rect 505468 80650 505520 80656
rect 506492 79422 506520 524418
rect 506572 447160 506624 447166
rect 506572 447102 506624 447108
rect 506480 79416 506532 79422
rect 506480 79358 506532 79364
rect 505284 65612 505336 65618
rect 505284 65554 505336 65560
rect 504088 65544 504140 65550
rect 504088 65486 504140 65492
rect 504364 60036 504416 60042
rect 504364 59978 504416 59984
rect 503812 55888 503864 55894
rect 503812 55830 503864 55836
rect 503720 14748 503772 14754
rect 503720 14690 503772 14696
rect 503628 4684 503680 4690
rect 503628 4626 503680 4632
rect 502984 3868 503036 3874
rect 502984 3810 503036 3816
rect 500960 604 501012 610
rect 500960 546 501012 552
rect 501236 604 501288 610
rect 501236 546 501288 552
rect 502432 604 502484 610
rect 502432 546 502484 552
rect 501248 480 501276 546
rect 502444 480 502472 546
rect 503640 480 503668 4626
rect 504376 3058 504404 59978
rect 506584 58682 506612 447102
rect 506756 432540 506808 432546
rect 506756 432482 506808 432488
rect 506664 420980 506716 420986
rect 506664 420922 506716 420928
rect 506676 62830 506704 420922
rect 506768 87650 506796 432482
rect 507136 393310 507164 601666
rect 507228 534070 507256 603094
rect 507860 602268 507912 602274
rect 507860 602210 507912 602216
rect 507308 601384 507360 601390
rect 507308 601326 507360 601332
rect 507320 587178 507348 601326
rect 507308 587172 507360 587178
rect 507308 587114 507360 587120
rect 507216 534064 507268 534070
rect 507216 534006 507268 534012
rect 507124 393304 507176 393310
rect 507124 393246 507176 393252
rect 506940 378208 506992 378214
rect 506940 378150 506992 378156
rect 506848 367124 506900 367130
rect 506848 367066 506900 367072
rect 506756 87644 506808 87650
rect 506756 87586 506808 87592
rect 506664 62824 506716 62830
rect 506664 62766 506716 62772
rect 506572 58676 506624 58682
rect 506572 58618 506624 58624
rect 505100 55956 505152 55962
rect 505100 55898 505152 55904
rect 504822 3360 504878 3369
rect 504822 3295 504878 3304
rect 504364 3052 504416 3058
rect 504364 2994 504416 3000
rect 504836 480 504864 3295
rect 505112 610 505140 55898
rect 506860 29646 506888 367066
rect 506952 43518 506980 378150
rect 507124 260908 507176 260914
rect 507124 260850 507176 260856
rect 507032 242956 507084 242962
rect 507032 242898 507084 242904
rect 507044 49026 507072 242898
rect 507136 93770 507164 260850
rect 507124 93764 507176 93770
rect 507124 93706 507176 93712
rect 507032 49020 507084 49026
rect 507032 48962 507084 48968
rect 506940 43512 506992 43518
rect 506940 43454 506992 43460
rect 506848 29640 506900 29646
rect 506848 29582 506900 29588
rect 507872 3398 507900 602210
rect 508516 499526 508544 606086
rect 509332 600840 509384 600846
rect 509332 600782 509384 600788
rect 508504 499520 508556 499526
rect 508504 499462 508556 499468
rect 507952 498228 508004 498234
rect 507952 498170 508004 498176
rect 507964 91934 507992 498170
rect 508044 461576 508096 461582
rect 508044 461518 508096 461524
rect 507952 91928 508004 91934
rect 507952 91870 508004 91876
rect 508056 89010 508084 461518
rect 508228 407176 508280 407182
rect 508228 407118 508280 407124
rect 508136 256760 508188 256766
rect 508136 256702 508188 256708
rect 508044 89004 508096 89010
rect 508044 88946 508096 88952
rect 507860 3392 507912 3398
rect 507860 3334 507912 3340
rect 507216 3052 507268 3058
rect 507216 2994 507268 3000
rect 505100 604 505152 610
rect 505100 546 505152 552
rect 506020 604 506072 610
rect 506020 546 506072 552
rect 506032 480 506060 546
rect 507228 480 507256 2994
rect 508148 610 508176 256702
rect 508240 84862 508268 407118
rect 508320 289876 508372 289882
rect 508320 289818 508372 289824
rect 508228 84856 508280 84862
rect 508228 84798 508280 84804
rect 508332 66910 508360 289818
rect 509240 171828 509292 171834
rect 509240 171770 509292 171776
rect 509252 170814 509280 171770
rect 509240 170808 509292 170814
rect 509240 170750 509292 170756
rect 508412 140820 508464 140826
rect 508412 140762 508464 140768
rect 508424 96218 508452 140762
rect 508504 133068 508556 133074
rect 508504 133010 508556 133016
rect 508516 101930 508544 133010
rect 509240 110492 509292 110498
rect 509240 110434 509292 110440
rect 509252 102882 509280 110434
rect 509240 102876 509292 102882
rect 509240 102818 509292 102824
rect 508504 101924 508556 101930
rect 508504 101866 508556 101872
rect 509344 98977 509372 600782
rect 509884 600364 509936 600370
rect 509884 600306 509936 600312
rect 509896 452606 509924 600306
rect 509884 452600 509936 452606
rect 509884 452542 509936 452548
rect 509608 443012 509660 443018
rect 509608 442954 509660 442960
rect 509516 440292 509568 440298
rect 509516 440234 509568 440240
rect 509424 425128 509476 425134
rect 509424 425070 509476 425076
rect 509330 98968 509386 98977
rect 509330 98903 509386 98912
rect 508412 96212 508464 96218
rect 508412 96154 508464 96160
rect 509238 69592 509294 69601
rect 509238 69527 509294 69536
rect 508320 66904 508372 66910
rect 508320 66846 508372 66852
rect 509252 626 509280 69527
rect 509436 18630 509464 425070
rect 509528 61402 509556 440234
rect 509620 64190 509648 442954
rect 509700 220924 509752 220930
rect 509700 220866 509752 220872
rect 509712 98734 509740 220866
rect 509792 125656 509844 125662
rect 509792 125598 509844 125604
rect 509804 101794 509832 125598
rect 509792 101788 509844 101794
rect 509792 101730 509844 101736
rect 509988 100298 510016 700402
rect 515404 638988 515456 638994
rect 515404 638930 515456 638936
rect 514944 606348 514996 606354
rect 514944 606290 514996 606296
rect 513564 604988 513616 604994
rect 513564 604930 513616 604936
rect 513380 604920 513432 604926
rect 513380 604862 513432 604868
rect 512092 603288 512144 603294
rect 510710 603256 510766 603265
rect 512092 603230 512144 603236
rect 510710 603191 510766 603200
rect 510620 601860 510672 601866
rect 510620 601802 510672 601808
rect 509976 100292 510028 100298
rect 509976 100234 510028 100240
rect 509700 98728 509752 98734
rect 509700 98670 509752 98676
rect 509608 64184 509660 64190
rect 509608 64126 509660 64132
rect 509516 61396 509568 61402
rect 509516 61338 509568 61344
rect 509424 18624 509476 18630
rect 509424 18566 509476 18572
rect 510632 6662 510660 601802
rect 510724 96082 510752 603191
rect 511356 600772 511408 600778
rect 511356 600714 511408 600720
rect 511264 592068 511316 592074
rect 511264 592010 511316 592016
rect 510804 469260 510856 469266
rect 510804 469202 510856 469208
rect 510816 99006 510844 469202
rect 510896 227792 510948 227798
rect 510896 227734 510948 227740
rect 510908 102134 510936 227734
rect 510988 143608 511040 143614
rect 510988 143550 511040 143556
rect 510896 102128 510948 102134
rect 510896 102070 510948 102076
rect 510804 99000 510856 99006
rect 510804 98942 510856 98948
rect 511000 96286 511028 143550
rect 511276 100502 511304 592010
rect 511368 171086 511396 600714
rect 511448 204332 511500 204338
rect 511448 204274 511500 204280
rect 511356 171080 511408 171086
rect 511356 171022 511408 171028
rect 511356 103556 511408 103562
rect 511356 103498 511408 103504
rect 511264 100496 511316 100502
rect 511264 100438 511316 100444
rect 510988 96280 511040 96286
rect 510988 96222 511040 96228
rect 510712 96076 510764 96082
rect 510712 96018 510764 96024
rect 511368 11898 511396 103498
rect 511460 100842 511488 204274
rect 511448 100836 511500 100842
rect 511448 100778 511500 100784
rect 511446 87544 511502 87553
rect 511446 87479 511502 87488
rect 511356 11892 511408 11898
rect 511356 11834 511408 11840
rect 510804 9240 510856 9246
rect 510804 9182 510856 9188
rect 510620 6656 510672 6662
rect 510620 6598 510672 6604
rect 508136 604 508188 610
rect 508136 546 508188 552
rect 508412 604 508464 610
rect 509252 598 509648 626
rect 508412 546 508464 552
rect 508424 480 508452 546
rect 509620 480 509648 598
rect 510816 480 510844 9182
rect 511460 4146 511488 87479
rect 512104 9042 512132 603230
rect 512828 596828 512880 596834
rect 512828 596770 512880 596776
rect 512840 570217 512868 596770
rect 512826 570208 512882 570217
rect 512826 570143 512882 570152
rect 512826 570072 512882 570081
rect 512826 570007 512882 570016
rect 512840 568585 512868 570007
rect 512826 568576 512882 568585
rect 512826 568511 512882 568520
rect 513010 568576 513066 568585
rect 513010 568511 513066 568520
rect 513024 558958 513052 568511
rect 512828 558952 512880 558958
rect 512828 558894 512880 558900
rect 513012 558952 513064 558958
rect 513012 558894 513064 558900
rect 512840 549273 512868 558894
rect 512826 549264 512882 549273
rect 512826 549199 512882 549208
rect 513010 549264 513066 549273
rect 513010 549199 513066 549208
rect 512644 545148 512696 545154
rect 512644 545090 512696 545096
rect 512184 322992 512236 322998
rect 512184 322934 512236 322940
rect 512092 9036 512144 9042
rect 512092 8978 512144 8984
rect 511448 4140 511500 4146
rect 511448 4082 511500 4088
rect 512196 4078 512224 322934
rect 512276 294024 512328 294030
rect 512276 293966 512328 293972
rect 512288 99142 512316 293966
rect 512460 223644 512512 223650
rect 512460 223586 512512 223592
rect 512368 165640 512420 165646
rect 512368 165582 512420 165588
rect 512276 99136 512328 99142
rect 512276 99078 512328 99084
rect 512184 4072 512236 4078
rect 512184 4014 512236 4020
rect 512380 3806 512408 165582
rect 512472 101522 512500 223586
rect 512552 209840 512604 209846
rect 512552 209782 512604 209788
rect 512460 101516 512512 101522
rect 512460 101458 512512 101464
rect 512564 98938 512592 209782
rect 512552 98932 512604 98938
rect 512552 98874 512604 98880
rect 512656 96490 512684 545090
rect 513024 531350 513052 549199
rect 512828 531344 512880 531350
rect 512828 531286 512880 531292
rect 513012 531344 513064 531350
rect 513012 531286 513064 531292
rect 512840 529922 512868 531286
rect 512828 529916 512880 529922
rect 512828 529858 512880 529864
rect 513012 529916 513064 529922
rect 513012 529858 513064 529864
rect 513024 512038 513052 529858
rect 512828 512032 512880 512038
rect 512828 511974 512880 511980
rect 513012 512032 513064 512038
rect 513012 511974 513064 511980
rect 512840 510610 512868 511974
rect 512828 510604 512880 510610
rect 512828 510546 512880 510552
rect 513012 510604 513064 510610
rect 513012 510546 513064 510552
rect 513024 500993 513052 510546
rect 512826 500984 512882 500993
rect 512826 500919 512882 500928
rect 513010 500984 513066 500993
rect 513010 500919 513066 500928
rect 512840 491298 512868 500919
rect 512828 491292 512880 491298
rect 512828 491234 512880 491240
rect 512828 481704 512880 481710
rect 512828 481646 512880 481652
rect 512840 471986 512868 481646
rect 512828 471980 512880 471986
rect 512828 471922 512880 471928
rect 512828 462392 512880 462398
rect 512828 462334 512880 462340
rect 512840 452538 512868 462334
rect 512828 452532 512880 452538
rect 512828 452474 512880 452480
rect 512828 443012 512880 443018
rect 512828 442954 512880 442960
rect 512840 433294 512868 442954
rect 512828 433288 512880 433294
rect 512828 433230 512880 433236
rect 512828 423700 512880 423706
rect 512828 423642 512880 423648
rect 512840 413982 512868 423642
rect 512828 413976 512880 413982
rect 512828 413918 512880 413924
rect 512828 404388 512880 404394
rect 512828 404330 512880 404336
rect 512840 394670 512868 404330
rect 512828 394664 512880 394670
rect 512828 394606 512880 394612
rect 512828 385144 512880 385150
rect 512828 385086 512880 385092
rect 512840 377074 512868 385086
rect 512840 377046 512960 377074
rect 512932 376802 512960 377046
rect 512840 376774 512960 376802
rect 512840 375290 512868 376774
rect 512828 375284 512880 375290
rect 512828 375226 512880 375232
rect 512828 365764 512880 365770
rect 512828 365706 512880 365712
rect 512840 357610 512868 365706
rect 512828 357604 512880 357610
rect 512828 357546 512880 357552
rect 512828 357468 512880 357474
rect 512828 357410 512880 357416
rect 512840 356046 512868 357410
rect 512828 356040 512880 356046
rect 512828 355982 512880 355988
rect 512828 346452 512880 346458
rect 512828 346394 512880 346400
rect 512840 336734 512868 346394
rect 512828 336728 512880 336734
rect 512828 336670 512880 336676
rect 512828 327140 512880 327146
rect 512828 327082 512880 327088
rect 512840 317422 512868 327082
rect 512828 317416 512880 317422
rect 512828 317358 512880 317364
rect 512920 317416 512972 317422
rect 512920 317358 512972 317364
rect 512932 299554 512960 317358
rect 512840 299526 512960 299554
rect 512840 298110 512868 299526
rect 512828 298104 512880 298110
rect 512828 298046 512880 298052
rect 512920 298104 512972 298110
rect 512920 298046 512972 298052
rect 512932 280242 512960 298046
rect 512840 280214 512960 280242
rect 512840 278769 512868 280214
rect 512826 278760 512882 278769
rect 512826 278695 512882 278704
rect 513010 278760 513066 278769
rect 513010 278695 513066 278704
rect 513024 269142 513052 278695
rect 512828 269136 512880 269142
rect 512828 269078 512880 269084
rect 513012 269136 513064 269142
rect 513012 269078 513064 269084
rect 512840 261066 512868 269078
rect 512840 261038 512960 261066
rect 512932 260930 512960 261038
rect 512840 260902 512960 260930
rect 512840 259457 512868 260902
rect 512826 259448 512882 259457
rect 512826 259383 512882 259392
rect 513010 259448 513066 259457
rect 513010 259383 513066 259392
rect 513024 249898 513052 259383
rect 512828 249892 512880 249898
rect 512828 249834 512880 249840
rect 513012 249892 513064 249898
rect 513012 249834 513064 249840
rect 512840 240145 512868 249834
rect 512826 240136 512882 240145
rect 512826 240071 512882 240080
rect 513010 240136 513066 240145
rect 513010 240071 513066 240080
rect 513024 230518 513052 240071
rect 512828 230512 512880 230518
rect 512828 230454 512880 230460
rect 513012 230512 513064 230518
rect 513012 230454 513064 230460
rect 512840 220833 512868 230454
rect 512826 220824 512882 220833
rect 512826 220759 512882 220768
rect 513010 220824 513066 220833
rect 513010 220759 513066 220768
rect 513024 211177 513052 220759
rect 512826 211168 512882 211177
rect 512826 211103 512882 211112
rect 513010 211168 513066 211177
rect 513010 211103 513066 211112
rect 512840 201482 512868 211103
rect 512828 201476 512880 201482
rect 512828 201418 512880 201424
rect 513012 201476 513064 201482
rect 513012 201418 513064 201424
rect 513024 191865 513052 201418
rect 512826 191856 512882 191865
rect 512826 191791 512882 191800
rect 513010 191856 513066 191865
rect 513010 191791 513066 191800
rect 512840 182170 512868 191791
rect 512828 182164 512880 182170
rect 512828 182106 512880 182112
rect 513012 182164 513064 182170
rect 513012 182106 513064 182112
rect 513024 172553 513052 182106
rect 512826 172544 512882 172553
rect 512826 172479 512882 172488
rect 513010 172544 513066 172553
rect 513010 172479 513066 172488
rect 512840 162858 512868 172479
rect 512828 162852 512880 162858
rect 512828 162794 512880 162800
rect 512828 153264 512880 153270
rect 512828 153206 512880 153212
rect 512840 143546 512868 153206
rect 512828 143540 512880 143546
rect 512828 143482 512880 143488
rect 512828 133952 512880 133958
rect 512828 133894 512880 133900
rect 512840 124166 512868 133894
rect 512828 124160 512880 124166
rect 512828 124102 512880 124108
rect 512828 114572 512880 114578
rect 512828 114514 512880 114520
rect 512840 104854 512868 114514
rect 512828 104848 512880 104854
rect 512828 104790 512880 104796
rect 513288 100768 513340 100774
rect 513288 100710 513340 100716
rect 513300 99346 513328 100710
rect 513288 99340 513340 99346
rect 513288 99282 513340 99288
rect 512644 96484 512696 96490
rect 512644 96426 512696 96432
rect 512736 95260 512788 95266
rect 512736 95202 512788 95208
rect 512748 87038 512776 95202
rect 512736 87032 512788 87038
rect 512736 86974 512788 86980
rect 512828 87032 512880 87038
rect 512828 86974 512880 86980
rect 512840 85542 512868 86974
rect 512828 85536 512880 85542
rect 512828 85478 512880 85484
rect 512828 75948 512880 75954
rect 512828 75890 512880 75896
rect 512840 66230 512868 75890
rect 512828 66224 512880 66230
rect 512828 66166 512880 66172
rect 512828 56636 512880 56642
rect 512828 56578 512880 56584
rect 512840 46918 512868 56578
rect 512828 46912 512880 46918
rect 512828 46854 512880 46860
rect 512828 37324 512880 37330
rect 512828 37266 512880 37272
rect 512840 27606 512868 37266
rect 512828 27600 512880 27606
rect 512828 27542 512880 27548
rect 512460 9716 512512 9722
rect 512460 9658 512512 9664
rect 512472 9602 512500 9658
rect 512472 9574 512592 9602
rect 512368 3800 512420 3806
rect 512368 3742 512420 3748
rect 512564 2786 512592 9574
rect 513196 4140 513248 4146
rect 513196 4082 513248 4088
rect 512000 2780 512052 2786
rect 512000 2722 512052 2728
rect 512552 2780 512604 2786
rect 512552 2722 512604 2728
rect 512012 480 512040 2722
rect 513208 480 513236 4082
rect 513392 3738 513420 604862
rect 513472 603764 513524 603770
rect 513472 603706 513524 603712
rect 513484 3942 513512 603706
rect 513576 6526 513604 604930
rect 514116 604580 514168 604586
rect 514116 604522 514168 604528
rect 514024 599684 514076 599690
rect 514024 599626 514076 599632
rect 513656 494080 513708 494086
rect 513656 494022 513708 494028
rect 513564 6520 513616 6526
rect 513564 6462 513616 6468
rect 513472 3936 513524 3942
rect 513472 3878 513524 3884
rect 513380 3732 513432 3738
rect 513380 3674 513432 3680
rect 513668 610 513696 494022
rect 513748 403028 513800 403034
rect 513748 402970 513800 402976
rect 513760 8294 513788 402970
rect 513840 345092 513892 345098
rect 513840 345034 513892 345040
rect 513852 101998 513880 345034
rect 514036 322930 514064 599626
rect 514128 440230 514156 604522
rect 514760 601928 514812 601934
rect 514760 601870 514812 601876
rect 514116 440224 514168 440230
rect 514116 440166 514168 440172
rect 514116 368552 514168 368558
rect 514116 368494 514168 368500
rect 514024 322924 514076 322930
rect 514024 322866 514076 322872
rect 513932 194608 513984 194614
rect 513932 194550 513984 194556
rect 513840 101992 513892 101998
rect 513840 101934 513892 101940
rect 513944 101726 513972 194550
rect 513932 101720 513984 101726
rect 513932 101662 513984 101668
rect 514128 100706 514156 368494
rect 514116 100700 514168 100706
rect 514116 100642 514168 100648
rect 513748 8288 513800 8294
rect 513748 8230 513800 8236
rect 514772 6594 514800 601870
rect 514852 564460 514904 564466
rect 514852 564402 514904 564408
rect 514864 22098 514892 564402
rect 514956 95849 514984 606290
rect 515036 545216 515088 545222
rect 515036 545158 515088 545164
rect 515048 96150 515076 545158
rect 515128 318844 515180 318850
rect 515128 318786 515180 318792
rect 515140 98802 515168 318786
rect 515312 267776 515364 267782
rect 515312 267718 515364 267724
rect 515220 193860 515272 193866
rect 515220 193802 515272 193808
rect 515128 98796 515180 98802
rect 515128 98738 515180 98744
rect 515036 96144 515088 96150
rect 515036 96086 515088 96092
rect 514942 95840 514998 95849
rect 514942 95775 514998 95784
rect 514852 22092 514904 22098
rect 514852 22034 514904 22040
rect 515232 6730 515260 193802
rect 515324 93294 515352 267718
rect 515416 100366 515444 638930
rect 520372 608660 520424 608666
rect 520372 608602 520424 608608
rect 517796 606076 517848 606082
rect 517796 606018 517848 606024
rect 516416 604852 516468 604858
rect 516416 604794 516468 604800
rect 515496 603560 515548 603566
rect 515496 603502 515548 603508
rect 516138 603528 516194 603537
rect 515508 311846 515536 603502
rect 516138 603463 516194 603472
rect 515496 311840 515548 311846
rect 515496 311782 515548 311788
rect 515404 100360 515456 100366
rect 515404 100302 515456 100308
rect 515312 93288 515364 93294
rect 515312 93230 515364 93236
rect 515220 6724 515272 6730
rect 515220 6666 515272 6672
rect 514760 6588 514812 6594
rect 514760 6530 514812 6536
rect 514666 5808 514722 5817
rect 514850 5808 514906 5817
rect 514722 5766 514850 5794
rect 514666 5743 514722 5752
rect 514850 5743 514906 5752
rect 516152 3777 516180 603463
rect 516324 603356 516376 603362
rect 516324 603298 516376 603304
rect 516232 600704 516284 600710
rect 516232 600646 516284 600652
rect 516244 6458 516272 600646
rect 516336 96422 516364 603298
rect 516428 97306 516456 604794
rect 516874 603936 516930 603945
rect 516874 603871 516930 603880
rect 516888 603770 516916 603871
rect 516876 603764 516928 603770
rect 516876 603706 516928 603712
rect 517612 603492 517664 603498
rect 517612 603434 517664 603440
rect 517518 601896 517574 601905
rect 517518 601831 517574 601840
rect 516508 476128 516560 476134
rect 516508 476070 516560 476076
rect 516416 97300 516468 97306
rect 516416 97242 516468 97248
rect 516324 96416 516376 96422
rect 516324 96358 516376 96364
rect 516520 96014 516548 476070
rect 516784 404388 516836 404394
rect 516784 404330 516836 404336
rect 516600 362976 516652 362982
rect 516600 362918 516652 362924
rect 516612 101561 516640 362918
rect 516692 234660 516744 234666
rect 516692 234602 516744 234608
rect 516598 101552 516654 101561
rect 516598 101487 516654 101496
rect 516508 96008 516560 96014
rect 516508 95950 516560 95956
rect 516704 93566 516732 234602
rect 516796 100638 516824 404330
rect 516784 100632 516836 100638
rect 516784 100574 516836 100580
rect 516692 93560 516744 93566
rect 516692 93502 516744 93508
rect 516324 11824 516376 11830
rect 516324 11766 516376 11772
rect 516232 6452 516284 6458
rect 516232 6394 516284 6400
rect 516138 3768 516194 3777
rect 516138 3703 516194 3712
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 513656 604 513708 610
rect 513656 546 513708 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 3470
rect 516336 3074 516364 11766
rect 517532 3482 517560 601831
rect 517624 3602 517652 603434
rect 517704 602472 517756 602478
rect 517704 602414 517756 602420
rect 517716 4010 517744 602414
rect 517808 97442 517836 606018
rect 517886 603392 517942 603401
rect 517886 603327 517942 603336
rect 517900 101697 517928 603327
rect 520278 602032 520334 602041
rect 520278 601967 520334 601976
rect 518164 600568 518216 600574
rect 518164 600510 518216 600516
rect 517980 567248 518032 567254
rect 517980 567190 518032 567196
rect 517886 101688 517942 101697
rect 517886 101623 517942 101632
rect 517992 98705 518020 567190
rect 518072 249824 518124 249830
rect 518072 249766 518124 249772
rect 517978 98696 518034 98705
rect 517978 98631 518034 98640
rect 517796 97436 517848 97442
rect 517796 97378 517848 97384
rect 518084 93226 518112 249766
rect 518072 93220 518124 93226
rect 518072 93162 518124 93168
rect 517704 4004 517756 4010
rect 517704 3946 517756 3952
rect 517612 3596 517664 3602
rect 517612 3538 517664 3544
rect 518176 3534 518204 600510
rect 518900 600432 518952 600438
rect 518900 600374 518952 600380
rect 518912 9110 518940 600374
rect 518992 549296 519044 549302
rect 518992 549238 519044 549244
rect 519004 99210 519032 549238
rect 519084 436144 519136 436150
rect 519084 436086 519136 436092
rect 518992 99204 519044 99210
rect 518992 99146 519044 99152
rect 519096 98666 519124 436086
rect 519176 380928 519228 380934
rect 519176 380870 519228 380876
rect 519188 101454 519216 380870
rect 519636 355360 519688 355366
rect 519636 355302 519688 355308
rect 519268 338156 519320 338162
rect 519268 338098 519320 338104
rect 519176 101448 519228 101454
rect 519176 101390 519228 101396
rect 519084 98660 519136 98666
rect 519084 98602 519136 98608
rect 519280 96354 519308 338098
rect 519360 274712 519412 274718
rect 519360 274654 519412 274660
rect 519268 96348 519320 96354
rect 519268 96290 519320 96296
rect 519372 90438 519400 274654
rect 519544 231872 519596 231878
rect 519544 231814 519596 231820
rect 519360 90432 519412 90438
rect 519360 90374 519412 90380
rect 519556 64870 519584 231814
rect 519648 231470 519676 355302
rect 519636 231464 519688 231470
rect 519636 231406 519688 231412
rect 519544 64864 519596 64870
rect 519544 64806 519596 64812
rect 518992 17264 519044 17270
rect 518992 17206 519044 17212
rect 518900 9104 518952 9110
rect 518900 9046 518952 9052
rect 518164 3528 518216 3534
rect 517532 3454 517928 3482
rect 518164 3470 518216 3476
rect 516336 3046 516732 3074
rect 516704 626 516732 3046
rect 516704 598 516824 626
rect 516796 480 516824 598
rect 517900 480 517928 3454
rect 519004 1578 519032 17206
rect 520292 3602 520320 601967
rect 520384 3670 520412 608602
rect 520476 100434 520504 700470
rect 522304 685908 522356 685914
rect 522304 685850 522356 685856
rect 521844 608728 521896 608734
rect 521844 608670 521896 608676
rect 521660 607368 521712 607374
rect 521660 607310 521712 607316
rect 520556 606280 520608 606286
rect 520556 606222 520608 606228
rect 520464 100428 520516 100434
rect 520464 100370 520516 100376
rect 520568 97374 520596 606222
rect 520648 560312 520700 560318
rect 520648 560254 520700 560260
rect 520660 99074 520688 560254
rect 520740 520328 520792 520334
rect 520740 520270 520792 520276
rect 520648 99068 520700 99074
rect 520648 99010 520700 99016
rect 520556 97368 520608 97374
rect 520556 97310 520608 97316
rect 520752 93362 520780 520270
rect 520832 398880 520884 398886
rect 520832 398822 520884 398828
rect 520844 95946 520872 398822
rect 520924 231464 520976 231470
rect 520924 231406 520976 231412
rect 520936 100774 520964 231406
rect 521566 200016 521622 200025
rect 521566 199951 521622 199960
rect 521580 190505 521608 199951
rect 521566 190496 521622 190505
rect 521566 190431 521622 190440
rect 520924 100768 520976 100774
rect 520924 100710 520976 100716
rect 520832 95940 520884 95946
rect 520832 95882 520884 95888
rect 520740 93356 520792 93362
rect 520740 93298 520792 93304
rect 520464 39364 520516 39370
rect 520464 39306 520516 39312
rect 520372 3664 520424 3670
rect 520372 3606 520424 3612
rect 520280 3596 520332 3602
rect 520280 3538 520332 3544
rect 520476 3482 520504 39306
rect 521672 8974 521700 607310
rect 521752 605056 521804 605062
rect 521752 604998 521804 605004
rect 521764 93634 521792 604998
rect 521856 100026 521884 608670
rect 521934 579592 521990 579601
rect 521934 579527 521990 579536
rect 521948 570217 521976 579527
rect 521934 570208 521990 570217
rect 521934 570143 521990 570152
rect 522118 560280 522174 560289
rect 522118 560215 522174 560224
rect 522132 550769 522160 560215
rect 522118 550760 522174 550769
rect 522118 550695 522174 550704
rect 522026 540968 522082 540977
rect 522026 540903 522082 540912
rect 521936 538280 521988 538286
rect 521936 538222 521988 538228
rect 521844 100020 521896 100026
rect 521844 99962 521896 99968
rect 521752 93628 521804 93634
rect 521752 93570 521804 93576
rect 521948 93430 521976 538222
rect 522040 531593 522068 540903
rect 522026 531584 522082 531593
rect 522026 531519 522082 531528
rect 522026 521656 522082 521665
rect 522026 521591 522082 521600
rect 522040 512281 522068 521591
rect 522026 512272 522082 512281
rect 522026 512207 522082 512216
rect 522026 502344 522082 502353
rect 522026 502279 522082 502288
rect 522040 492697 522068 502279
rect 522026 492688 522082 492697
rect 522026 492623 522082 492632
rect 522028 483064 522080 483070
rect 522028 483006 522080 483012
rect 521936 93424 521988 93430
rect 521936 93366 521988 93372
rect 522040 93158 522068 483006
rect 522118 463448 522174 463457
rect 522118 463383 522174 463392
rect 522132 454073 522160 463383
rect 522118 454064 522174 454073
rect 522118 453999 522174 454008
rect 522120 429208 522172 429214
rect 522120 429150 522172 429156
rect 522132 93702 522160 429150
rect 522210 424960 522266 424969
rect 522210 424895 522266 424904
rect 522224 415449 522252 424895
rect 522210 415440 522266 415449
rect 522210 415375 522266 415384
rect 522210 405512 522266 405521
rect 522210 405447 522266 405456
rect 522224 396137 522252 405447
rect 522210 396128 522266 396137
rect 522210 396063 522266 396072
rect 522210 386200 522266 386209
rect 522210 386135 522266 386144
rect 522224 376825 522252 386135
rect 522210 376816 522266 376825
rect 522210 376751 522266 376760
rect 522316 375358 522344 685850
rect 523040 605940 523092 605946
rect 523040 605882 523092 605888
rect 522304 375352 522356 375358
rect 522304 375294 522356 375300
rect 522210 357368 522266 357377
rect 522210 357303 522266 357312
rect 522224 350577 522252 357303
rect 522210 350568 522266 350577
rect 522210 350503 522266 350512
rect 522210 347576 522266 347585
rect 522210 347511 522266 347520
rect 522224 338201 522252 347511
rect 522210 338192 522266 338201
rect 522210 338127 522266 338136
rect 522210 328400 522266 328409
rect 522210 328335 522266 328344
rect 522224 319025 522252 328335
rect 522210 319016 522266 319025
rect 522210 318951 522266 318960
rect 522210 308952 522266 308961
rect 522210 308887 522266 308896
rect 522224 302161 522252 308887
rect 522210 302152 522266 302161
rect 522210 302087 522266 302096
rect 522210 289640 522266 289649
rect 522210 289575 522266 289584
rect 522224 280401 522252 289575
rect 522210 280392 522266 280401
rect 522210 280327 522266 280336
rect 522210 270464 522266 270473
rect 522210 270399 522266 270408
rect 522224 261089 522252 270399
rect 522210 261080 522266 261089
rect 522210 261015 522266 261024
rect 522210 251152 522266 251161
rect 522210 251087 522266 251096
rect 522224 241777 522252 251087
rect 522210 241768 522266 241777
rect 522210 241703 522266 241712
rect 522210 222184 522266 222193
rect 522210 222119 522266 222128
rect 522224 212673 522252 222119
rect 522210 212664 522266 212673
rect 522210 212599 522266 212608
rect 522210 212528 522266 212537
rect 522210 212463 522266 212472
rect 522224 206281 522252 212463
rect 522210 206272 522266 206281
rect 522210 206207 522266 206216
rect 522210 173904 522266 173913
rect 522210 173839 522266 173848
rect 522224 164257 522252 173839
rect 522210 164248 522266 164257
rect 522210 164183 522266 164192
rect 522302 135144 522358 135153
rect 522302 135079 522358 135088
rect 522316 125633 522344 135079
rect 522302 125624 522358 125633
rect 522302 125559 522358 125568
rect 522210 115832 522266 115841
rect 522210 115767 522266 115776
rect 522224 106321 522252 115767
rect 522210 106312 522266 106321
rect 522210 106247 522266 106256
rect 522120 93696 522172 93702
rect 522120 93638 522172 93644
rect 522028 93152 522080 93158
rect 522028 93094 522080 93100
rect 521660 8968 521712 8974
rect 521660 8910 521712 8916
rect 521476 3596 521528 3602
rect 521476 3538 521528 3544
rect 520292 3454 520504 3482
rect 519004 1550 519124 1578
rect 519096 480 519124 1550
rect 520292 480 520320 3454
rect 521488 480 521516 3538
rect 522672 3460 522724 3466
rect 522672 3402 522724 3408
rect 522684 480 522712 3402
rect 523052 3346 523080 605882
rect 525708 603764 525760 603770
rect 525708 603706 525760 603712
rect 525720 603673 525748 603706
rect 525706 603664 525762 603673
rect 525706 603599 525762 603608
rect 524420 602200 524472 602206
rect 524420 602142 524472 602148
rect 523132 598324 523184 598330
rect 523132 598266 523184 598272
rect 523144 94722 523172 598266
rect 523224 587172 523276 587178
rect 523224 587114 523276 587120
rect 523236 97578 523264 587114
rect 523316 473408 523368 473414
rect 523316 473350 523368 473356
rect 523328 99278 523356 473350
rect 523408 382968 523460 382974
rect 523408 382910 523460 382916
rect 523420 102814 523448 382910
rect 523408 102808 523460 102814
rect 523408 102750 523460 102756
rect 523316 99272 523368 99278
rect 523316 99214 523368 99220
rect 523224 97572 523276 97578
rect 523224 97514 523276 97520
rect 523132 94716 523184 94722
rect 523132 94658 523184 94664
rect 524432 3346 524460 602142
rect 527192 171834 527220 703520
rect 543476 700330 543504 703520
rect 559668 700330 559696 703520
rect 529204 700324 529256 700330
rect 529204 700266 529256 700272
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 543556 700324 543608 700330
rect 543556 700266 543608 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 529216 554742 529244 700266
rect 543568 699718 543596 700266
rect 543004 699712 543056 699718
rect 543004 699654 543056 699660
rect 543556 699712 543608 699718
rect 543556 699654 543608 699660
rect 543016 610638 543044 699654
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 543004 610632 543056 610638
rect 543004 610574 543056 610580
rect 554044 606212 554096 606218
rect 554044 606154 554096 606160
rect 540886 603800 540942 603809
rect 540886 603735 540942 603744
rect 540900 603702 540928 603735
rect 533988 603696 534040 603702
rect 533986 603664 533988 603673
rect 540888 603696 540940 603702
rect 534040 603664 534042 603673
rect 540888 603638 540940 603644
rect 533986 603599 534042 603608
rect 531964 603424 532016 603430
rect 531964 603366 532016 603372
rect 529204 554736 529256 554742
rect 529204 554678 529256 554684
rect 527824 340944 527876 340950
rect 527824 340886 527876 340892
rect 527180 171828 527232 171834
rect 527180 171770 527232 171776
rect 527180 57316 527232 57322
rect 527180 57258 527232 57264
rect 525800 15904 525852 15910
rect 525800 15846 525852 15852
rect 525812 3346 525840 15846
rect 526442 5808 526498 5817
rect 526442 5743 526498 5752
rect 526456 5545 526484 5743
rect 526442 5536 526498 5545
rect 526442 5471 526498 5480
rect 527192 3346 527220 57258
rect 527836 4826 527864 340886
rect 531976 229090 532004 603366
rect 552664 603220 552716 603226
rect 552664 603162 552716 603168
rect 543004 601996 543056 602002
rect 543004 601938 543056 601944
rect 532700 600500 532752 600506
rect 532700 600442 532752 600448
rect 531964 229084 532016 229090
rect 531964 229026 532016 229032
rect 531964 107704 532016 107710
rect 531964 107646 532016 107652
rect 528560 86284 528612 86290
rect 528560 86226 528612 86232
rect 527824 4820 527876 4826
rect 527824 4762 527876 4768
rect 528572 3466 528600 86226
rect 531320 20120 531372 20126
rect 531320 20062 531372 20068
rect 528652 14884 528704 14890
rect 528652 14826 528704 14832
rect 528560 3460 528612 3466
rect 528560 3402 528612 3408
rect 523052 3318 523908 3346
rect 524432 3318 525104 3346
rect 525812 3318 526300 3346
rect 527192 3318 527496 3346
rect 523880 480 523908 3318
rect 525076 480 525104 3318
rect 526272 480 526300 3318
rect 527468 480 527496 3318
rect 528664 480 528692 14826
rect 529940 11756 529992 11762
rect 529940 11698 529992 11704
rect 529952 3482 529980 11698
rect 531332 3618 531360 20062
rect 531976 6458 532004 107646
rect 531964 6452 532016 6458
rect 531964 6394 532016 6400
rect 531332 3590 532280 3618
rect 529848 3460 529900 3466
rect 529952 3454 531084 3482
rect 529848 3402 529900 3408
rect 529860 480 529888 3402
rect 531056 480 531084 3454
rect 532252 480 532280 3590
rect 532712 3482 532740 600442
rect 534080 598256 534132 598262
rect 534080 598198 534132 598204
rect 534092 3482 534120 598198
rect 540244 586560 540296 586566
rect 540244 586502 540296 586508
rect 538864 571396 538916 571402
rect 538864 571338 538916 571344
rect 536840 547188 536892 547194
rect 536840 547130 536892 547136
rect 535734 4040 535790 4049
rect 535734 3975 535790 3984
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3975
rect 536852 2378 536880 547130
rect 538876 124166 538904 571338
rect 540256 299470 540284 586502
rect 540244 299464 540296 299470
rect 540244 299406 540296 299412
rect 540244 285728 540296 285734
rect 540244 285670 540296 285676
rect 540256 218006 540284 285670
rect 540244 218000 540296 218006
rect 540244 217942 540296 217948
rect 540244 212560 540296 212566
rect 540244 212502 540296 212508
rect 538864 124160 538916 124166
rect 538864 124102 538916 124108
rect 538220 43444 538272 43450
rect 538220 43386 538272 43392
rect 536930 6216 536986 6225
rect 536930 6151 536986 6160
rect 536840 2372 536892 2378
rect 536840 2314 536892 2320
rect 536944 480 536972 6151
rect 538232 3482 538260 43386
rect 539600 26920 539652 26926
rect 539600 26862 539652 26868
rect 539612 3482 539640 26862
rect 540256 8974 540284 212502
rect 540886 181384 540942 181393
rect 540886 181319 540942 181328
rect 540900 181121 540928 181319
rect 540886 181112 540942 181121
rect 540886 181047 540942 181056
rect 540980 49156 541032 49162
rect 540980 49098 541032 49104
rect 540244 8968 540296 8974
rect 540244 8910 540296 8916
rect 540992 3482 541020 49098
rect 542912 3528 542964 3534
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542912 3470 542964 3476
rect 538128 2372 538180 2378
rect 538128 2314 538180 2320
rect 538140 480 538168 2314
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3470
rect 543016 3330 543044 601938
rect 543740 600976 543792 600982
rect 543740 600918 543792 600924
rect 543752 3482 543780 600918
rect 549904 385076 549956 385082
rect 549904 385018 549956 385024
rect 545120 282940 545172 282946
rect 545120 282882 545172 282888
rect 545132 3482 545160 282882
rect 547144 245676 547196 245682
rect 547144 245618 547196 245624
rect 546592 18760 546644 18766
rect 546592 18702 546644 18708
rect 546604 3482 546632 18702
rect 547156 18018 547184 245618
rect 549916 41410 549944 385018
rect 552676 135250 552704 603162
rect 554056 276010 554084 606154
rect 573364 606008 573416 606014
rect 573364 605950 573416 605956
rect 554780 604648 554832 604654
rect 554780 604590 554832 604596
rect 558918 604616 558974 604625
rect 554044 276004 554096 276010
rect 554044 275946 554096 275952
rect 554044 187740 554096 187746
rect 554044 187682 554096 187688
rect 552756 151836 552808 151842
rect 552756 151778 552808 151784
rect 552664 135244 552716 135250
rect 552664 135186 552716 135192
rect 549904 41404 549956 41410
rect 549904 41346 549956 41352
rect 550640 25560 550692 25566
rect 550640 25502 550692 25508
rect 547144 18012 547196 18018
rect 547144 17954 547196 17960
rect 549260 18012 549312 18018
rect 549260 17954 549312 17960
rect 548892 4820 548944 4826
rect 548892 4762 548944 4768
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 546604 3454 547736 3482
rect 543004 3324 543056 3330
rect 543004 3266 543056 3272
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546500 3324 546552 3330
rect 546500 3266 546552 3272
rect 546512 480 546540 3266
rect 547708 480 547736 3454
rect 548904 480 548932 4762
rect 549272 3482 549300 17954
rect 550652 3482 550680 25502
rect 552020 22772 552072 22778
rect 552020 22714 552072 22720
rect 552032 3482 552060 22714
rect 552768 7614 552796 151778
rect 553400 72480 553452 72486
rect 553400 72422 553452 72428
rect 553124 29232 553176 29238
rect 553122 29200 553124 29209
rect 553176 29200 553178 29209
rect 553122 29135 553178 29144
rect 552756 7608 552808 7614
rect 552756 7550 552808 7556
rect 553412 3482 553440 72422
rect 554056 4826 554084 187682
rect 554044 4820 554096 4826
rect 554044 4762 554096 4768
rect 554792 3534 554820 604590
rect 558918 604551 558974 604560
rect 556160 600636 556212 600642
rect 556160 600578 556212 600584
rect 554872 6384 554924 6390
rect 554872 6326 554924 6332
rect 554780 3528 554832 3534
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 554780 3470 554832 3476
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554884 3346 554912 6326
rect 555976 3528 556028 3534
rect 555976 3470 556028 3476
rect 556172 3482 556200 600578
rect 558184 316056 558236 316062
rect 558184 315998 558236 316004
rect 558196 85542 558224 315998
rect 558184 85536 558236 85542
rect 558184 85478 558236 85484
rect 558368 6316 558420 6322
rect 558368 6258 558420 6264
rect 554792 3318 554912 3346
rect 554792 480 554820 3318
rect 555988 480 556016 3470
rect 556172 3454 557212 3482
rect 557184 480 557212 3454
rect 558380 480 558408 6258
rect 558932 3482 558960 604551
rect 563702 604480 563758 604489
rect 563702 604415 563758 604424
rect 560944 579692 560996 579698
rect 560944 579634 560996 579640
rect 560956 100570 560984 579634
rect 560944 100564 560996 100570
rect 560944 100506 560996 100512
rect 563058 93120 563114 93129
rect 563058 93055 563114 93064
rect 560206 29336 560262 29345
rect 560206 29271 560262 29280
rect 560220 29238 560248 29271
rect 560208 29232 560260 29238
rect 560208 29174 560260 29180
rect 560300 14476 560352 14482
rect 560300 14418 560352 14424
rect 560312 3482 560340 14418
rect 561956 6248 562008 6254
rect 561956 6190 562008 6196
rect 558932 3454 559604 3482
rect 560312 3454 560800 3482
rect 559576 480 559604 3454
rect 560772 480 560800 3454
rect 561968 480 561996 6190
rect 563072 3482 563100 93055
rect 563716 17950 563744 604415
rect 572626 603800 572682 603809
rect 572810 603800 572866 603809
rect 572682 603758 572810 603786
rect 572626 603735 572682 603744
rect 572810 603735 572866 603744
rect 569960 602132 570012 602138
rect 569960 602074 570012 602080
rect 569316 556232 569368 556238
rect 569316 556174 569368 556180
rect 565084 541680 565136 541686
rect 565084 541622 565136 541628
rect 565096 510610 565124 541622
rect 565084 510604 565136 510610
rect 565084 510546 565136 510552
rect 567844 485852 567896 485858
rect 567844 485794 567896 485800
rect 565084 462392 565136 462398
rect 565084 462334 565136 462340
rect 565096 96626 565124 462334
rect 567856 306338 567884 485794
rect 569224 357468 569276 357474
rect 569224 357410 569276 357416
rect 567844 306332 567896 306338
rect 567844 306274 567896 306280
rect 567844 251252 567896 251258
rect 567844 251194 567896 251200
rect 567856 97986 567884 251194
rect 569236 100881 569264 357410
rect 569328 335306 569356 556174
rect 569316 335300 569368 335306
rect 569316 335242 569368 335248
rect 569222 100872 569278 100881
rect 569222 100807 569278 100816
rect 567844 97980 567896 97986
rect 567844 97922 567896 97928
rect 565084 96620 565136 96626
rect 565084 96562 565136 96568
rect 567200 94512 567252 94518
rect 567200 94454 567252 94460
rect 564440 85536 564492 85542
rect 564440 85478 564492 85484
rect 563704 17944 563756 17950
rect 563704 17886 563756 17892
rect 564348 7608 564400 7614
rect 564348 7550 564400 7556
rect 563072 3454 563192 3482
rect 563164 480 563192 3454
rect 564360 480 564388 7550
rect 564452 3482 564480 85478
rect 565820 44872 565872 44878
rect 565820 44814 565872 44820
rect 565832 3482 565860 44814
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567212 3346 567240 94454
rect 569040 6180 569092 6186
rect 569040 6122 569092 6128
rect 567212 3318 567884 3346
rect 567856 480 567884 3318
rect 569052 480 569080 6122
rect 569972 3346 570000 602074
rect 571984 487212 572036 487218
rect 571984 487154 572036 487160
rect 571340 11892 571392 11898
rect 571340 11834 571392 11840
rect 571352 3482 571380 11834
rect 571996 5574 572024 487154
rect 572628 6452 572680 6458
rect 572628 6394 572680 6400
rect 571984 5568 572036 5574
rect 571984 5510 572036 5516
rect 571352 3454 571472 3482
rect 569972 3318 570276 3346
rect 570248 480 570276 3318
rect 571444 480 571472 3454
rect 572640 480 572668 6394
rect 573376 3466 573404 605950
rect 580264 602404 580316 602410
rect 580264 602346 580316 602352
rect 579894 592512 579950 592521
rect 579894 592447 579950 592456
rect 579908 592074 579936 592447
rect 579896 592068 579948 592074
rect 579896 592010 579948 592016
rect 574100 582412 574152 582418
rect 574100 582354 574152 582360
rect 573456 389224 573508 389230
rect 573456 389166 573508 389172
rect 573468 158710 573496 389166
rect 573456 158704 573508 158710
rect 573456 158646 573508 158652
rect 573824 8968 573876 8974
rect 573824 8910 573876 8916
rect 573364 3460 573416 3466
rect 573364 3402 573416 3408
rect 573836 480 573864 8910
rect 574112 3346 574140 582354
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 579894 545592 579950 545601
rect 579894 545527 579950 545536
rect 579908 545154 579936 545527
rect 579896 545148 579948 545154
rect 579896 545090 579948 545096
rect 580172 534064 580224 534070
rect 580172 534006 580224 534012
rect 580184 533905 580212 534006
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580172 510604 580224 510610
rect 580172 510546 580224 510552
rect 580184 510377 580212 510546
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580172 499520 580224 499526
rect 580172 499462 580224 499468
rect 580184 498681 580212 499462
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580172 452600 580224 452606
rect 580172 452542 580224 452548
rect 580184 451761 580212 452542
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 579620 440224 579672 440230
rect 579620 440166 579672 440172
rect 579632 439929 579660 440166
rect 579618 439920 579674 439929
rect 579618 439855 579674 439864
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580172 393304 580224 393310
rect 580172 393246 580224 393252
rect 580184 393009 580212 393246
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 580184 357474 580212 357847
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 580276 346089 580304 602346
rect 580356 599616 580408 599622
rect 580356 599558 580408 599564
rect 580368 416537 580396 599558
rect 580354 416528 580410 416537
rect 580354 416463 580410 416472
rect 580262 346080 580318 346089
rect 580262 346015 580318 346024
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 251258 580212 252175
rect 580172 251252 580224 251258
rect 580172 251194 580224 251200
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580184 204338 580212 205255
rect 580172 204332 580224 204338
rect 580172 204274 580224 204280
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 580262 111480 580318 111489
rect 580262 111415 580318 111424
rect 580276 102105 580304 111415
rect 580262 102096 580318 102105
rect 580262 102031 580318 102040
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 574744 33856 574796 33862
rect 574744 33798 574796 33804
rect 574756 3602 574784 33798
rect 581092 28280 581144 28286
rect 581092 28222 581144 28228
rect 576860 21480 576912 21486
rect 576860 21422 576912 21428
rect 576216 5568 576268 5574
rect 576216 5510 576268 5516
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 574112 3318 575060 3346
rect 575032 480 575060 3318
rect 576228 480 576256 5510
rect 576872 610 576900 21422
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 578608 4820 578660 4826
rect 578608 4762 578660 4768
rect 576860 604 576912 610
rect 576860 546 576912 552
rect 577412 604 577464 610
rect 577412 546 577464 552
rect 577424 480 577452 546
rect 578620 480 578648 4762
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3470
rect 581104 610 581132 28222
rect 581092 604 581144 610
rect 581092 546 581144 552
rect 582196 604 582248 610
rect 582196 546 582248 552
rect 582208 480 582236 546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 2870 595992 2926 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 3422 538600 3478 538656
rect 3146 509904 3202 509960
rect 3422 495488 3478 495544
rect 3790 481072 3846 481128
rect 3422 437960 3478 438016
rect 3238 423680 3294 423736
rect 3330 394984 3386 395040
rect 3422 380568 3478 380624
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 3422 308760 3478 308816
rect 3422 294344 3478 294400
rect 3422 280064 3478 280120
rect 3422 278840 3478 278896
rect 3422 265648 3478 265704
rect 3422 251252 3478 251288
rect 3422 251232 3424 251252
rect 3424 251232 3476 251252
rect 3476 251232 3478 251252
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 3422 208120 3478 208176
rect 3146 193840 3202 193896
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3514 136312 3570 136368
rect 3422 122032 3478 122088
rect 4066 107652 4068 107672
rect 4068 107652 4120 107672
rect 4120 107652 4122 107672
rect 4066 107616 4122 107652
rect 3422 93200 3478 93256
rect 3422 80008 3478 80064
rect 3422 78920 3478 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3146 21392 3202 21448
rect 3422 7112 3478 7168
rect 5262 2760 5318 2816
rect 13082 600480 13138 600536
rect 13634 30912 13690 30968
rect 16026 8880 16082 8936
rect 24674 600616 24730 600672
rect 23110 3712 23166 3768
rect 24766 102040 24822 102096
rect 35806 595448 35862 595504
rect 33046 24112 33102 24168
rect 48226 601840 48282 601896
rect 46846 9016 46902 9072
rect 52366 601704 52422 601760
rect 53746 600344 53802 600400
rect 55218 4800 55274 4856
rect 59174 601024 59230 601080
rect 59174 101632 59230 101688
rect 60646 602248 60702 602304
rect 64234 39208 64290 39264
rect 64602 11600 64658 11656
rect 67086 604016 67142 604072
rect 66994 578176 67050 578232
rect 66994 572600 67050 572656
rect 66994 534248 67050 534304
rect 66994 531528 67050 531584
rect 66534 521600 66590 521656
rect 66534 512216 66590 512272
rect 66626 510312 66682 510368
rect 66626 500928 66682 500984
rect 66994 491136 67050 491192
rect 66994 483656 67050 483712
rect 66994 478760 67050 478816
rect 66994 469376 67050 469432
rect 66902 469104 66958 469160
rect 66902 459720 66958 459776
rect 66718 446392 66774 446448
rect 66718 434696 66774 434752
rect 66994 434560 67050 434616
rect 66994 429800 67050 429856
rect 66902 398928 66958 398984
rect 66902 396072 66958 396128
rect 66994 383424 67050 383480
rect 66994 374040 67050 374096
rect 66718 336504 66774 336560
rect 66902 328344 66958 328400
rect 66718 327256 66774 327312
rect 66902 323584 66958 323640
rect 66994 299240 67050 299296
rect 66994 289992 67050 290048
rect 66902 280064 66958 280120
rect 66902 270680 66958 270736
rect 66718 201320 66774 201376
rect 66718 195472 66774 195528
rect 67086 240080 67142 240136
rect 67086 222400 67142 222456
rect 67086 205944 67142 206000
rect 67086 205400 67142 205456
rect 67086 191528 67142 191584
rect 67086 174120 67142 174176
rect 67086 114416 67142 114472
rect 67086 113328 67142 113384
rect 67086 103264 67142 103320
rect 67086 89664 67142 89720
rect 67270 72392 67326 72448
rect 67270 67632 67326 67688
rect 67086 57840 67142 57896
rect 67086 50904 67142 50960
rect 67454 100408 67510 100464
rect 69662 3848 69718 3904
rect 67178 3440 67234 3496
rect 71410 599936 71466 599992
rect 72330 190440 72386 190496
rect 71686 3576 71742 3632
rect 71318 3304 71374 3360
rect 74170 600752 74226 600808
rect 73066 190440 73122 190496
rect 72882 101360 72938 101416
rect 73802 101496 73858 101552
rect 73066 9152 73122 9208
rect 73250 3848 73306 3904
rect 73066 3440 73122 3496
rect 73250 3440 73306 3496
rect 75182 102720 75238 102776
rect 76470 205944 76526 206000
rect 76470 205400 76526 205456
rect 76930 101904 76986 101960
rect 78678 599528 78734 599584
rect 78678 595720 78734 595776
rect 78678 592184 78734 592240
rect 78954 577496 79010 577552
rect 78770 573960 78826 574016
rect 78678 570152 78734 570208
rect 78678 566616 78734 566672
rect 78678 562808 78734 562864
rect 78678 555736 78734 555792
rect 78678 526360 78734 526416
rect 78862 519016 78918 519072
rect 78678 511672 78734 511728
rect 78678 508136 78734 508192
rect 78678 504600 78734 504656
rect 79046 500792 79102 500848
rect 78678 497256 78734 497312
rect 78678 486104 78734 486160
rect 78678 479032 78734 479088
rect 78678 471688 78734 471744
rect 78678 460536 78734 460592
rect 78678 457000 78734 457056
rect 78678 449656 78734 449712
rect 78678 446120 78734 446176
rect 78678 442312 78734 442368
rect 78494 438776 78550 438832
rect 78402 394984 78458 395040
rect 78218 307128 78274 307184
rect 78126 303592 78182 303648
rect 77942 197784 77998 197840
rect 77206 100544 77262 100600
rect 78034 161064 78090 161120
rect 77206 90344 77262 90400
rect 75458 3712 75514 3768
rect 78586 434968 78642 435024
rect 78678 431432 78734 431488
rect 78678 427896 78734 427952
rect 78678 420552 78734 420608
rect 78678 416780 78680 416800
rect 78680 416780 78732 416800
rect 78732 416780 78734 416800
rect 78678 416744 78734 416780
rect 78678 413208 78734 413264
rect 78678 405864 78734 405920
rect 78678 402328 78734 402384
rect 78678 398520 78734 398576
rect 78678 387640 78734 387696
rect 78678 383832 78734 383888
rect 78678 369416 78734 369472
rect 78678 362072 78734 362128
rect 78678 358264 78734 358320
rect 78678 351192 78734 351248
rect 78678 347384 78734 347440
rect 78678 336504 78734 336560
rect 78678 332696 78734 332752
rect 78678 329160 78734 329216
rect 78678 325624 78734 325680
rect 78678 321816 78734 321872
rect 78678 318280 78734 318336
rect 78678 310936 78734 310992
rect 79230 300056 79286 300112
rect 78678 296248 78734 296304
rect 78678 292712 78734 292768
rect 78678 281580 78734 281616
rect 78678 281560 78680 281580
rect 78680 281560 78732 281580
rect 78732 281560 78734 281580
rect 78678 278024 78734 278080
rect 78678 274488 78734 274544
rect 78678 267144 78734 267200
rect 78678 263336 78734 263392
rect 78678 252456 78734 252512
rect 78678 248920 78734 248976
rect 78678 241576 78734 241632
rect 78678 237768 78734 237824
rect 78678 234232 78734 234288
rect 78678 230424 78734 230480
rect 78678 223352 78734 223408
rect 78678 212200 78734 212256
rect 78678 208664 78734 208720
rect 78678 193976 78734 194032
rect 78678 190476 78680 190496
rect 78680 190476 78732 190496
rect 78732 190476 78734 190496
rect 78678 190440 78734 190476
rect 79230 186632 79286 186688
rect 78678 183096 78734 183152
rect 78678 179288 78734 179344
rect 78678 172216 78734 172272
rect 78678 164872 78734 164928
rect 78678 157528 78734 157584
rect 78678 153720 78734 153776
rect 78678 150184 78734 150240
rect 78678 146648 78734 146704
rect 78678 131960 78734 132016
rect 78678 128152 78734 128208
rect 79138 113736 79194 113792
rect 78678 109928 78734 109984
rect 79598 559272 79654 559328
rect 79874 530168 79930 530224
rect 79506 493448 79562 493504
rect 79874 391176 79930 391232
rect 79782 343848 79838 343904
rect 79690 259800 79746 259856
rect 79598 219544 79654 219600
rect 79414 187720 79470 187776
rect 79506 142840 79562 142896
rect 79414 124616 79470 124672
rect 80702 601296 80758 601352
rect 80702 600888 80758 600944
rect 80978 482568 81034 482624
rect 80886 340040 80942 340096
rect 80794 201320 80850 201376
rect 81438 464344 81494 464400
rect 81530 409400 81586 409456
rect 81714 380296 81770 380352
rect 81622 314472 81678 314528
rect 81622 270680 81678 270736
rect 81714 216008 81770 216064
rect 81806 168408 81862 168464
rect 82082 155216 82138 155272
rect 83370 601296 83426 601352
rect 93766 605920 93822 605976
rect 88338 602248 88394 602304
rect 83370 600344 83426 600400
rect 92386 601296 92442 601352
rect 103702 604424 103758 604480
rect 267646 700304 267702 700360
rect 169758 683168 169814 683224
rect 170126 683168 170182 683224
rect 188342 674056 188398 674112
rect 173898 673956 173900 673976
rect 173900 673956 173952 673976
rect 173952 673956 173954 673976
rect 173898 673920 173954 673956
rect 154578 673804 154634 673840
rect 154578 673784 154580 673804
rect 154580 673784 154632 673804
rect 154632 673784 154634 673804
rect 166906 673784 166962 673840
rect 178314 673784 178370 673840
rect 188342 673784 188398 673840
rect 162214 673512 162270 673568
rect 166906 673512 166962 673568
rect 118790 603880 118846 603936
rect 118606 603744 118662 603800
rect 104898 601840 104954 601896
rect 138294 604560 138350 604616
rect 138110 603880 138166 603936
rect 137926 603744 137982 603800
rect 149610 603880 149666 603936
rect 149702 603744 149758 603800
rect 157982 604696 158038 604752
rect 168286 605956 168288 605976
rect 168288 605956 168340 605976
rect 168340 605956 168342 605976
rect 168286 605920 168342 605956
rect 170310 603472 170366 603528
rect 185214 605920 185270 605976
rect 190090 604832 190146 604888
rect 196070 604016 196126 604072
rect 195886 603744 195942 603800
rect 219806 606056 219862 606112
rect 212262 603472 212318 603528
rect 494794 700304 494850 700360
rect 293958 607416 294014 607472
rect 281446 607280 281502 607336
rect 267094 601840 267150 601896
rect 289818 604052 289820 604072
rect 289820 604052 289872 604072
rect 289872 604052 289874 604072
rect 289818 604016 289874 604052
rect 286414 602112 286470 602168
rect 288990 602112 289046 602168
rect 298742 604832 298798 604888
rect 309138 604016 309194 604072
rect 299386 603744 299442 603800
rect 330942 607552 330998 607608
rect 315946 601976 316002 602032
rect 318706 603744 318762 603800
rect 318798 602248 318854 602304
rect 328458 604052 328460 604072
rect 328460 604052 328512 604072
rect 328512 604052 328514 604072
rect 328458 604016 328514 604052
rect 335910 606192 335966 606248
rect 338026 603744 338082 603800
rect 347778 604052 347780 604072
rect 347780 604052 347832 604072
rect 347832 604052 347834 604072
rect 347778 604016 347834 604052
rect 350630 603608 350686 603664
rect 346398 602384 346454 602440
rect 357346 603880 357402 603936
rect 369674 603744 369730 603800
rect 369950 603744 370006 603800
rect 379426 603744 379482 603800
rect 379610 603608 379666 603664
rect 397734 606464 397790 606520
rect 385222 606328 385278 606384
rect 392766 604968 392822 605024
rect 439686 604152 439742 604208
rect 429750 603336 429806 603392
rect 444378 603608 444434 603664
rect 442078 603336 442134 603392
rect 449162 603764 449218 603800
rect 449162 603744 449164 603764
rect 449164 603744 449216 603764
rect 449216 603744 449218 603764
rect 447046 603200 447102 603256
rect 449622 603200 449678 603256
rect 463606 604152 463662 604208
rect 463606 603880 463662 603936
rect 488998 604016 489054 604072
rect 483018 603900 483074 603936
rect 483018 603880 483020 603900
rect 483020 603880 483072 603900
rect 483072 603880 483074 603900
rect 473266 603744 473322 603800
rect 473266 603608 473322 603664
rect 481822 602012 481824 602032
rect 481824 602012 481876 602032
rect 481876 602012 481878 602032
rect 481822 601976 481878 602012
rect 491574 603336 491630 603392
rect 492770 603900 492826 603936
rect 492770 603880 492772 603900
rect 492772 603880 492824 603900
rect 492824 603880 492826 603900
rect 498934 603064 498990 603120
rect 367650 601704 367706 601760
rect 427726 601704 427782 601760
rect 162858 601296 162914 601352
rect 195334 601296 195390 601352
rect 207202 601296 207258 601352
rect 249706 601296 249762 601352
rect 278778 601296 278834 601352
rect 296074 601296 296130 601352
rect 306010 601296 306066 601352
rect 402886 601296 402942 601352
rect 405462 601296 405518 601352
rect 415398 601296 415454 601352
rect 435086 601296 435142 601352
rect 476946 601296 477002 601352
rect 486330 601296 486386 601352
rect 496266 601296 496322 601352
rect 501510 600244 501512 600264
rect 501512 600244 501564 600264
rect 501564 600244 501566 600264
rect 501510 600208 501566 600244
rect 501510 589464 501566 589520
rect 82634 452920 82690 452976
rect 82634 175344 82690 175400
rect 82542 138760 82598 138816
rect 82634 134952 82690 135008
rect 82174 120536 82230 120592
rect 81990 117000 82046 117056
rect 82634 106700 82636 106720
rect 82636 106700 82688 106720
rect 82688 106700 82690 106720
rect 82634 106664 82690 106700
rect 502338 535336 502394 535392
rect 501786 526360 501842 526416
rect 501878 524728 501934 524784
rect 501786 522824 501842 522880
rect 501878 522280 501934 522336
rect 502062 507728 502118 507784
rect 502062 498344 502118 498400
rect 501970 481480 502026 481536
rect 501970 471960 502026 472016
rect 502062 471824 502118 471880
rect 502062 462576 502118 462632
rect 501970 458904 502026 458960
rect 501970 452648 502026 452704
rect 502338 451288 502394 451344
rect 502062 442856 502118 442912
rect 502062 433336 502118 433392
rect 501694 430616 501750 430672
rect 501878 430480 501934 430536
rect 502062 428440 502118 428496
rect 501970 415384 502026 415440
rect 502062 413888 502118 413944
rect 502062 404504 502118 404560
rect 502062 394576 502118 394632
rect 502062 385192 502118 385248
rect 502062 360848 502118 360904
rect 502062 356088 502118 356144
rect 502246 354592 502302 354648
rect 502246 345208 502302 345264
rect 502062 335280 502118 335336
rect 501694 327528 501750 327584
rect 502062 325760 502118 325816
rect 501602 321408 501658 321464
rect 501602 312024 501658 312080
rect 501602 308216 501658 308272
rect 501510 137808 501566 137864
rect 501510 136584 501566 136640
rect 108946 102584 109002 102640
rect 109130 102584 109186 102640
rect 118422 102584 118478 102640
rect 118606 102584 118662 102640
rect 125506 102584 125562 102640
rect 133694 102584 133750 102640
rect 133878 102584 133934 102640
rect 84014 102448 84070 102504
rect 133970 102448 134026 102504
rect 84106 75112 84162 75168
rect 85578 101904 85634 101960
rect 88338 102040 88394 102096
rect 87326 100408 87382 100464
rect 89994 101632 90050 101688
rect 89902 77288 89958 77344
rect 90086 77288 90142 77344
rect 99194 26832 99250 26888
rect 116122 101496 116178 101552
rect 115754 50224 115810 50280
rect 124494 100544 124550 100600
rect 120078 98912 120134 98968
rect 131210 101360 131266 101416
rect 129738 98640 129794 98696
rect 135166 79328 135222 79384
rect 133694 2760 133750 2816
rect 135258 5772 135314 5808
rect 135258 5752 135260 5772
rect 135260 5752 135312 5772
rect 135312 5752 135314 5772
rect 141790 100680 141846 100736
rect 138018 86944 138074 87000
rect 140778 86944 140834 87000
rect 140502 77152 140558 77208
rect 140778 77152 140834 77208
rect 140502 67632 140558 67688
rect 140778 67632 140834 67688
rect 140686 44784 140742 44840
rect 145010 5616 145066 5672
rect 148966 36488 149022 36544
rect 161478 97824 161534 97880
rect 164146 95784 164202 95840
rect 162766 5888 162822 5944
rect 162766 5480 162822 5536
rect 163042 5480 163098 5536
rect 162950 5344 163006 5400
rect 171414 100680 171470 100736
rect 169390 3984 169446 4040
rect 176566 101360 176622 101416
rect 176750 102584 176806 102640
rect 182178 5652 182180 5672
rect 182180 5652 182232 5672
rect 182232 5652 182234 5672
rect 182178 5616 182234 5652
rect 193678 100816 193734 100872
rect 190366 46144 190422 46200
rect 198370 96600 198426 96656
rect 198738 96600 198794 96656
rect 199934 5752 199990 5808
rect 307666 102584 307722 102640
rect 274546 102448 274602 102504
rect 201590 5924 201592 5944
rect 201592 5924 201644 5944
rect 201644 5924 201646 5944
rect 201590 5888 201646 5924
rect 212262 101496 212318 101552
rect 209686 87624 209742 87680
rect 211066 5924 211068 5944
rect 211068 5924 211120 5944
rect 211120 5924 211122 5944
rect 211066 5888 211122 5924
rect 213918 86264 213974 86320
rect 220634 6024 220690 6080
rect 220634 5344 220690 5400
rect 237286 98640 237342 98696
rect 242806 97144 242862 97200
rect 248326 72392 248382 72448
rect 253754 9288 253810 9344
rect 263414 86264 263470 86320
rect 259366 6024 259422 6080
rect 259366 5616 259422 5672
rect 263322 3576 263378 3632
rect 266174 71168 266230 71224
rect 266358 71304 266414 71360
rect 273902 5752 273958 5808
rect 273902 5480 273958 5536
rect 280250 77152 280306 77208
rect 280434 77152 280490 77208
rect 282826 5752 282882 5808
rect 283010 5752 283066 5808
rect 289726 98912 289782 98968
rect 295522 7520 295578 7576
rect 299110 3440 299166 3496
rect 304906 97280 304962 97336
rect 309138 94424 309194 94480
rect 319994 95920 320050 95976
rect 317326 51720 317382 51776
rect 324226 101768 324282 101824
rect 322846 101632 322902 101688
rect 325238 6296 325294 6352
rect 330850 5752 330906 5808
rect 330942 5616 330998 5672
rect 331218 98776 331274 98832
rect 340786 57160 340842 57216
rect 344926 98776 344982 98832
rect 346674 9288 346730 9344
rect 350446 5616 350502 5672
rect 350630 5616 350686 5672
rect 357346 96056 357402 96112
rect 369214 9016 369270 9072
rect 375286 5752 375342 5808
rect 375286 5480 375342 5536
rect 381174 3440 381230 3496
rect 386418 11736 386474 11792
rect 389178 53080 389234 53136
rect 390650 9152 390706 9208
rect 395434 9016 395490 9072
rect 394606 6024 394662 6080
rect 394606 5616 394662 5672
rect 406382 99048 406438 99104
rect 400126 50360 400182 50416
rect 403714 6432 403770 6488
rect 409878 35128 409934 35184
rect 407302 6296 407358 6352
rect 409878 29144 409934 29200
rect 414018 29008 414074 29064
rect 411166 19352 411222 19408
rect 411350 19352 411406 19408
rect 415398 6568 415454 6624
rect 415398 6024 415454 6080
rect 483018 102176 483074 102232
rect 423402 96600 423458 96656
rect 423586 96600 423642 96656
rect 422206 82048 422262 82104
rect 424966 6568 425022 6624
rect 424966 6024 425022 6080
rect 426438 66816 426494 66872
rect 425150 6568 425206 6624
rect 433430 47504 433486 47560
rect 437570 71032 437626 71088
rect 438122 5772 438178 5808
rect 438122 5752 438124 5772
rect 438124 5752 438176 5772
rect 438176 5752 438178 5772
rect 445482 96600 445538 96656
rect 445666 96600 445722 96656
rect 442906 5772 442962 5808
rect 442906 5752 442908 5772
rect 442908 5752 442960 5772
rect 442960 5752 442962 5772
rect 448518 86128 448574 86184
rect 447046 5752 447102 5808
rect 447230 5616 447286 5672
rect 451370 3712 451426 3768
rect 450174 3576 450230 3632
rect 454038 90480 454094 90536
rect 458178 59880 458234 59936
rect 468482 5888 468538 5944
rect 468482 5480 468538 5536
rect 464434 3848 464490 3904
rect 465630 2760 465686 2816
rect 471518 6704 471574 6760
rect 480166 96464 480222 96520
rect 483018 97280 483074 97336
rect 481638 77832 481694 77888
rect 481822 5924 481824 5944
rect 481824 5924 481876 5944
rect 481876 5924 481878 5944
rect 481822 5888 481878 5924
rect 484490 96600 484546 96656
rect 488630 96600 488686 96656
rect 492862 102040 492918 102096
rect 492862 96056 492918 96112
rect 495254 102040 495310 102096
rect 494150 101904 494206 101960
rect 491206 5924 491208 5944
rect 491208 5924 491260 5944
rect 491260 5924 491262 5944
rect 491206 5888 491262 5924
rect 489366 3984 489422 4040
rect 490562 3712 490618 3768
rect 499118 100680 499174 100736
rect 499118 67632 499174 67688
rect 499210 66952 499266 67008
rect 499210 60016 499266 60072
rect 499210 55120 499266 55176
rect 499210 45736 499266 45792
rect 496358 45464 496414 45520
rect 499210 45464 499266 45520
rect 496358 40704 496414 40760
rect 499210 40704 499266 40760
rect 498382 28736 498438 28792
rect 498382 21120 498438 21176
rect 500498 87624 500554 87680
rect 500498 82048 500554 82104
rect 500038 45464 500094 45520
rect 500038 39208 500094 39264
rect 501786 279112 501842 279168
rect 501694 271904 501750 271960
rect 501970 228792 502026 228848
rect 501970 220904 502026 220960
rect 501878 183912 501934 183968
rect 501970 126928 502026 126984
rect 501878 122712 501934 122768
rect 501878 121896 501934 121952
rect 501970 119312 502026 119368
rect 502430 414840 502486 414896
rect 502522 411032 502578 411088
rect 502430 312568 502486 312624
rect 502614 352552 502670 352608
rect 502706 264968 502762 265024
rect 503626 254360 503682 254416
rect 503626 253816 503682 253872
rect 502890 217640 502946 217696
rect 502798 159160 502854 159216
rect 503902 593816 503958 593872
rect 503902 586508 503904 586528
rect 503904 586508 503956 586528
rect 503956 586508 503958 586528
rect 503902 586472 503958 586508
rect 503902 582664 503958 582720
rect 504454 575592 504510 575648
rect 503902 571784 503958 571840
rect 504362 569880 504418 569936
rect 503902 568248 503958 568304
rect 503902 564460 503958 564496
rect 503902 564440 503904 564460
rect 503904 564440 503956 564460
rect 503956 564440 503958 564460
rect 503902 560904 503958 560960
rect 503902 553560 503958 553616
rect 503902 550024 503958 550080
rect 503902 546216 503958 546272
rect 504546 569880 504602 569936
rect 503902 542680 503958 542736
rect 503902 538872 503958 538928
rect 503902 524476 503958 524512
rect 503902 524456 503904 524476
rect 503904 524456 503956 524476
rect 503956 524456 503958 524476
rect 503902 520648 503958 520704
rect 503902 498888 503958 498944
rect 503902 495080 503958 495136
rect 504178 492632 504234 492688
rect 504362 492632 504418 492688
rect 503902 487736 503958 487792
rect 503902 484200 503958 484256
rect 503902 476856 503958 476912
rect 503902 473356 503904 473376
rect 503904 473356 503956 473376
rect 503956 473356 503958 473376
rect 503902 473320 503958 473356
rect 503902 469512 503958 469568
rect 504454 473320 504510 473376
rect 504638 473320 504694 473376
rect 503902 462168 503958 462224
rect 504178 454008 504234 454064
rect 504362 454008 504418 454064
rect 503902 447752 503958 447808
rect 503902 443944 503958 444000
rect 503902 440408 503958 440464
rect 503902 436600 503958 436656
rect 503902 433064 503958 433120
rect 503902 429256 503958 429312
rect 503902 425720 503958 425776
rect 503902 422184 503958 422240
rect 503902 407496 503958 407552
rect 503902 403688 503958 403744
rect 503902 400152 503958 400208
rect 505098 396616 505154 396672
rect 504454 396072 504510 396128
rect 504638 396072 504694 396128
rect 503902 389272 503958 389328
rect 503902 385464 503958 385520
rect 503902 381928 503958 381984
rect 503902 378156 503904 378176
rect 503904 378156 503956 378176
rect 503956 378156 503958 378176
rect 503902 378120 503958 378156
rect 503902 374584 503958 374640
rect 503902 371048 503958 371104
rect 503810 181192 503866 181248
rect 503810 177384 503866 177440
rect 503718 173984 503774 174040
rect 503718 170040 503774 170096
rect 503718 166504 503774 166560
rect 503718 151836 503774 151872
rect 503718 151816 503720 151836
rect 503720 151816 503772 151836
rect 503772 151816 503774 151836
rect 503718 148008 503774 148064
rect 503074 133592 503130 133648
rect 503258 111560 503314 111616
rect 503350 108024 503406 108080
rect 503994 367240 504050 367296
rect 503994 363704 504050 363760
rect 503994 359896 504050 359952
rect 504086 345480 504142 345536
rect 504086 341672 504142 341728
rect 504086 338156 504142 338192
rect 504086 338136 504088 338156
rect 504088 338136 504140 338156
rect 504140 338136 504142 338156
rect 504086 334328 504142 334384
rect 504086 323448 504142 323504
rect 504086 319912 504142 319968
rect 504086 316104 504142 316160
rect 504086 305224 504142 305280
rect 504086 294344 504142 294400
rect 504086 290536 504142 290592
rect 504086 287000 504142 287056
rect 504178 283328 504234 283384
rect 504086 283192 504142 283248
rect 504178 280336 504234 280392
rect 504086 275848 504142 275904
rect 504086 268776 504142 268832
rect 504086 261432 504142 261488
rect 504086 257624 504142 257680
rect 504086 250280 504142 250336
rect 504086 246744 504142 246800
rect 504086 243208 504142 243264
rect 504086 235864 504142 235920
rect 504086 232056 504142 232112
rect 504086 228520 504142 228576
rect 504086 224712 504142 224768
rect 504086 221176 504142 221232
rect 504086 213832 504142 213888
rect 504086 210296 504142 210352
rect 504086 202952 504142 203008
rect 503994 151136 504050 151192
rect 503994 118904 504050 118960
rect 504178 195608 504234 195664
rect 504270 194384 504326 194440
rect 504178 188264 504234 188320
rect 504270 186224 504326 186280
rect 504270 185272 504326 185328
rect 504178 185136 504234 185192
rect 504270 184728 504326 184784
rect 504178 176568 504234 176624
rect 504178 175344 504234 175400
rect 504178 173576 504234 173632
rect 504362 175072 504418 175128
rect 504362 165824 504418 165880
rect 504454 162696 504510 162752
rect 504546 144472 504602 144528
rect 504546 140936 504602 140992
rect 504546 126248 504602 126304
rect 504546 104216 504602 104272
rect 505190 392808 505246 392864
rect 505282 356360 505338 356416
rect 505374 330792 505430 330848
rect 505466 301416 505522 301472
rect 505558 254088 505614 254144
rect 505650 180920 505706 180976
rect 505742 129784 505798 129840
rect 504822 3304 504878 3360
rect 509330 98912 509386 98968
rect 509238 69536 509294 69592
rect 510710 603200 510766 603256
rect 511446 87488 511502 87544
rect 512826 570152 512882 570208
rect 512826 570016 512882 570072
rect 512826 568520 512882 568576
rect 513010 568520 513066 568576
rect 512826 549208 512882 549264
rect 513010 549208 513066 549264
rect 512826 500928 512882 500984
rect 513010 500928 513066 500984
rect 512826 278704 512882 278760
rect 513010 278704 513066 278760
rect 512826 259392 512882 259448
rect 513010 259392 513066 259448
rect 512826 240080 512882 240136
rect 513010 240080 513066 240136
rect 512826 220768 512882 220824
rect 513010 220768 513066 220824
rect 512826 211112 512882 211168
rect 513010 211112 513066 211168
rect 512826 191800 512882 191856
rect 513010 191800 513066 191856
rect 512826 172488 512882 172544
rect 513010 172488 513066 172544
rect 514942 95784 514998 95840
rect 516138 603472 516194 603528
rect 514666 5752 514722 5808
rect 514850 5752 514906 5808
rect 516874 603880 516930 603936
rect 517518 601840 517574 601896
rect 516598 101496 516654 101552
rect 516138 3712 516194 3768
rect 517886 603336 517942 603392
rect 520278 601976 520334 602032
rect 517886 101632 517942 101688
rect 517978 98640 518034 98696
rect 521566 199960 521622 200016
rect 521566 190440 521622 190496
rect 521934 579536 521990 579592
rect 521934 570152 521990 570208
rect 522118 560224 522174 560280
rect 522118 550704 522174 550760
rect 522026 540912 522082 540968
rect 522026 531528 522082 531584
rect 522026 521600 522082 521656
rect 522026 512216 522082 512272
rect 522026 502288 522082 502344
rect 522026 492632 522082 492688
rect 522118 463392 522174 463448
rect 522118 454008 522174 454064
rect 522210 424904 522266 424960
rect 522210 415384 522266 415440
rect 522210 405456 522266 405512
rect 522210 396072 522266 396128
rect 522210 386144 522266 386200
rect 522210 376760 522266 376816
rect 522210 357312 522266 357368
rect 522210 350512 522266 350568
rect 522210 347520 522266 347576
rect 522210 338136 522266 338192
rect 522210 328344 522266 328400
rect 522210 318960 522266 319016
rect 522210 308896 522266 308952
rect 522210 302096 522266 302152
rect 522210 289584 522266 289640
rect 522210 280336 522266 280392
rect 522210 270408 522266 270464
rect 522210 261024 522266 261080
rect 522210 251096 522266 251152
rect 522210 241712 522266 241768
rect 522210 222128 522266 222184
rect 522210 212608 522266 212664
rect 522210 212472 522266 212528
rect 522210 206216 522266 206272
rect 522210 173848 522266 173904
rect 522210 164192 522266 164248
rect 522302 135088 522358 135144
rect 522302 125568 522358 125624
rect 522210 115776 522266 115832
rect 522210 106256 522266 106312
rect 525706 603608 525762 603664
rect 580170 686296 580226 686352
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 540886 603744 540942 603800
rect 533986 603644 533988 603664
rect 533988 603644 534040 603664
rect 534040 603644 534042 603664
rect 533986 603608 534042 603644
rect 526442 5752 526498 5808
rect 526442 5480 526498 5536
rect 535734 3984 535790 4040
rect 536930 6160 536986 6216
rect 540886 181328 540942 181384
rect 540886 181056 540942 181112
rect 553122 29180 553124 29200
rect 553124 29180 553176 29200
rect 553176 29180 553178 29200
rect 553122 29144 553178 29180
rect 558918 604560 558974 604616
rect 563702 604424 563758 604480
rect 563058 93064 563114 93120
rect 560206 29280 560262 29336
rect 572626 603744 572682 603800
rect 572810 603744 572866 603800
rect 569222 100816 569278 100872
rect 579894 592456 579950 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 579894 545536 579950 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580170 451696 580226 451752
rect 579618 439864 579674 439920
rect 580170 404776 580226 404832
rect 580170 392944 580226 393000
rect 580170 369552 580226 369608
rect 580170 357856 580226 357912
rect 580354 416472 580410 416528
rect 580262 346024 580318 346080
rect 580170 322632 580226 322688
rect 580170 310800 580226 310856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 252184 580226 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 580170 205264 580226 205320
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 580262 111424 580318 111480
rect 580262 102040 580318 102096
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 579802 17584 579858 17640
<< metal3 >>
rect 68870 700300 68876 700364
rect 68940 700362 68946 700364
rect 267641 700362 267707 700365
rect 68940 700360 267707 700362
rect 68940 700304 267646 700360
rect 267702 700304 267707 700360
rect 68940 700302 267707 700304
rect 68940 700300 68946 700302
rect 267641 700299 267707 700302
rect 486366 700300 486372 700364
rect 486436 700362 486442 700364
rect 494789 700362 494855 700365
rect 486436 700360 494855 700362
rect 486436 700304 494794 700360
rect 494850 700304 494855 700360
rect 486436 700302 494855 700304
rect 486436 700300 486442 700302
rect 494789 700299 494855 700302
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 519486 697172 519492 697236
rect 519556 697234 519562 697236
rect 519556 697174 528570 697234
rect 519556 697172 519562 697174
rect 528510 697098 528570 697174
rect 538262 697174 547890 697234
rect 528510 697038 538138 697098
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 547830 697098 547890 697174
rect 557582 697174 567210 697234
rect 547830 697038 557458 697098
rect 538078 696902 538322 696962
rect 557398 696962 557458 697038
rect 557582 696962 557642 697174
rect 567150 697098 567210 697174
rect 567150 697038 576778 697098
rect 557398 696902 557642 696962
rect 576718 696962 576778 697038
rect 583342 696962 583402 697990
rect 583520 697900 584960 697990
rect 576718 696902 583402 696962
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 169753 683226 169819 683229
rect 170121 683226 170187 683229
rect 169753 683224 170187 683226
rect 169753 683168 169758 683224
rect 169814 683168 170126 683224
rect 170182 683168 170187 683224
rect 169753 683166 170187 683168
rect 169753 683163 169819 683166
rect 170121 683163 170187 683166
rect -960 682274 480 682364
rect -960 682214 674 682274
rect -960 682124 480 682214
rect 614 681866 674 682214
rect 512678 681866 512684 681868
rect 614 681806 512684 681866
rect 512678 681804 512684 681806
rect 512748 681804 512754 681868
rect 583520 674658 584960 674748
rect 583342 674598 584960 674658
rect 183502 674052 183508 674116
rect 183572 674114 183578 674116
rect 188337 674114 188403 674117
rect 183572 674112 188403 674114
rect 183572 674056 188342 674112
rect 188398 674056 188403 674112
rect 183572 674054 188403 674056
rect 183572 674052 183578 674054
rect 188337 674051 188403 674054
rect 173893 673978 173959 673981
rect 167318 673976 173959 673978
rect 167318 673920 173898 673976
rect 173954 673920 173959 673976
rect 167318 673918 173959 673920
rect 154573 673842 154639 673845
rect 79918 673782 84210 673842
rect 79918 673706 79978 673782
rect 70350 673646 79978 673706
rect 84150 673706 84210 673782
rect 93902 673782 103530 673842
rect 84150 673646 93778 673706
rect 70158 673508 70164 673572
rect 70228 673570 70234 673572
rect 70350 673570 70410 673646
rect 70228 673510 70410 673570
rect 93718 673570 93778 673646
rect 93902 673570 93962 673782
rect 103470 673706 103530 673782
rect 113222 673782 122850 673842
rect 103470 673646 113098 673706
rect 93718 673510 93962 673570
rect 113038 673570 113098 673646
rect 113222 673570 113282 673782
rect 122790 673706 122850 673782
rect 132542 673782 142170 673842
rect 122790 673646 132418 673706
rect 113038 673510 113282 673570
rect 132358 673570 132418 673646
rect 132542 673570 132602 673782
rect 142110 673706 142170 673782
rect 151862 673840 154639 673842
rect 151862 673784 154578 673840
rect 154634 673784 154639 673840
rect 151862 673782 154639 673784
rect 142110 673646 151738 673706
rect 132358 673510 132602 673570
rect 151678 673570 151738 673646
rect 151862 673570 151922 673782
rect 154573 673779 154639 673782
rect 166901 673842 166967 673845
rect 167318 673842 167378 673918
rect 173893 673915 173959 673918
rect 166901 673840 167378 673842
rect 166901 673784 166906 673840
rect 166962 673784 167378 673840
rect 166901 673782 167378 673784
rect 178309 673842 178375 673845
rect 183502 673842 183508 673844
rect 178309 673840 183508 673842
rect 178309 673784 178314 673840
rect 178370 673784 183508 673840
rect 178309 673782 183508 673784
rect 166901 673779 166967 673782
rect 178309 673779 178375 673782
rect 183502 673780 183508 673782
rect 183572 673780 183578 673844
rect 188337 673842 188403 673845
rect 188337 673840 200130 673842
rect 188337 673784 188342 673840
rect 188398 673784 200130 673840
rect 188337 673782 200130 673784
rect 188337 673779 188403 673782
rect 200070 673706 200130 673782
rect 209822 673782 219450 673842
rect 200070 673646 209698 673706
rect 151678 673510 151922 673570
rect 162209 673570 162275 673573
rect 166901 673570 166967 673573
rect 162209 673568 166967 673570
rect 162209 673512 162214 673568
rect 162270 673512 166906 673568
rect 166962 673512 166967 673568
rect 162209 673510 166967 673512
rect 209638 673570 209698 673646
rect 209822 673570 209882 673782
rect 219390 673706 219450 673782
rect 229142 673782 238770 673842
rect 219390 673646 229018 673706
rect 209638 673510 209882 673570
rect 228958 673570 229018 673646
rect 229142 673570 229202 673782
rect 238710 673706 238770 673782
rect 248462 673782 258090 673842
rect 238710 673646 248338 673706
rect 228958 673510 229202 673570
rect 248278 673570 248338 673646
rect 248462 673570 248522 673782
rect 258030 673706 258090 673782
rect 267782 673782 277410 673842
rect 258030 673646 267658 673706
rect 248278 673510 248522 673570
rect 267598 673570 267658 673646
rect 267782 673570 267842 673782
rect 277350 673706 277410 673782
rect 287102 673782 296730 673842
rect 277350 673646 286978 673706
rect 267598 673510 267842 673570
rect 286918 673570 286978 673646
rect 287102 673570 287162 673782
rect 296670 673706 296730 673782
rect 306422 673782 316050 673842
rect 296670 673646 306298 673706
rect 286918 673510 287162 673570
rect 306238 673570 306298 673646
rect 306422 673570 306482 673782
rect 315990 673706 316050 673782
rect 325742 673782 335370 673842
rect 315990 673646 325618 673706
rect 306238 673510 306482 673570
rect 325558 673570 325618 673646
rect 325742 673570 325802 673782
rect 335310 673706 335370 673782
rect 345062 673782 354690 673842
rect 335310 673646 344938 673706
rect 325558 673510 325802 673570
rect 344878 673570 344938 673646
rect 345062 673570 345122 673782
rect 354630 673706 354690 673782
rect 364382 673782 374010 673842
rect 354630 673646 364258 673706
rect 344878 673510 345122 673570
rect 364198 673570 364258 673646
rect 364382 673570 364442 673782
rect 373950 673706 374010 673782
rect 383702 673782 393330 673842
rect 373950 673646 383578 673706
rect 364198 673510 364442 673570
rect 383518 673570 383578 673646
rect 383702 673570 383762 673782
rect 393270 673706 393330 673782
rect 403022 673782 412650 673842
rect 393270 673646 402898 673706
rect 383518 673510 383762 673570
rect 402838 673570 402898 673646
rect 403022 673570 403082 673782
rect 412590 673706 412650 673782
rect 431910 673782 441538 673842
rect 412590 673646 422218 673706
rect 402838 673510 403082 673570
rect 422158 673570 422218 673646
rect 431910 673570 431970 673782
rect 422158 673510 431970 673570
rect 441478 673570 441538 673782
rect 441662 673782 451290 673842
rect 441662 673570 441722 673782
rect 451230 673706 451290 673782
rect 460982 673782 470610 673842
rect 451230 673646 460858 673706
rect 441478 673510 441722 673570
rect 460798 673570 460858 673646
rect 460982 673570 461042 673782
rect 470550 673706 470610 673782
rect 480302 673782 489930 673842
rect 470550 673646 480178 673706
rect 460798 673510 461042 673570
rect 480118 673570 480178 673646
rect 480302 673570 480362 673782
rect 489870 673706 489930 673782
rect 499622 673782 509250 673842
rect 489870 673646 499498 673706
rect 480118 673510 480362 673570
rect 499438 673570 499498 673646
rect 499622 673570 499682 673782
rect 509190 673706 509250 673782
rect 518942 673782 528570 673842
rect 509190 673646 518818 673706
rect 499438 673510 499682 673570
rect 518758 673570 518818 673646
rect 518942 673570 519002 673782
rect 528510 673706 528570 673782
rect 538262 673782 547890 673842
rect 528510 673646 538138 673706
rect 518758 673510 519002 673570
rect 538078 673570 538138 673646
rect 538262 673570 538322 673782
rect 547830 673706 547890 673782
rect 557582 673782 567210 673842
rect 547830 673646 557458 673706
rect 538078 673510 538322 673570
rect 557398 673570 557458 673646
rect 557582 673570 557642 673782
rect 567150 673706 567210 673782
rect 583342 673706 583402 674598
rect 583520 674508 584960 674598
rect 567150 673646 576778 673706
rect 557398 673510 557642 673570
rect 576718 673570 576778 673646
rect 576902 673646 583402 673706
rect 576902 673570 576962 673646
rect 576718 673510 576962 673570
rect 70228 673508 70234 673510
rect 162209 673507 162275 673510
rect 166901 673507 166967 673510
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 330937 607610 331003 607613
rect 489862 607610 489868 607612
rect 330937 607608 489868 607610
rect 330937 607552 330942 607608
rect 330998 607552 489868 607608
rect 330937 607550 489868 607552
rect 330937 607547 331003 607550
rect 489862 607548 489868 607550
rect 489932 607548 489938 607612
rect 293953 607474 294019 607477
rect 487838 607474 487844 607476
rect 293953 607472 487844 607474
rect 293953 607416 293958 607472
rect 294014 607416 487844 607472
rect 293953 607414 487844 607416
rect 293953 607411 294019 607414
rect 487838 607412 487844 607414
rect 487908 607412 487914 607476
rect 281441 607338 281507 607341
rect 491150 607338 491156 607340
rect 281441 607336 491156 607338
rect 281441 607280 281446 607336
rect 281502 607280 491156 607336
rect 281441 607278 491156 607280
rect 281441 607275 281507 607278
rect 491150 607276 491156 607278
rect 491220 607276 491226 607340
rect 428222 606658 428228 606660
rect 389222 606598 428228 606658
rect 389222 606522 389282 606598
rect 428222 606596 428228 606598
rect 428292 606596 428298 606660
rect 437790 606596 437796 606660
rect 437860 606658 437866 606660
rect 458766 606658 458772 606660
rect 437860 606598 458772 606658
rect 437860 606596 437866 606598
rect 458766 606596 458772 606598
rect 458836 606596 458842 606660
rect 380206 606462 389282 606522
rect 397729 606522 397795 606525
rect 500902 606522 500908 606524
rect 397729 606520 500908 606522
rect 397729 606464 397734 606520
rect 397790 606464 500908 606520
rect 397729 606462 500908 606464
rect 380206 606386 380266 606462
rect 397729 606459 397795 606462
rect 500902 606460 500908 606462
rect 500972 606460 500978 606524
rect 331262 606326 380266 606386
rect 385217 606386 385283 606389
rect 502374 606386 502380 606388
rect 385217 606384 502380 606386
rect 385217 606328 385222 606384
rect 385278 606328 502380 606384
rect 385217 606326 502380 606328
rect 235942 606188 235948 606252
rect 236012 606250 236018 606252
rect 244406 606250 244412 606252
rect 236012 606190 244412 606250
rect 236012 606188 236018 606190
rect 244406 606188 244412 606190
rect 244476 606188 244482 606252
rect 253974 606188 253980 606252
rect 254044 606250 254050 606252
rect 272926 606250 272932 606252
rect 254044 606190 272932 606250
rect 254044 606188 254050 606190
rect 272926 606188 272932 606190
rect 272996 606188 273002 606252
rect 273294 606188 273300 606252
rect 273364 606250 273370 606252
rect 331262 606250 331322 606326
rect 385217 606323 385283 606326
rect 502374 606324 502380 606326
rect 502444 606324 502450 606388
rect 273364 606190 331322 606250
rect 335905 606250 335971 606253
rect 507894 606250 507900 606252
rect 335905 606248 507900 606250
rect 335905 606192 335910 606248
rect 335966 606192 507900 606248
rect 335905 606190 507900 606192
rect 273364 606188 273370 606190
rect 335905 606187 335971 606190
rect 507894 606188 507900 606190
rect 507964 606188 507970 606252
rect 118918 606052 118924 606116
rect 118988 606114 118994 606116
rect 128670 606114 128676 606116
rect 118988 606054 128676 606114
rect 118988 606052 118994 606054
rect 128670 606052 128676 606054
rect 128740 606052 128746 606116
rect 138422 606052 138428 606116
rect 138492 606114 138498 606116
rect 157190 606114 157196 606116
rect 138492 606054 157196 606114
rect 138492 606052 138498 606054
rect 157190 606052 157196 606054
rect 157260 606052 157266 606116
rect 176878 606052 176884 606116
rect 176948 606114 176954 606116
rect 195830 606114 195836 606116
rect 176948 606054 195836 606114
rect 176948 606052 176954 606054
rect 195830 606052 195836 606054
rect 195900 606052 195906 606116
rect 196566 606052 196572 606116
rect 196636 606114 196642 606116
rect 207054 606114 207060 606116
rect 196636 606054 207060 606114
rect 196636 606052 196642 606054
rect 207054 606052 207060 606054
rect 207124 606052 207130 606116
rect 219801 606114 219867 606117
rect 499430 606114 499436 606116
rect 219801 606112 499436 606114
rect 219801 606056 219806 606112
rect 219862 606056 499436 606112
rect 219801 606054 499436 606056
rect 219801 606051 219867 606054
rect 499430 606052 499436 606054
rect 499500 606052 499506 606116
rect 93761 605978 93827 605981
rect 168281 605978 168347 605981
rect 93761 605976 168347 605978
rect 93761 605920 93766 605976
rect 93822 605920 168286 605976
rect 168342 605920 168347 605976
rect 93761 605918 168347 605920
rect 93761 605915 93827 605918
rect 168281 605915 168347 605918
rect 185209 605978 185275 605981
rect 516726 605978 516732 605980
rect 185209 605976 516732 605978
rect 185209 605920 185214 605976
rect 185270 605920 516732 605976
rect 185209 605918 516732 605920
rect 185209 605915 185275 605918
rect 516726 605916 516732 605918
rect 516796 605916 516802 605980
rect 89110 605508 89116 605572
rect 89180 605570 89186 605572
rect 90214 605570 90220 605572
rect 89180 605510 90220 605570
rect 89180 605508 89186 605510
rect 90214 605508 90220 605510
rect 90284 605508 90290 605572
rect 109718 605508 109724 605572
rect 109788 605570 109794 605572
rect 118550 605570 118556 605572
rect 109788 605510 118556 605570
rect 109788 605508 109794 605510
rect 118550 605508 118556 605510
rect 118620 605508 118626 605572
rect 157742 605508 157748 605572
rect 157812 605570 157818 605572
rect 176510 605570 176516 605572
rect 157812 605510 176516 605570
rect 157812 605508 157818 605510
rect 176510 605508 176516 605510
rect 176580 605508 176586 605572
rect 392761 605026 392827 605029
rect 492806 605026 492812 605028
rect 392761 605024 492812 605026
rect 392761 604968 392766 605024
rect 392822 604968 492812 605024
rect 392761 604966 492812 604968
rect 392761 604963 392827 604966
rect 492806 604964 492812 604966
rect 492876 604964 492882 605028
rect 67398 604828 67404 604892
rect 67468 604890 67474 604892
rect 190085 604890 190151 604893
rect 67468 604888 190151 604890
rect 67468 604832 190090 604888
rect 190146 604832 190151 604888
rect 67468 604830 190151 604832
rect 67468 604828 67474 604830
rect 190085 604827 190151 604830
rect 298737 604890 298803 604893
rect 491886 604890 491892 604892
rect 298737 604888 491892 604890
rect 298737 604832 298742 604888
rect 298798 604832 491892 604888
rect 298737 604830 491892 604832
rect 298737 604827 298803 604830
rect 491886 604828 491892 604830
rect 491956 604828 491962 604892
rect 157977 604754 158043 604757
rect 496854 604754 496860 604756
rect 157977 604752 496860 604754
rect 157977 604696 157982 604752
rect 158038 604696 496860 604752
rect 157977 604694 496860 604696
rect 157977 604691 158043 604694
rect 496854 604692 496860 604694
rect 496924 604692 496930 604756
rect 138289 604618 138355 604621
rect 558913 604618 558979 604621
rect 138289 604616 558979 604618
rect 138289 604560 138294 604616
rect 138350 604560 558918 604616
rect 558974 604560 558979 604616
rect 138289 604558 558979 604560
rect 138289 604555 138355 604558
rect 558913 604555 558979 604558
rect 103697 604482 103763 604485
rect 563697 604482 563763 604485
rect 103697 604480 563763 604482
rect 103697 604424 103702 604480
rect 103758 604424 563702 604480
rect 563758 604424 563763 604480
rect 103697 604422 563763 604424
rect 103697 604419 103763 604422
rect 563697 604419 563763 604422
rect 108430 604148 108436 604212
rect 108500 604210 108506 604212
rect 109718 604210 109724 604212
rect 108500 604150 109724 604210
rect 108500 604148 108506 604150
rect 109718 604148 109724 604150
rect 109788 604148 109794 604212
rect 147438 604148 147444 604212
rect 147508 604210 147514 604212
rect 157926 604210 157932 604212
rect 147508 604150 157932 604210
rect 147508 604148 147514 604150
rect 157926 604148 157932 604150
rect 157996 604148 158002 604212
rect 223614 604148 223620 604212
rect 223684 604210 223690 604212
rect 224902 604210 224908 604212
rect 223684 604150 224908 604210
rect 223684 604148 223690 604150
rect 224902 604148 224908 604150
rect 224972 604148 224978 604212
rect 263358 604148 263364 604212
rect 263428 604210 263434 604212
rect 264462 604210 264468 604212
rect 263428 604150 264468 604210
rect 263428 604148 263434 604150
rect 264462 604148 264468 604150
rect 264532 604148 264538 604212
rect 281206 604148 281212 604212
rect 281276 604210 281282 604212
rect 283046 604210 283052 604212
rect 281276 604150 283052 604210
rect 281276 604148 281282 604150
rect 283046 604148 283052 604150
rect 283116 604148 283122 604212
rect 378542 604148 378548 604212
rect 378612 604210 378618 604212
rect 389030 604210 389036 604212
rect 378612 604150 389036 604210
rect 378612 604148 378618 604150
rect 389030 604148 389036 604150
rect 389100 604148 389106 604212
rect 414422 604148 414428 604212
rect 414492 604210 414498 604212
rect 421598 604210 421604 604212
rect 414492 604150 421604 604210
rect 414492 604148 414498 604150
rect 421598 604148 421604 604150
rect 421668 604148 421674 604212
rect 437238 604148 437244 604212
rect 437308 604210 437314 604212
rect 439681 604210 439747 604213
rect 437308 604208 439747 604210
rect 437308 604152 439686 604208
rect 439742 604152 439747 604208
rect 437308 604150 439747 604152
rect 437308 604148 437314 604150
rect 439681 604147 439747 604150
rect 453982 604148 453988 604212
rect 454052 604210 454058 604212
rect 463601 604210 463667 604213
rect 583520 604210 584960 604300
rect 454052 604208 463667 604210
rect 454052 604152 463606 604208
rect 463662 604152 463667 604208
rect 454052 604150 463667 604152
rect 454052 604148 454058 604150
rect 463601 604147 463667 604150
rect 583342 604150 584960 604210
rect 67081 604074 67147 604077
rect 67081 604072 70594 604074
rect 67081 604016 67086 604072
rect 67142 604016 70594 604072
rect 67081 604014 70594 604016
rect 67081 604011 67147 604014
rect 70534 603938 70594 604014
rect 86902 604012 86908 604076
rect 86972 604074 86978 604076
rect 86972 604014 87338 604074
rect 86972 604012 86978 604014
rect 87278 603938 87338 604014
rect 99974 604014 109234 604074
rect 99974 603938 100034 604014
rect 70534 603878 75930 603938
rect 87278 603878 100034 603938
rect 75870 603836 75930 603878
rect 75870 603802 76114 603836
rect 86902 603802 86908 603804
rect 75870 603776 86908 603802
rect 76054 603742 86908 603776
rect 86902 603740 86908 603742
rect 86972 603740 86978 603804
rect 109174 603802 109234 604014
rect 153142 604012 153148 604076
rect 153212 604074 153218 604076
rect 196065 604074 196131 604077
rect 289813 604074 289879 604077
rect 309133 604074 309199 604077
rect 328453 604074 328519 604077
rect 347773 604074 347839 604077
rect 153212 604014 158178 604074
rect 153212 604012 153218 604014
rect 118785 603938 118851 603941
rect 138105 603938 138171 603941
rect 149605 603938 149671 603941
rect 118785 603936 129106 603938
rect 118785 603880 118790 603936
rect 118846 603880 129106 603936
rect 118785 603878 129106 603880
rect 118785 603875 118851 603878
rect 118601 603802 118667 603805
rect 109174 603800 118667 603802
rect 109174 603744 118606 603800
rect 118662 603744 118667 603800
rect 109174 603742 118667 603744
rect 129046 603802 129106 603878
rect 138105 603936 149671 603938
rect 138105 603880 138110 603936
rect 138166 603880 149610 603936
rect 149666 603880 149671 603936
rect 138105 603878 149671 603880
rect 158118 603938 158178 604014
rect 172286 604014 186514 604074
rect 172286 603938 172346 604014
rect 158118 603878 172346 603938
rect 138105 603875 138171 603878
rect 149605 603875 149671 603878
rect 137921 603802 137987 603805
rect 129046 603800 137987 603802
rect 129046 603744 137926 603800
rect 137982 603744 137987 603800
rect 129046 603742 137987 603744
rect 118601 603739 118667 603742
rect 137921 603739 137987 603742
rect 149697 603802 149763 603805
rect 153142 603802 153148 603804
rect 149697 603800 153148 603802
rect 149697 603744 149702 603800
rect 149758 603744 153148 603800
rect 149697 603742 153148 603744
rect 149697 603739 149763 603742
rect 153142 603740 153148 603742
rect 153212 603740 153218 603804
rect 186454 603802 186514 604014
rect 196065 604072 205834 604074
rect 196065 604016 196070 604072
rect 196126 604016 205834 604072
rect 196065 604014 205834 604016
rect 196065 604011 196131 604014
rect 195881 603802 195947 603805
rect 186454 603800 195947 603802
rect 186454 603744 195886 603800
rect 195942 603744 195947 603800
rect 186454 603742 195947 603744
rect 205774 603802 205834 604014
rect 215158 604014 225154 604074
rect 215158 603802 215218 604014
rect 205774 603742 215218 603802
rect 225094 603802 225154 604014
rect 234478 604014 244474 604074
rect 234478 603802 234538 604014
rect 225094 603742 234538 603802
rect 244414 603802 244474 604014
rect 253798 604014 263794 604074
rect 253798 603802 253858 604014
rect 244414 603742 253858 603802
rect 263734 603802 263794 604014
rect 282870 604072 289879 604074
rect 282870 604016 289818 604072
rect 289874 604016 289879 604072
rect 282870 604014 289879 604016
rect 282870 603802 282930 604014
rect 289813 604011 289879 604014
rect 302190 604072 309199 604074
rect 302190 604016 309138 604072
rect 309194 604016 309199 604072
rect 302190 604014 309199 604016
rect 263734 603742 282930 603802
rect 299381 603802 299447 603805
rect 302190 603802 302250 604014
rect 309133 604011 309199 604014
rect 321510 604072 328519 604074
rect 321510 604016 328458 604072
rect 328514 604016 328519 604072
rect 321510 604014 328519 604016
rect 299381 603800 302250 603802
rect 299381 603744 299386 603800
rect 299442 603744 302250 603800
rect 299381 603742 302250 603744
rect 318701 603802 318767 603805
rect 321510 603802 321570 604014
rect 328453 604011 328519 604014
rect 340830 604072 347839 604074
rect 340830 604016 347778 604072
rect 347834 604016 347839 604072
rect 340830 604014 347839 604016
rect 318701 603800 321570 603802
rect 318701 603744 318706 603800
rect 318762 603744 321570 603800
rect 318701 603742 321570 603744
rect 338021 603802 338087 603805
rect 340830 603802 340890 604014
rect 347773 604011 347839 604014
rect 488574 604012 488580 604076
rect 488644 604074 488650 604076
rect 488993 604074 489059 604077
rect 488644 604072 489059 604074
rect 488644 604016 488998 604072
rect 489054 604016 489059 604072
rect 488644 604014 489059 604016
rect 488644 604012 488650 604014
rect 488993 604011 489059 604014
rect 553350 604014 563162 604074
rect 357341 603938 357407 603941
rect 357341 603936 360210 603938
rect 357341 603880 357346 603936
rect 357402 603880 360210 603936
rect 357341 603878 360210 603880
rect 357341 603875 357407 603878
rect 338021 603800 340890 603802
rect 338021 603744 338026 603800
rect 338082 603744 340890 603800
rect 338021 603742 340890 603744
rect 360150 603802 360210 603878
rect 384982 603876 384988 603940
rect 385052 603938 385058 603940
rect 463601 603938 463667 603941
rect 483013 603938 483079 603941
rect 385052 603878 399034 603938
rect 385052 603876 385058 603878
rect 369669 603802 369735 603805
rect 360150 603800 369735 603802
rect 360150 603744 369674 603800
rect 369730 603744 369735 603800
rect 360150 603742 369735 603744
rect 195881 603739 195947 603742
rect 299381 603739 299447 603742
rect 318701 603739 318767 603742
rect 338021 603739 338087 603742
rect 369669 603739 369735 603742
rect 369945 603802 370011 603805
rect 379421 603802 379487 603805
rect 369945 603800 379487 603802
rect 369945 603744 369950 603800
rect 370006 603744 379426 603800
rect 379482 603744 379487 603800
rect 369945 603742 379487 603744
rect 369945 603739 370011 603742
rect 379421 603739 379487 603742
rect 70894 603604 70900 603668
rect 70964 603666 70970 603668
rect 350625 603666 350691 603669
rect 70964 603664 350691 603666
rect 70964 603608 350630 603664
rect 350686 603608 350691 603664
rect 70964 603606 350691 603608
rect 70964 603604 70970 603606
rect 350625 603603 350691 603606
rect 379605 603666 379671 603669
rect 384982 603666 384988 603668
rect 379605 603664 384988 603666
rect 379605 603608 379610 603664
rect 379666 603608 384988 603664
rect 379605 603606 384988 603608
rect 379605 603603 379671 603606
rect 384982 603604 384988 603606
rect 385052 603604 385058 603668
rect 398974 603666 399034 603878
rect 404494 603878 437674 603938
rect 404494 603802 404554 603878
rect 404310 603742 404554 603802
rect 404310 603666 404370 603742
rect 398974 603606 404370 603666
rect 437614 603666 437674 603878
rect 463601 603936 466194 603938
rect 463601 603880 463606 603936
rect 463662 603880 466194 603936
rect 463601 603878 466194 603880
rect 463601 603875 463667 603878
rect 449157 603802 449223 603805
rect 453982 603802 453988 603804
rect 449157 603800 453988 603802
rect 449157 603744 449162 603800
rect 449218 603744 453988 603800
rect 449157 603742 453988 603744
rect 449157 603739 449223 603742
rect 453982 603740 453988 603742
rect 454052 603740 454058 603804
rect 466134 603802 466194 603878
rect 476254 603936 483079 603938
rect 476254 603880 483018 603936
rect 483074 603880 483079 603936
rect 476254 603878 483079 603880
rect 473261 603802 473327 603805
rect 476254 603802 476314 603878
rect 483013 603875 483079 603878
rect 492765 603938 492831 603941
rect 516869 603938 516935 603941
rect 492765 603936 516935 603938
rect 492765 603880 492770 603936
rect 492826 603880 516874 603936
rect 516930 603880 516935 603936
rect 492765 603878 516935 603880
rect 492765 603875 492831 603878
rect 516869 603875 516935 603878
rect 466134 603800 473327 603802
rect 466134 603744 473266 603800
rect 473322 603744 473327 603800
rect 466134 603742 473327 603744
rect 473261 603739 473327 603742
rect 476070 603742 476314 603802
rect 540881 603802 540947 603805
rect 553350 603802 553410 604014
rect 540881 603800 553410 603802
rect 540881 603744 540886 603800
rect 540942 603744 553410 603800
rect 540881 603742 553410 603744
rect 563102 603802 563162 604014
rect 583342 603938 583402 604150
rect 583520 604060 584960 604150
rect 582238 603878 583402 603938
rect 572621 603802 572687 603805
rect 563102 603800 572687 603802
rect 563102 603744 572626 603800
rect 572682 603744 572687 603800
rect 563102 603742 572687 603744
rect 444373 603666 444439 603669
rect 437614 603664 444439 603666
rect 437614 603608 444378 603664
rect 444434 603608 444439 603664
rect 437614 603606 444439 603608
rect 444373 603603 444439 603606
rect 473261 603666 473327 603669
rect 476070 603666 476130 603742
rect 540881 603739 540947 603742
rect 572621 603739 572687 603742
rect 572805 603802 572871 603805
rect 582238 603802 582298 603878
rect 572805 603800 582298 603802
rect 572805 603744 572810 603800
rect 572866 603744 582298 603800
rect 572805 603742 582298 603744
rect 572805 603739 572871 603742
rect 473261 603664 476130 603666
rect 473261 603608 473266 603664
rect 473322 603608 476130 603664
rect 473261 603606 476130 603608
rect 525701 603666 525767 603669
rect 533981 603666 534047 603669
rect 525701 603664 534047 603666
rect 525701 603608 525706 603664
rect 525762 603608 533986 603664
rect 534042 603608 534047 603664
rect 525701 603606 534047 603608
rect 473261 603603 473327 603606
rect 525701 603603 525767 603606
rect 533981 603603 534047 603606
rect 89662 603468 89668 603532
rect 89732 603530 89738 603532
rect 170305 603530 170371 603533
rect 89732 603528 170371 603530
rect 89732 603472 170310 603528
rect 170366 603472 170371 603528
rect 89732 603470 170371 603472
rect 89732 603468 89738 603470
rect 170305 603467 170371 603470
rect 212257 603530 212323 603533
rect 516133 603530 516199 603533
rect 212257 603528 516199 603530
rect 212257 603472 212262 603528
rect 212318 603472 516138 603528
rect 516194 603472 516199 603528
rect 212257 603470 516199 603472
rect 212257 603467 212323 603470
rect 516133 603467 516199 603470
rect 72366 603332 72372 603396
rect 72436 603394 72442 603396
rect 429745 603394 429811 603397
rect 72436 603392 429811 603394
rect 72436 603336 429750 603392
rect 429806 603336 429811 603392
rect 72436 603334 429811 603336
rect 72436 603332 72442 603334
rect 429745 603331 429811 603334
rect 442073 603394 442139 603397
rect 485998 603394 486004 603396
rect 442073 603392 486004 603394
rect 442073 603336 442078 603392
rect 442134 603336 486004 603392
rect 442073 603334 486004 603336
rect 442073 603331 442139 603334
rect 485998 603332 486004 603334
rect 486068 603332 486074 603396
rect 491569 603394 491635 603397
rect 517881 603394 517947 603397
rect 491569 603392 517947 603394
rect 491569 603336 491574 603392
rect 491630 603336 517886 603392
rect 517942 603336 517947 603392
rect 491569 603334 517947 603336
rect 491569 603331 491635 603334
rect 517881 603331 517947 603334
rect 82854 603196 82860 603260
rect 82924 603258 82930 603260
rect 447041 603258 447107 603261
rect 82924 603256 447107 603258
rect 82924 603200 447046 603256
rect 447102 603200 447107 603256
rect 82924 603198 447107 603200
rect 82924 603196 82930 603198
rect 447041 603195 447107 603198
rect 449617 603258 449683 603261
rect 510705 603258 510771 603261
rect 449617 603256 510771 603258
rect 449617 603200 449622 603256
rect 449678 603200 510710 603256
rect 510766 603200 510771 603256
rect 449617 603198 510771 603200
rect 449617 603195 449683 603198
rect 510705 603195 510771 603198
rect 495934 603060 495940 603124
rect 496004 603122 496010 603124
rect 498929 603122 498995 603125
rect 496004 603120 498995 603122
rect 496004 603064 498934 603120
rect 498990 603064 498995 603120
rect 496004 603062 498995 603064
rect 496004 603060 496010 603062
rect 498929 603059 498995 603062
rect 496854 602924 496860 602988
rect 496924 602924 496930 602988
rect 496862 602850 496922 602924
rect 497222 602850 497228 602852
rect 496862 602790 497228 602850
rect 497222 602788 497228 602790
rect 497292 602788 497298 602852
rect 346393 602442 346459 602445
rect 482870 602442 482876 602444
rect 346393 602440 482876 602442
rect 346393 602384 346398 602440
rect 346454 602384 482876 602440
rect 346393 602382 482876 602384
rect 346393 602379 346459 602382
rect 482870 602380 482876 602382
rect 482940 602380 482946 602444
rect 60641 602306 60707 602309
rect 88333 602306 88399 602309
rect 60641 602304 88399 602306
rect 60641 602248 60646 602304
rect 60702 602248 88338 602304
rect 88394 602248 88399 602304
rect 60641 602246 88399 602248
rect 60641 602243 60707 602246
rect 88333 602243 88399 602246
rect 318793 602306 318859 602309
rect 492622 602306 492628 602308
rect 318793 602304 492628 602306
rect 318793 602248 318798 602304
rect 318854 602248 492628 602304
rect 318793 602246 492628 602248
rect 318793 602243 318859 602246
rect 492622 602244 492628 602246
rect 492692 602244 492698 602308
rect 72550 602108 72556 602172
rect 72620 602170 72626 602172
rect 286409 602170 286475 602173
rect 72620 602168 286475 602170
rect 72620 602112 286414 602168
rect 286470 602112 286475 602168
rect 72620 602110 286475 602112
rect 72620 602108 72626 602110
rect 286409 602107 286475 602110
rect 288985 602170 289051 602173
rect 488574 602170 488580 602172
rect 288985 602168 488580 602170
rect 288985 602112 288990 602168
rect 289046 602112 488580 602168
rect 288985 602110 488580 602112
rect 288985 602107 289051 602110
rect 488574 602108 488580 602110
rect 488644 602108 488650 602172
rect 75126 601972 75132 602036
rect 75196 602034 75202 602036
rect 315941 602034 316007 602037
rect 75196 602032 316007 602034
rect 75196 601976 315946 602032
rect 316002 601976 316007 602032
rect 75196 601974 316007 601976
rect 75196 601972 75202 601974
rect 315941 601971 316007 601974
rect 481817 602034 481883 602037
rect 520273 602034 520339 602037
rect 481817 602032 520339 602034
rect 481817 601976 481822 602032
rect 481878 601976 520278 602032
rect 520334 601976 520339 602032
rect 481817 601974 520339 601976
rect 481817 601971 481883 601974
rect 520273 601971 520339 601974
rect 48221 601898 48287 601901
rect 104893 601898 104959 601901
rect 48221 601896 104959 601898
rect 48221 601840 48226 601896
rect 48282 601840 104898 601896
rect 104954 601840 104959 601896
rect 48221 601838 104959 601840
rect 48221 601835 48287 601838
rect 104893 601835 104959 601838
rect 267089 601898 267155 601901
rect 517513 601898 517579 601901
rect 267089 601896 517579 601898
rect 267089 601840 267094 601896
rect 267150 601840 517518 601896
rect 517574 601840 517579 601896
rect 267089 601838 517579 601840
rect 267089 601835 267155 601838
rect 517513 601835 517579 601838
rect 52361 601762 52427 601765
rect 367645 601762 367711 601765
rect 52361 601760 367711 601762
rect 52361 601704 52366 601760
rect 52422 601704 367650 601760
rect 367706 601704 367711 601760
rect 52361 601702 367711 601704
rect 52361 601699 52427 601702
rect 367645 601699 367711 601702
rect 427721 601762 427787 601765
rect 501638 601762 501644 601764
rect 427721 601760 501644 601762
rect 427721 601704 427726 601760
rect 427782 601704 501644 601760
rect 427721 601702 501644 601704
rect 427721 601699 427787 601702
rect 501638 601700 501644 601702
rect 501708 601700 501714 601764
rect 75862 601292 75868 601356
rect 75932 601354 75938 601356
rect 80697 601354 80763 601357
rect 75932 601352 80763 601354
rect 75932 601296 80702 601352
rect 80758 601296 80763 601352
rect 75932 601294 80763 601296
rect 75932 601292 75938 601294
rect 80697 601291 80763 601294
rect 83365 601354 83431 601357
rect 92381 601354 92447 601357
rect 83365 601352 92447 601354
rect 83365 601296 83370 601352
rect 83426 601296 92386 601352
rect 92442 601296 92447 601352
rect 83365 601294 92447 601296
rect 83365 601291 83431 601294
rect 92381 601291 92447 601294
rect 162853 601356 162919 601357
rect 162853 601352 162900 601356
rect 162964 601354 162970 601356
rect 195329 601354 195395 601357
rect 200614 601354 200620 601356
rect 162853 601296 162858 601352
rect 162853 601292 162900 601296
rect 162964 601294 163010 601354
rect 195329 601352 200620 601354
rect 195329 601296 195334 601352
rect 195390 601296 200620 601352
rect 195329 601294 200620 601296
rect 162964 601292 162970 601294
rect 162853 601291 162919 601292
rect 195329 601291 195395 601294
rect 200614 601292 200620 601294
rect 200684 601292 200690 601356
rect 200798 601292 200804 601356
rect 200868 601354 200874 601356
rect 207197 601354 207263 601357
rect 200868 601352 207263 601354
rect 200868 601296 207202 601352
rect 207258 601296 207263 601352
rect 200868 601294 207263 601296
rect 200868 601292 200874 601294
rect 207197 601291 207263 601294
rect 249701 601354 249767 601357
rect 258758 601354 258764 601356
rect 249701 601352 258764 601354
rect 249701 601296 249706 601352
rect 249762 601296 258764 601352
rect 249701 601294 258764 601296
rect 249701 601291 249767 601294
rect 258758 601292 258764 601294
rect 258828 601292 258834 601356
rect 260782 601292 260788 601356
rect 260852 601354 260858 601356
rect 270350 601354 270356 601356
rect 260852 601294 270356 601354
rect 260852 601292 260858 601294
rect 270350 601292 270356 601294
rect 270420 601292 270426 601356
rect 270534 601292 270540 601356
rect 270604 601354 270610 601356
rect 278773 601354 278839 601357
rect 296069 601354 296135 601357
rect 270604 601352 278839 601354
rect 270604 601296 278778 601352
rect 278834 601296 278839 601352
rect 270604 601294 278839 601296
rect 270604 601292 270610 601294
rect 278773 601291 278839 601294
rect 291702 601352 296135 601354
rect 291702 601296 296074 601352
rect 296130 601296 296135 601352
rect 291702 601294 296135 601296
rect 86902 601156 86908 601220
rect 86972 601218 86978 601220
rect 86972 601158 87154 601218
rect 86972 601156 86978 601158
rect 59169 601082 59235 601085
rect 75862 601082 75868 601084
rect 59169 601080 75868 601082
rect 59169 601024 59174 601080
rect 59230 601024 75868 601080
rect 59169 601022 75868 601024
rect 59169 601019 59235 601022
rect 75862 601020 75868 601022
rect 75932 601020 75938 601084
rect 87094 601082 87154 601158
rect 135110 601156 135116 601220
rect 135180 601218 135186 601220
rect 135180 601158 135362 601218
rect 135180 601156 135186 601158
rect 87094 601022 113098 601082
rect 80697 600946 80763 600949
rect 86902 600946 86908 600948
rect 80697 600944 86908 600946
rect 80697 600888 80702 600944
rect 80758 600888 86908 600944
rect 80697 600886 86908 600888
rect 80697 600883 80763 600886
rect 86902 600884 86908 600886
rect 86972 600884 86978 600948
rect 113038 600946 113098 601022
rect 124254 601020 124260 601084
rect 124324 601082 124330 601084
rect 135302 601082 135362 601158
rect 153142 601156 153148 601220
rect 153212 601218 153218 601220
rect 153212 601158 158178 601218
rect 153212 601156 153218 601158
rect 158118 601082 158178 601158
rect 167678 601156 167684 601220
rect 167748 601218 167754 601220
rect 172278 601218 172284 601220
rect 167748 601158 172284 601218
rect 167748 601156 167754 601158
rect 172278 601156 172284 601158
rect 172348 601156 172354 601220
rect 175966 601158 176762 601218
rect 175966 601082 176026 601158
rect 124324 601022 132418 601082
rect 135302 601022 149714 601082
rect 158118 601022 176026 601082
rect 176702 601082 176762 601158
rect 176702 601022 188170 601082
rect 124324 601020 124330 601022
rect 124070 600946 124076 600948
rect 113038 600886 124076 600946
rect 124070 600884 124076 600886
rect 124140 600884 124146 600948
rect 132358 600946 132418 601022
rect 135110 600946 135116 600948
rect 132358 600886 135116 600946
rect 135110 600884 135116 600886
rect 135180 600884 135186 600948
rect 149654 600946 149714 601022
rect 153142 600946 153148 600948
rect 149654 600886 153148 600946
rect 153142 600884 153148 600886
rect 153212 600884 153218 600948
rect 172278 600884 172284 600948
rect 172348 600884 172354 600948
rect 188110 600946 188170 601022
rect 205590 601022 205834 601082
rect 195830 600946 195836 600948
rect 188110 600886 195836 600946
rect 195830 600884 195836 600886
rect 195900 600884 195906 600948
rect 202822 600884 202828 600948
rect 202892 600946 202898 600948
rect 205590 600946 205650 601022
rect 202892 600886 205650 600946
rect 205774 600946 205834 601022
rect 215334 601020 215340 601084
rect 215404 601082 215410 601084
rect 215404 601022 226994 601082
rect 215404 601020 215410 601022
rect 215150 600946 215156 600948
rect 205774 600886 215156 600946
rect 202892 600884 202898 600886
rect 215150 600884 215156 600886
rect 215220 600884 215226 600948
rect 226934 600946 226994 601022
rect 234654 601020 234660 601084
rect 234724 601082 234730 601084
rect 234724 601022 246314 601082
rect 234724 601020 234730 601022
rect 234470 600946 234476 600948
rect 226934 600886 234476 600946
rect 234470 600884 234476 600886
rect 234540 600884 234546 600948
rect 246254 600946 246314 601022
rect 253974 601020 253980 601084
rect 254044 601082 254050 601084
rect 260782 601082 260788 601084
rect 254044 601022 260788 601082
rect 254044 601020 254050 601022
rect 260782 601020 260788 601022
rect 260852 601020 260858 601084
rect 270350 601020 270356 601084
rect 270420 601020 270426 601084
rect 253790 600946 253796 600948
rect 246254 600886 253796 600946
rect 253790 600884 253796 600886
rect 253860 600884 253866 600948
rect 270358 600946 270418 601020
rect 270534 600946 270540 600948
rect 270358 600886 270540 600946
rect 270534 600884 270540 600886
rect 270604 600884 270610 600948
rect 74165 600810 74231 600813
rect 167678 600810 167684 600812
rect 74165 600808 167684 600810
rect 74165 600752 74170 600808
rect 74226 600752 167684 600808
rect 74165 600750 167684 600752
rect 74165 600747 74231 600750
rect 167678 600748 167684 600750
rect 167748 600748 167754 600812
rect 172286 600810 172346 600884
rect 291702 600810 291762 601294
rect 296069 601291 296135 601294
rect 301446 601292 301452 601356
rect 301516 601354 301522 601356
rect 306005 601354 306071 601357
rect 301516 601352 306071 601354
rect 301516 601296 306010 601352
rect 306066 601296 306071 601352
rect 301516 601294 306071 601296
rect 301516 601292 301522 601294
rect 306005 601291 306071 601294
rect 402881 601354 402947 601357
rect 405038 601354 405044 601356
rect 402881 601352 405044 601354
rect 402881 601296 402886 601352
rect 402942 601296 405044 601352
rect 402881 601294 405044 601296
rect 402881 601291 402947 601294
rect 405038 601292 405044 601294
rect 405108 601292 405114 601356
rect 405457 601354 405523 601357
rect 409086 601354 409092 601356
rect 405457 601352 409092 601354
rect 405457 601296 405462 601352
rect 405518 601296 409092 601352
rect 405457 601294 409092 601296
rect 405457 601291 405523 601294
rect 409086 601292 409092 601294
rect 409156 601292 409162 601356
rect 415393 601354 415459 601357
rect 435081 601354 435147 601357
rect 476941 601356 477007 601357
rect 415393 601352 415962 601354
rect 415393 601296 415398 601352
rect 415454 601296 415962 601352
rect 415393 601294 415962 601296
rect 415393 601291 415459 601294
rect 172286 600750 291762 600810
rect 415902 600810 415962 601294
rect 435081 601352 436202 601354
rect 435081 601296 435086 601352
rect 435142 601296 436202 601352
rect 435081 601294 436202 601296
rect 435081 601291 435147 601294
rect 436142 600946 436202 601294
rect 476941 601352 476988 601356
rect 477052 601354 477058 601356
rect 476941 601296 476946 601352
rect 476941 601292 476988 601296
rect 477052 601294 477098 601354
rect 477052 601292 477058 601294
rect 486182 601292 486188 601356
rect 486252 601354 486258 601356
rect 486325 601354 486391 601357
rect 486252 601352 486391 601354
rect 486252 601296 486330 601352
rect 486386 601296 486391 601352
rect 486252 601294 486391 601296
rect 486252 601292 486258 601294
rect 476941 601291 477007 601292
rect 486325 601291 486391 601294
rect 494830 601292 494836 601356
rect 494900 601354 494906 601356
rect 496261 601354 496327 601357
rect 494900 601352 496327 601354
rect 494900 601296 496266 601352
rect 496322 601296 496327 601352
rect 494900 601294 496327 601296
rect 494900 601292 494906 601294
rect 496261 601291 496327 601294
rect 497590 600946 497596 600948
rect 436142 600886 497596 600946
rect 497590 600884 497596 600886
rect 497660 600884 497666 600948
rect 498326 600810 498332 600812
rect 415902 600750 498332 600810
rect 498326 600748 498332 600750
rect 498396 600748 498402 600812
rect 24669 600674 24735 600677
rect 167678 600674 167684 600676
rect 24669 600672 167684 600674
rect 24669 600616 24674 600672
rect 24730 600616 167684 600672
rect 24669 600614 167684 600616
rect 24669 600611 24735 600614
rect 167678 600612 167684 600614
rect 167748 600612 167754 600676
rect 172278 600612 172284 600676
rect 172348 600674 172354 600676
rect 200798 600674 200804 600676
rect 172348 600614 200804 600674
rect 172348 600612 172354 600614
rect 200798 600612 200804 600614
rect 200868 600612 200874 600676
rect 258758 600612 258764 600676
rect 258828 600674 258834 600676
rect 495382 600674 495388 600676
rect 258828 600614 495388 600674
rect 258828 600612 258834 600614
rect 495382 600612 495388 600614
rect 495452 600612 495458 600676
rect 13077 600538 13143 600541
rect 301446 600538 301452 600540
rect 13077 600536 301452 600538
rect 13077 600480 13082 600536
rect 13138 600480 301452 600536
rect 13077 600478 301452 600480
rect 13077 600475 13143 600478
rect 301446 600476 301452 600478
rect 301516 600476 301522 600540
rect 409086 600476 409092 600540
rect 409156 600538 409162 600540
rect 494278 600538 494284 600540
rect 409156 600478 494284 600538
rect 409156 600476 409162 600478
rect 494278 600476 494284 600478
rect 494348 600476 494354 600540
rect 53741 600402 53807 600405
rect 83365 600402 83431 600405
rect 53741 600400 83431 600402
rect 53741 600344 53746 600400
rect 53802 600344 83370 600400
rect 83426 600344 83431 600400
rect 53741 600342 83431 600344
rect 53741 600339 53807 600342
rect 83365 600339 83431 600342
rect 200614 600340 200620 600404
rect 200684 600402 200690 600404
rect 511206 600402 511212 600404
rect 200684 600342 511212 600402
rect 200684 600340 200690 600342
rect 511206 600340 511212 600342
rect 511276 600340 511282 600404
rect 82854 600266 82860 600268
rect 80654 600206 82860 600266
rect 75678 600068 75684 600132
rect 75748 600130 75754 600132
rect 80654 600130 80714 600206
rect 82854 600204 82860 600206
rect 82924 600204 82930 600268
rect 167678 600204 167684 600268
rect 167748 600266 167754 600268
rect 172278 600266 172284 600268
rect 167748 600206 172284 600266
rect 167748 600204 167754 600206
rect 172278 600204 172284 600206
rect 172348 600204 172354 600268
rect 195830 600204 195836 600268
rect 195900 600266 195906 600268
rect 202638 600266 202644 600268
rect 195900 600206 202644 600266
rect 195900 600204 195906 600206
rect 202638 600204 202644 600206
rect 202708 600204 202714 600268
rect 499798 600204 499804 600268
rect 499868 600266 499874 600268
rect 501505 600266 501571 600269
rect 499868 600264 501571 600266
rect 499868 600208 501510 600264
rect 501566 600208 501571 600264
rect 499868 600206 501571 600208
rect 499868 600204 499874 600206
rect 501505 600203 501571 600206
rect 75748 600070 80714 600130
rect 75748 600068 75754 600070
rect 80830 600068 80836 600132
rect 80900 600130 80906 600132
rect 89662 600130 89668 600132
rect 80900 600070 89668 600130
rect 80900 600068 80906 600070
rect 89662 600068 89668 600070
rect 89732 600068 89738 600132
rect 487838 600068 487844 600132
rect 487908 600130 487914 600132
rect 488206 600130 488212 600132
rect 487908 600070 488212 600130
rect 487908 600068 487914 600070
rect 488206 600068 488212 600070
rect 488276 600068 488282 600132
rect 71405 599994 71471 599997
rect 162894 599994 162900 599996
rect 71405 599992 162900 599994
rect 71405 599936 71410 599992
rect 71466 599936 162900 599992
rect 71405 599934 162900 599936
rect 71405 599931 71471 599934
rect 162894 599932 162900 599934
rect 162964 599932 162970 599996
rect 405038 599932 405044 599996
rect 405108 599932 405114 599996
rect 482870 599932 482876 599996
rect 482940 599994 482946 599996
rect 489862 599994 489868 599996
rect 482940 599934 489868 599994
rect 482940 599932 482946 599934
rect 489862 599932 489868 599934
rect 489932 599932 489938 599996
rect 491150 599932 491156 599996
rect 491220 599994 491226 599996
rect 493174 599994 493180 599996
rect 491220 599934 493180 599994
rect 491220 599932 491226 599934
rect 493174 599932 493180 599934
rect 493244 599932 493250 599996
rect 78673 599586 78739 599589
rect 78673 599584 82156 599586
rect 78673 599528 78678 599584
rect 78734 599528 82156 599584
rect 78673 599526 82156 599528
rect 78673 599523 78739 599526
rect 405046 599452 405106 599932
rect 405038 599388 405044 599452
rect 405108 599388 405114 599452
rect 511574 598028 511580 598092
rect 511644 598090 511650 598092
rect 515254 598090 515260 598092
rect 511644 598030 515260 598090
rect 511644 598028 511650 598030
rect 515254 598028 515260 598030
rect 515324 598028 515330 598092
rect 501646 596594 501706 597380
rect 501646 596534 501890 596594
rect 501830 596322 501890 596534
rect 513414 596322 513420 596324
rect 501830 596262 513420 596322
rect 513414 596260 513420 596262
rect 513484 596260 513490 596324
rect -960 596050 480 596140
rect 2865 596050 2931 596053
rect -960 596048 2931 596050
rect -960 595992 2870 596048
rect 2926 595992 2931 596048
rect -960 595990 2931 595992
rect -960 595900 480 595990
rect 2865 595987 2931 595990
rect 78673 595778 78739 595781
rect 78673 595776 82156 595778
rect 78673 595720 78678 595776
rect 78734 595720 82156 595776
rect 78673 595718 82156 595720
rect 78673 595715 78739 595718
rect 35801 595506 35867 595509
rect 82486 595506 82492 595508
rect 35801 595504 82492 595506
rect 35801 595448 35806 595504
rect 35862 595448 82492 595504
rect 35801 595446 82492 595448
rect 35801 595443 35867 595446
rect 82486 595444 82492 595446
rect 82556 595444 82562 595508
rect 503897 593874 503963 593877
rect 501860 593872 503963 593874
rect 501860 593816 503902 593872
rect 503958 593816 503963 593872
rect 501860 593814 503963 593816
rect 503897 593811 503963 593814
rect 579889 592514 579955 592517
rect 583520 592514 584960 592604
rect 579889 592512 584960 592514
rect 579889 592456 579894 592512
rect 579950 592456 584960 592512
rect 579889 592454 584960 592456
rect 579889 592451 579955 592454
rect 583520 592364 584960 592454
rect 78673 592242 78739 592245
rect 78673 592240 82156 592242
rect 78673 592184 78678 592240
rect 78734 592184 82156 592240
rect 78673 592182 82156 592184
rect 78673 592179 78739 592182
rect 522062 592106 522068 592108
rect 521886 592046 522068 592106
rect 521886 591836 521946 592046
rect 522062 592044 522068 592046
rect 522132 592044 522138 592108
rect 521878 591772 521884 591836
rect 521948 591772 521954 591836
rect 501462 589525 501522 590036
rect 501462 589520 501571 589525
rect 501462 589464 501510 589520
rect 501566 589464 501571 589520
rect 501462 589462 501571 589464
rect 501505 589459 501571 589462
rect 501638 589324 501644 589388
rect 501708 589324 501714 589388
rect 501646 589114 501706 589324
rect 501822 589114 501828 589116
rect 501646 589054 501828 589114
rect 501822 589052 501828 589054
rect 501892 589052 501898 589116
rect 78438 588372 78444 588436
rect 78508 588434 78514 588436
rect 78508 588374 82156 588434
rect 78508 588372 78514 588374
rect 503897 586530 503963 586533
rect 501860 586528 503963 586530
rect 501860 586472 503902 586528
rect 503958 586472 503963 586528
rect 501860 586470 503963 586472
rect 503897 586467 503963 586470
rect 503897 582722 503963 582725
rect 501860 582720 503963 582722
rect 501860 582664 503902 582720
rect 503958 582664 503963 582720
rect 501860 582662 503963 582664
rect 503897 582659 503963 582662
rect 66846 582388 66852 582452
rect 66916 582388 66922 582452
rect 521878 582388 521884 582452
rect 521948 582388 521954 582452
rect 66854 582178 66914 582388
rect 67030 582178 67036 582180
rect 66854 582118 67036 582178
rect 67030 582116 67036 582118
rect 67100 582116 67106 582180
rect 521886 582178 521946 582388
rect 522062 582178 522068 582180
rect 521886 582118 522068 582178
rect 522062 582116 522068 582118
rect 522132 582116 522138 582180
rect -960 581620 480 581860
rect 81382 581300 81388 581364
rect 81452 581362 81458 581364
rect 81452 581302 82156 581362
rect 81452 581300 81458 581302
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 501638 579668 501644 579732
rect 501708 579668 501714 579732
rect 501646 579596 501706 579668
rect 501638 579532 501644 579596
rect 501708 579532 501714 579596
rect 521929 579594 521995 579597
rect 522062 579594 522068 579596
rect 521929 579592 522068 579594
rect 521929 579536 521934 579592
rect 521990 579536 522068 579592
rect 521929 579534 522068 579536
rect 521929 579531 521995 579534
rect 522062 579532 522068 579534
rect 522132 579532 522138 579596
rect 505502 579186 505508 579188
rect 501860 579126 505508 579186
rect 505502 579124 505508 579126
rect 505572 579124 505578 579188
rect 66989 578236 67055 578237
rect 66989 578234 67036 578236
rect 66944 578232 67036 578234
rect 66944 578176 66994 578232
rect 66944 578174 67036 578176
rect 66989 578172 67036 578174
rect 67100 578172 67106 578236
rect 66989 578171 67055 578172
rect 78949 577554 79015 577557
rect 78949 577552 82156 577554
rect 78949 577496 78954 577552
rect 79010 577496 82156 577552
rect 78949 577494 82156 577496
rect 78949 577491 79015 577494
rect 504449 575650 504515 575653
rect 501860 575648 504515 575650
rect 501860 575592 504454 575648
rect 504510 575592 504515 575648
rect 501860 575590 504515 575592
rect 504449 575587 504515 575590
rect 78765 574018 78831 574021
rect 78765 574016 82156 574018
rect 78765 573960 78770 574016
rect 78826 573960 82156 574016
rect 78765 573958 82156 573960
rect 78765 573955 78831 573958
rect 66989 572660 67055 572661
rect 66989 572656 67036 572660
rect 67100 572658 67106 572660
rect 66989 572600 66994 572656
rect 66989 572596 67036 572600
rect 67100 572598 67146 572658
rect 67100 572596 67106 572598
rect 66989 572595 67055 572596
rect 503897 571842 503963 571845
rect 501860 571840 503963 571842
rect 501860 571784 503902 571840
rect 503958 571784 503963 571840
rect 501860 571782 503963 571784
rect 503897 571779 503963 571782
rect 78673 570210 78739 570213
rect 512821 570210 512887 570213
rect 521929 570210 521995 570213
rect 78673 570208 82156 570210
rect 78673 570152 78678 570208
rect 78734 570152 82156 570208
rect 78673 570150 82156 570152
rect 512686 570208 512887 570210
rect 512686 570152 512826 570208
rect 512882 570152 512887 570208
rect 512686 570150 512887 570152
rect 78673 570147 78739 570150
rect 512686 570074 512746 570150
rect 512821 570147 512887 570150
rect 521886 570208 521995 570210
rect 521886 570152 521934 570208
rect 521990 570152 521995 570208
rect 521886 570147 521995 570152
rect 512821 570074 512887 570077
rect 521886 570076 521946 570147
rect 512686 570072 512887 570074
rect 512686 570016 512826 570072
rect 512882 570016 512887 570072
rect 512686 570014 512887 570016
rect 512821 570011 512887 570014
rect 521878 570012 521884 570076
rect 521948 570012 521954 570076
rect 504357 569938 504423 569941
rect 504541 569938 504607 569941
rect 504357 569936 504607 569938
rect 504357 569880 504362 569936
rect 504418 569880 504546 569936
rect 504602 569880 504607 569936
rect 504357 569878 504607 569880
rect 504357 569875 504423 569878
rect 504541 569875 504607 569878
rect 583520 568836 584960 569076
rect 512821 568578 512887 568581
rect 513005 568578 513071 568581
rect 512821 568576 513071 568578
rect 512821 568520 512826 568576
rect 512882 568520 513010 568576
rect 513066 568520 513071 568576
rect 512821 568518 513071 568520
rect 512821 568515 512887 568518
rect 513005 568515 513071 568518
rect 503897 568306 503963 568309
rect 501860 568304 503963 568306
rect 501860 568248 503902 568304
rect 503958 568248 503963 568304
rect 501860 568246 503963 568248
rect 503897 568243 503963 568246
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 78673 566674 78739 566677
rect 78673 566672 82156 566674
rect 78673 566616 78678 566672
rect 78734 566616 82156 566672
rect 78673 566614 82156 566616
rect 78673 566611 78739 566614
rect 503897 564498 503963 564501
rect 501860 564496 503963 564498
rect 501860 564440 503902 564496
rect 503958 564440 503963 564496
rect 501860 564438 503963 564440
rect 503897 564435 503963 564438
rect 521878 563076 521884 563140
rect 521948 563076 521954 563140
rect 78673 562866 78739 562869
rect 521886 562866 521946 563076
rect 522062 562866 522068 562868
rect 78673 562864 82156 562866
rect 78673 562808 78678 562864
rect 78734 562808 82156 562864
rect 78673 562806 82156 562808
rect 521886 562806 522068 562866
rect 78673 562803 78739 562806
rect 522062 562804 522068 562806
rect 522132 562804 522138 562868
rect 503897 560962 503963 560965
rect 501860 560960 503963 560962
rect 501860 560904 503902 560960
rect 503958 560904 503963 560960
rect 501860 560902 503963 560904
rect 503897 560899 503963 560902
rect 522113 560284 522179 560285
rect 522062 560282 522068 560284
rect 522022 560222 522068 560282
rect 522132 560280 522179 560284
rect 522174 560224 522179 560280
rect 522062 560220 522068 560222
rect 522132 560220 522179 560224
rect 522113 560219 522179 560220
rect 79593 559330 79659 559333
rect 79593 559328 82156 559330
rect 79593 559272 79598 559328
rect 79654 559272 82156 559328
rect 79593 559270 82156 559272
rect 79593 559267 79659 559270
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 506422 557154 506428 557156
rect 501860 557094 506428 557154
rect 506422 557092 506428 557094
rect 506492 557092 506498 557156
rect 583520 557140 584960 557230
rect 78673 555794 78739 555797
rect 78673 555792 82156 555794
rect 78673 555736 78678 555792
rect 78734 555736 82156 555792
rect 78673 555734 82156 555736
rect 78673 555731 78739 555734
rect 501638 554916 501644 554980
rect 501708 554916 501714 554980
rect 501646 554842 501706 554916
rect 501822 554842 501828 554844
rect 501646 554782 501828 554842
rect 501822 554780 501828 554782
rect 501892 554780 501898 554844
rect 503897 553618 503963 553621
rect 501860 553616 503963 553618
rect 501860 553560 503902 553616
rect 503958 553560 503963 553616
rect 501860 553558 503963 553560
rect 503897 553555 503963 553558
rect 66846 553420 66852 553484
rect 66916 553420 66922 553484
rect 66854 553210 66914 553420
rect 67030 553210 67036 553212
rect -960 553074 480 553164
rect 66854 553150 67036 553210
rect 67030 553148 67036 553150
rect 67100 553148 67106 553212
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 77150 551924 77156 551988
rect 77220 551986 77226 551988
rect 77220 551926 82156 551986
rect 77220 551924 77226 551926
rect 522113 550762 522179 550765
rect 522246 550762 522252 550764
rect 522113 550760 522252 550762
rect 522113 550704 522118 550760
rect 522174 550704 522252 550760
rect 522113 550702 522252 550704
rect 522113 550699 522179 550702
rect 522246 550700 522252 550702
rect 522316 550700 522322 550764
rect 503897 550082 503963 550085
rect 501860 550080 503963 550082
rect 501860 550024 503902 550080
rect 503958 550024 503963 550080
rect 501860 550022 503963 550024
rect 503897 550019 503963 550022
rect 512821 549266 512887 549269
rect 513005 549266 513071 549269
rect 512821 549264 513071 549266
rect 512821 549208 512826 549264
rect 512882 549208 513010 549264
rect 513066 549208 513071 549264
rect 512821 549206 513071 549208
rect 512821 549203 512887 549206
rect 513005 549203 513071 549206
rect 78254 548388 78260 548452
rect 78324 548450 78330 548452
rect 78324 548390 82156 548450
rect 78324 548388 78330 548390
rect 503897 546274 503963 546277
rect 501860 546272 503963 546274
rect 501860 546216 503902 546272
rect 503958 546216 503963 546272
rect 501860 546214 503963 546216
rect 503897 546211 503963 546214
rect 579889 545594 579955 545597
rect 583520 545594 584960 545684
rect 579889 545592 584960 545594
rect 579889 545536 579894 545592
rect 579950 545536 584960 545592
rect 579889 545534 584960 545536
rect 579889 545531 579955 545534
rect 583520 545444 584960 545534
rect 67030 543900 67036 543964
rect 67100 543900 67106 543964
rect 67038 543556 67098 543900
rect 74206 543764 74212 543828
rect 74276 543826 74282 543828
rect 82126 543826 82186 544612
rect 522246 543962 522252 543964
rect 74276 543766 82186 543826
rect 522070 543902 522252 543962
rect 74276 543764 74282 543766
rect 522070 543692 522130 543902
rect 522246 543900 522252 543902
rect 522316 543900 522322 543964
rect 522062 543628 522068 543692
rect 522132 543628 522138 543692
rect 67030 543492 67036 543556
rect 67100 543492 67106 543556
rect 503897 542738 503963 542741
rect 501860 542736 503963 542738
rect 501860 542680 503902 542736
rect 503958 542680 503963 542736
rect 501860 542678 503963 542680
rect 503897 542675 503963 542678
rect 74390 541044 74396 541108
rect 74460 541106 74466 541108
rect 74460 541046 82156 541106
rect 74460 541044 74466 541046
rect 522021 540972 522087 540973
rect 522021 540970 522068 540972
rect 521976 540968 522068 540970
rect 521976 540912 522026 540968
rect 521976 540910 522068 540912
rect 522021 540908 522068 540910
rect 522132 540908 522138 540972
rect 522021 540907 522087 540908
rect 503897 538930 503963 538933
rect 501860 538928 503963 538930
rect 501860 538872 503902 538928
rect 503958 538872 503963 538928
rect 501860 538870 503963 538872
rect 503897 538867 503963 538870
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 76230 537236 76236 537300
rect 76300 537298 76306 537300
rect 76300 537238 82156 537298
rect 76300 537236 76306 537238
rect 502333 535394 502399 535397
rect 501860 535392 502399 535394
rect 501860 535336 502338 535392
rect 502394 535336 502399 535392
rect 501860 535334 502399 535336
rect 502333 535331 502399 535334
rect 66989 534308 67055 534309
rect 66989 534306 67036 534308
rect 66944 534304 67036 534306
rect 66944 534248 66994 534304
rect 66944 534246 67036 534248
rect 66989 534244 67036 534246
rect 67100 534244 67106 534308
rect 66989 534243 67055 534244
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 81198 533700 81204 533764
rect 81268 533762 81274 533764
rect 81268 533702 82156 533762
rect 583520 533748 584960 533838
rect 81268 533700 81274 533702
rect 66989 531586 67055 531589
rect 504214 531586 504220 531588
rect 66989 531584 67098 531586
rect 66989 531528 66994 531584
rect 67050 531528 67098 531584
rect 66989 531523 67098 531528
rect 501860 531526 504220 531586
rect 504214 531524 504220 531526
rect 504284 531524 504290 531588
rect 522021 531586 522087 531589
rect 521886 531584 522087 531586
rect 521886 531528 522026 531584
rect 522082 531528 522087 531584
rect 521886 531526 522087 531528
rect 67038 531452 67098 531523
rect 521886 531452 521946 531526
rect 522021 531523 522087 531526
rect 67030 531388 67036 531452
rect 67100 531388 67106 531452
rect 521878 531388 521884 531452
rect 521948 531388 521954 531452
rect 79869 530226 79935 530229
rect 79869 530224 82156 530226
rect 79869 530168 79874 530224
rect 79930 530168 82156 530224
rect 79869 530166 82156 530168
rect 79869 530163 79935 530166
rect 78673 526418 78739 526421
rect 78673 526416 82156 526418
rect 78673 526360 78678 526416
rect 78734 526360 82156 526416
rect 78673 526358 82156 526360
rect 78673 526355 78739 526358
rect 501270 526356 501276 526420
rect 501340 526418 501346 526420
rect 501781 526418 501847 526421
rect 501340 526416 501847 526418
rect 501340 526360 501786 526416
rect 501842 526360 501847 526416
rect 501340 526358 501847 526360
rect 501340 526356 501346 526358
rect 501781 526355 501847 526358
rect 67030 524786 67036 524788
rect 66670 524726 67036 524786
rect -960 524092 480 524332
rect 66670 524244 66730 524726
rect 67030 524724 67036 524726
rect 67100 524724 67106 524788
rect 501873 524786 501939 524789
rect 502006 524786 502012 524788
rect 501873 524784 502012 524786
rect 501873 524728 501878 524784
rect 501934 524728 502012 524784
rect 501873 524726 502012 524728
rect 501873 524723 501939 524726
rect 502006 524724 502012 524726
rect 502076 524724 502082 524788
rect 503897 524514 503963 524517
rect 501860 524512 503963 524514
rect 501860 524456 503902 524512
rect 503958 524456 503963 524512
rect 501860 524454 503963 524456
rect 503897 524451 503963 524454
rect 521878 524452 521884 524516
rect 521948 524452 521954 524516
rect 66662 524180 66668 524244
rect 66732 524180 66738 524244
rect 521886 524242 521946 524452
rect 522062 524242 522068 524244
rect 521886 524182 522068 524242
rect 522062 524180 522068 524182
rect 522132 524180 522138 524244
rect 79726 522820 79732 522884
rect 79796 522882 79802 522884
rect 79796 522822 82156 522882
rect 79796 522820 79802 522822
rect 501270 522820 501276 522884
rect 501340 522882 501346 522884
rect 501781 522882 501847 522885
rect 501340 522880 501847 522882
rect 501340 522824 501786 522880
rect 501842 522824 501847 522880
rect 501340 522822 501847 522824
rect 501340 522820 501346 522822
rect 501781 522819 501847 522822
rect 501873 522340 501939 522341
rect 501822 522338 501828 522340
rect 501782 522278 501828 522338
rect 501892 522336 501939 522340
rect 501934 522280 501939 522336
rect 501822 522276 501828 522278
rect 501892 522276 501939 522280
rect 501873 522275 501939 522276
rect 583520 521916 584960 522156
rect 66529 521658 66595 521661
rect 522021 521660 522087 521661
rect 66662 521658 66668 521660
rect 66529 521656 66668 521658
rect 66529 521600 66534 521656
rect 66590 521600 66668 521656
rect 66529 521598 66668 521600
rect 66529 521595 66595 521598
rect 66662 521596 66668 521598
rect 66732 521596 66738 521660
rect 522021 521658 522068 521660
rect 521976 521656 522068 521658
rect 521976 521600 522026 521656
rect 521976 521598 522068 521600
rect 522021 521596 522068 521598
rect 522132 521596 522138 521660
rect 522021 521595 522087 521596
rect 503897 520706 503963 520709
rect 501860 520704 503963 520706
rect 501860 520648 503902 520704
rect 503958 520648 503963 520704
rect 501860 520646 503963 520648
rect 503897 520643 503963 520646
rect 78857 519074 78923 519077
rect 78857 519072 82156 519074
rect 78857 519016 78862 519072
rect 78918 519016 82156 519072
rect 78857 519014 82156 519016
rect 78857 519011 78923 519014
rect 502558 517170 502564 517172
rect 501860 517110 502564 517170
rect 502558 517108 502564 517110
rect 502628 517108 502634 517172
rect 81566 515476 81572 515540
rect 81636 515538 81642 515540
rect 81636 515478 82156 515538
rect 81636 515476 81642 515478
rect 505686 513362 505692 513364
rect 501860 513302 505692 513362
rect 505686 513300 505692 513302
rect 505756 513300 505762 513364
rect 66529 512274 66595 512277
rect 522021 512274 522087 512277
rect 66486 512272 66595 512274
rect 66486 512216 66534 512272
rect 66590 512216 66595 512272
rect 66486 512211 66595 512216
rect 521886 512272 522087 512274
rect 521886 512216 522026 512272
rect 522082 512216 522087 512272
rect 521886 512214 522087 512216
rect 66486 512140 66546 512211
rect 521886 512140 521946 512214
rect 522021 512211 522087 512214
rect 66478 512076 66484 512140
rect 66548 512076 66554 512140
rect 521878 512076 521884 512140
rect 521948 512076 521954 512140
rect 78673 511730 78739 511733
rect 78673 511728 82156 511730
rect 78673 511672 78678 511728
rect 78734 511672 82156 511728
rect 78673 511670 82156 511672
rect 78673 511667 78739 511670
rect 66478 510444 66484 510508
rect 66548 510444 66554 510508
rect 66486 510370 66546 510444
rect 66621 510370 66687 510373
rect 66486 510368 66687 510370
rect 66486 510312 66626 510368
rect 66682 510312 66687 510368
rect 66486 510310 66687 510312
rect 66621 510307 66687 510310
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3141 509962 3207 509965
rect -960 509960 3207 509962
rect -960 509904 3146 509960
rect 3202 509904 3207 509960
rect -960 509902 3207 509904
rect -960 509812 480 509902
rect 3141 509899 3207 509902
rect 502742 509826 502748 509828
rect 501860 509766 502748 509826
rect 502742 509764 502748 509766
rect 502812 509764 502818 509828
rect 78673 508194 78739 508197
rect 78673 508192 82156 508194
rect 78673 508136 78678 508192
rect 78734 508136 82156 508192
rect 78673 508134 82156 508136
rect 78673 508131 78739 508134
rect 502057 507788 502123 507789
rect 502006 507724 502012 507788
rect 502076 507786 502123 507788
rect 502076 507784 502168 507786
rect 502118 507728 502168 507784
rect 502076 507726 502168 507728
rect 502076 507724 502123 507726
rect 502057 507723 502123 507724
rect 501462 505612 501522 505988
rect 501454 505548 501460 505612
rect 501524 505548 501530 505612
rect 521878 505202 521884 505204
rect 521702 505142 521884 505202
rect 521702 504932 521762 505142
rect 521878 505140 521884 505142
rect 521948 505140 521954 505204
rect 521694 504868 521700 504932
rect 521764 504868 521770 504932
rect 78673 504658 78739 504661
rect 78673 504656 82156 504658
rect 78673 504600 78678 504656
rect 78734 504600 82156 504656
rect 78673 504598 82156 504600
rect 78673 504595 78739 504598
rect 510654 502482 510660 502484
rect 501860 502422 510660 502482
rect 510654 502420 510660 502422
rect 510724 502420 510730 502484
rect 521694 502284 521700 502348
rect 521764 502346 521770 502348
rect 522021 502346 522087 502349
rect 521764 502344 522087 502346
rect 521764 502288 522026 502344
rect 522082 502288 522087 502344
rect 521764 502286 522087 502288
rect 521764 502284 521770 502286
rect 522021 502283 522087 502286
rect 66621 500986 66687 500989
rect 67030 500986 67036 500988
rect 66621 500984 67036 500986
rect 66621 500928 66626 500984
rect 66682 500928 67036 500984
rect 66621 500926 67036 500928
rect 66621 500923 66687 500926
rect 67030 500924 67036 500926
rect 67100 500924 67106 500988
rect 512821 500986 512887 500989
rect 513005 500986 513071 500989
rect 512821 500984 513071 500986
rect 512821 500928 512826 500984
rect 512882 500928 513010 500984
rect 513066 500928 513071 500984
rect 512821 500926 513071 500928
rect 512821 500923 512887 500926
rect 513005 500923 513071 500926
rect 79041 500850 79107 500853
rect 79041 500848 82156 500850
rect 79041 500792 79046 500848
rect 79102 500792 82156 500848
rect 79041 500790 82156 500792
rect 79041 500787 79107 500790
rect 503897 498946 503963 498949
rect 501860 498944 503963 498946
rect 501860 498888 503902 498944
rect 503958 498888 503963 498944
rect 501860 498886 503963 498888
rect 503897 498883 503963 498886
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect 502057 498402 502123 498405
rect 502014 498400 502123 498402
rect 502014 498344 502062 498400
rect 502118 498344 502123 498400
rect 502014 498339 502123 498344
rect 502014 498268 502074 498339
rect 502006 498204 502012 498268
rect 502076 498204 502082 498268
rect 78673 497314 78739 497317
rect 78673 497312 82156 497314
rect 78673 497256 78678 497312
rect 78734 497256 82156 497312
rect 78673 497254 82156 497256
rect 78673 497251 78739 497254
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 503897 495138 503963 495141
rect 501860 495136 503963 495138
rect 501860 495080 503902 495136
rect 503958 495080 503963 495136
rect 501860 495078 503963 495080
rect 503897 495075 503963 495078
rect 79501 493506 79567 493509
rect 79501 493504 82156 493506
rect 79501 493448 79506 493504
rect 79562 493448 82156 493504
rect 79501 493446 82156 493448
rect 79501 493443 79567 493446
rect 504173 492690 504239 492693
rect 504357 492690 504423 492693
rect 504173 492688 504423 492690
rect 504173 492632 504178 492688
rect 504234 492632 504362 492688
rect 504418 492632 504423 492688
rect 504173 492630 504423 492632
rect 504173 492627 504239 492630
rect 504357 492627 504423 492630
rect 521878 492628 521884 492692
rect 521948 492690 521954 492692
rect 522021 492690 522087 492693
rect 521948 492688 522087 492690
rect 521948 492632 522026 492688
rect 522082 492632 522087 492688
rect 521948 492630 522087 492632
rect 521948 492628 521954 492630
rect 522021 492627 522087 492630
rect 66989 491196 67055 491197
rect 66989 491194 67036 491196
rect 66944 491192 67036 491194
rect 66944 491136 66994 491192
rect 66944 491134 67036 491136
rect 66989 491132 67036 491134
rect 67100 491132 67106 491196
rect 66989 491131 67055 491132
rect 501462 491060 501522 491572
rect 501454 490996 501460 491060
rect 501524 490996 501530 491060
rect 79542 489908 79548 489972
rect 79612 489970 79618 489972
rect 79612 489910 82156 489970
rect 79612 489908 79618 489910
rect 503897 487794 503963 487797
rect 501860 487792 503963 487794
rect 501860 487736 503902 487792
rect 503958 487736 503963 487792
rect 501860 487734 503963 487736
rect 503897 487731 503963 487734
rect 501638 487460 501644 487524
rect 501708 487522 501714 487524
rect 502006 487522 502012 487524
rect 501708 487462 502012 487522
rect 501708 487460 501714 487462
rect 502006 487460 502012 487462
rect 502076 487460 502082 487524
rect 33726 487188 33732 487252
rect 33796 487250 33802 487252
rect 46790 487250 46796 487252
rect 33796 487190 46796 487250
rect 33796 487188 33802 487190
rect 46790 487188 46796 487190
rect 46860 487188 46866 487252
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 78673 486162 78739 486165
rect 78673 486160 82156 486162
rect 78673 486104 78678 486160
rect 78734 486104 82156 486160
rect 78673 486102 82156 486104
rect 78673 486099 78739 486102
rect 17902 485828 17908 485892
rect 17972 485890 17978 485892
rect 27470 485890 27476 485892
rect 17972 485830 27476 485890
rect 17972 485828 17978 485830
rect 27470 485828 27476 485830
rect 27540 485828 27546 485892
rect 521878 485890 521884 485892
rect 521702 485830 521884 485890
rect 521702 485620 521762 485830
rect 521878 485828 521884 485830
rect 521948 485828 521954 485892
rect 521694 485556 521700 485620
rect 521764 485556 521770 485620
rect 503897 484258 503963 484261
rect 501860 484256 503963 484258
rect 501860 484200 503902 484256
rect 503958 484200 503963 484256
rect 501860 484198 503963 484200
rect 503897 484195 503963 484198
rect 66989 483716 67055 483717
rect 66989 483714 67036 483716
rect 66944 483712 67036 483714
rect 66944 483656 66994 483712
rect 66944 483654 67036 483656
rect 66989 483652 67036 483654
rect 67100 483652 67106 483716
rect 66989 483651 67055 483652
rect 80973 482626 81039 482629
rect 80973 482624 82156 482626
rect 80973 482568 80978 482624
rect 81034 482568 82156 482624
rect 80973 482566 82156 482568
rect 80973 482563 81039 482566
rect 501965 481540 502031 481541
rect 501965 481538 502012 481540
rect 501920 481536 502012 481538
rect 501920 481480 501970 481536
rect 501920 481478 502012 481480
rect 501965 481476 502012 481478
rect 502076 481476 502082 481540
rect 501965 481475 502031 481476
rect -960 481130 480 481220
rect 3785 481130 3851 481133
rect -960 481128 3851 481130
rect -960 481072 3790 481128
rect 3846 481072 3851 481128
rect -960 481070 3851 481072
rect -960 480980 480 481070
rect 3785 481067 3851 481070
rect 505870 480450 505876 480452
rect 501860 480390 505876 480450
rect 505870 480388 505876 480390
rect 505940 480388 505946 480452
rect 78673 479090 78739 479093
rect 78673 479088 82156 479090
rect 78673 479032 78678 479088
rect 78734 479032 82156 479088
rect 78673 479030 82156 479032
rect 78673 479027 78739 479030
rect 66989 478820 67055 478821
rect 66989 478818 67036 478820
rect 66944 478816 67036 478818
rect 66944 478760 66994 478816
rect 66944 478758 67036 478760
rect 66989 478756 67036 478758
rect 67100 478756 67106 478820
rect 66989 478755 67055 478756
rect 503897 476914 503963 476917
rect 501860 476912 503963 476914
rect 501860 476856 503902 476912
rect 503958 476856 503963 476912
rect 501860 476854 503963 476856
rect 503897 476851 503963 476854
rect 521694 476036 521700 476100
rect 521764 476098 521770 476100
rect 522430 476098 522436 476100
rect 521764 476038 522436 476098
rect 521764 476036 521770 476038
rect 522430 476036 522436 476038
rect 522500 476036 522506 476100
rect 82494 475012 82554 475252
rect 82486 474948 82492 475012
rect 82556 474948 82562 475012
rect 583520 474996 584960 475236
rect 503897 473378 503963 473381
rect 501860 473376 503963 473378
rect 501860 473320 503902 473376
rect 503958 473320 503963 473376
rect 501860 473318 503963 473320
rect 503897 473315 503963 473318
rect 504449 473378 504515 473381
rect 504633 473378 504699 473381
rect 504449 473376 504699 473378
rect 504449 473320 504454 473376
rect 504510 473320 504638 473376
rect 504694 473320 504699 473376
rect 504449 473318 504699 473320
rect 504449 473315 504515 473318
rect 504633 473315 504699 473318
rect 501965 472020 502031 472021
rect 501965 472016 502012 472020
rect 502076 472018 502082 472020
rect 501965 471960 501970 472016
rect 501965 471956 502012 471960
rect 502076 471958 502122 472018
rect 502076 471956 502082 471958
rect 501965 471955 502031 471956
rect 502057 471884 502123 471885
rect 502006 471820 502012 471884
rect 502076 471882 502123 471884
rect 502076 471880 502168 471882
rect 502118 471824 502168 471880
rect 502076 471822 502168 471824
rect 502076 471820 502123 471822
rect 502057 471819 502123 471820
rect 78673 471746 78739 471749
rect 78673 471744 82156 471746
rect 78673 471688 78678 471744
rect 78734 471688 82156 471744
rect 78673 471686 82156 471688
rect 78673 471683 78739 471686
rect 503897 469570 503963 469573
rect 501860 469568 503963 469570
rect 501860 469512 503902 469568
rect 503958 469512 503963 469568
rect 501860 469510 503963 469512
rect 503897 469507 503963 469510
rect 66989 469436 67055 469437
rect 66989 469432 67036 469436
rect 67100 469434 67106 469436
rect 66989 469376 66994 469432
rect 66989 469372 67036 469376
rect 67100 469374 67146 469434
rect 67100 469372 67106 469374
rect 66989 469371 67055 469372
rect 66897 469162 66963 469165
rect 67030 469162 67036 469164
rect 66897 469160 67036 469162
rect 66897 469104 66902 469160
rect 66958 469104 67036 469160
rect 66897 469102 67036 469104
rect 66897 469099 66963 469102
rect 67030 469100 67036 469102
rect 67100 469100 67106 469164
rect 82494 467668 82554 467908
rect 82486 467604 82492 467668
rect 82556 467604 82562 467668
rect -960 466700 480 466940
rect 522430 466578 522436 466580
rect 522254 466518 522436 466578
rect 522254 466308 522314 466518
rect 522430 466516 522436 466518
rect 522500 466516 522506 466580
rect 522246 466244 522252 466308
rect 522316 466244 522322 466308
rect 506606 466034 506612 466036
rect 501860 465974 506612 466034
rect 506606 465972 506612 465974
rect 506676 465972 506682 466036
rect 81433 464402 81499 464405
rect 81433 464400 82156 464402
rect 81433 464344 81438 464400
rect 81494 464344 82156 464400
rect 81433 464342 82156 464344
rect 81433 464339 81499 464342
rect 522246 463524 522252 463588
rect 522316 463524 522322 463588
rect 522113 463450 522179 463453
rect 522254 463450 522314 463524
rect 522113 463448 522314 463450
rect 522113 463392 522118 463448
rect 522174 463392 522314 463448
rect 522113 463390 522314 463392
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 522113 463387 522179 463390
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 502057 462636 502123 462637
rect 502006 462634 502012 462636
rect 501966 462574 502012 462634
rect 502076 462632 502123 462636
rect 502118 462576 502123 462632
rect 502006 462572 502012 462574
rect 502076 462572 502123 462576
rect 502057 462571 502123 462572
rect 503897 462226 503963 462229
rect 501860 462224 503963 462226
rect 501860 462168 503902 462224
rect 503958 462168 503963 462224
rect 501860 462166 503963 462168
rect 503897 462163 503963 462166
rect 78673 460594 78739 460597
rect 78673 460592 82156 460594
rect 78673 460536 78678 460592
rect 78734 460536 82156 460592
rect 78673 460534 82156 460536
rect 78673 460531 78739 460534
rect 66897 459778 66963 459781
rect 66854 459776 66963 459778
rect 66854 459720 66902 459776
rect 66958 459720 66963 459776
rect 66854 459715 66963 459720
rect 66854 459644 66914 459715
rect 66846 459580 66852 459644
rect 66916 459580 66922 459644
rect 501638 458900 501644 458964
rect 501708 458962 501714 458964
rect 501965 458962 502031 458965
rect 501708 458960 502031 458962
rect 501708 458904 501970 458960
rect 502026 458904 502031 458960
rect 501708 458902 502031 458904
rect 501708 458900 501714 458902
rect 501965 458899 502031 458902
rect 501646 458284 501706 458660
rect 501638 458220 501644 458284
rect 501708 458220 501714 458284
rect 78673 457058 78739 457061
rect 78673 457056 82156 457058
rect 78673 457000 78678 457056
rect 78734 457000 82156 457056
rect 78673 456998 82156 457000
rect 78673 456995 78739 456998
rect 506790 454882 506796 454884
rect 501860 454822 506796 454882
rect 506790 454820 506796 454822
rect 506860 454820 506866 454884
rect 504173 454066 504239 454069
rect 504357 454066 504423 454069
rect 504173 454064 504423 454066
rect 504173 454008 504178 454064
rect 504234 454008 504362 454064
rect 504418 454008 504423 454064
rect 504173 454006 504423 454008
rect 504173 454003 504239 454006
rect 504357 454003 504423 454006
rect 521878 454004 521884 454068
rect 521948 454066 521954 454068
rect 522113 454066 522179 454069
rect 521948 454064 522179 454066
rect 521948 454008 522118 454064
rect 522174 454008 522179 454064
rect 521948 454006 522179 454008
rect 521948 454004 521954 454006
rect 522113 454003 522179 454006
rect 82678 452981 82738 453492
rect 82629 452976 82738 452981
rect 82629 452920 82634 452976
rect 82690 452920 82738 452976
rect 82629 452918 82738 452920
rect 82629 452915 82695 452918
rect 501965 452708 502031 452709
rect 501965 452704 502012 452708
rect 502076 452706 502082 452708
rect 501965 452648 501970 452704
rect 501965 452644 502012 452648
rect 502076 452646 502122 452706
rect 502076 452644 502082 452646
rect 501965 452643 502031 452644
rect 10174 452570 10180 452572
rect -960 452434 480 452524
rect 614 452510 10180 452570
rect 614 452434 674 452510
rect 10174 452508 10180 452510
rect 10244 452508 10250 452572
rect -960 452374 674 452434
rect -960 452284 480 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 502333 451346 502399 451349
rect 501860 451344 502399 451346
rect 501860 451288 502338 451344
rect 502394 451288 502399 451344
rect 501860 451286 502399 451288
rect 502333 451283 502399 451286
rect 78673 449714 78739 449717
rect 78673 449712 82156 449714
rect 78673 449656 78678 449712
rect 78734 449656 82156 449712
rect 78673 449654 82156 449656
rect 78673 449651 78739 449654
rect 503897 447810 503963 447813
rect 501860 447808 503963 447810
rect 501860 447752 503902 447808
rect 503958 447752 503963 447808
rect 501860 447750 503963 447752
rect 503897 447747 503963 447750
rect 521878 447204 521884 447268
rect 521948 447204 521954 447268
rect 521886 446994 521946 447204
rect 522062 446994 522068 446996
rect 521886 446934 522068 446994
rect 522062 446932 522068 446934
rect 522132 446932 522138 446996
rect 66713 446450 66779 446453
rect 67030 446450 67036 446452
rect 66713 446448 67036 446450
rect 66713 446392 66718 446448
rect 66774 446392 67036 446448
rect 66713 446390 67036 446392
rect 66713 446387 66779 446390
rect 67030 446388 67036 446390
rect 67100 446388 67106 446452
rect 78673 446178 78739 446181
rect 78673 446176 82156 446178
rect 78673 446120 78678 446176
rect 78734 446120 82156 446176
rect 78673 446118 82156 446120
rect 78673 446115 78739 446118
rect 503897 444002 503963 444005
rect 501860 444000 503963 444002
rect 501860 443944 503902 444000
rect 503958 443944 503963 444000
rect 501860 443942 503963 443944
rect 503897 443939 503963 443942
rect 502057 442916 502123 442917
rect 502006 442852 502012 442916
rect 502076 442914 502123 442916
rect 502076 442912 502168 442914
rect 502118 442856 502168 442912
rect 502076 442854 502168 442856
rect 502076 442852 502123 442854
rect 502057 442851 502123 442852
rect 78673 442370 78739 442373
rect 78673 442368 82156 442370
rect 78673 442312 78678 442368
rect 78734 442312 82156 442368
rect 78673 442310 82156 442312
rect 78673 442307 78739 442310
rect 503897 440466 503963 440469
rect 501860 440464 503963 440466
rect 501860 440408 503902 440464
rect 503958 440408 503963 440464
rect 501860 440406 503963 440408
rect 503897 440403 503963 440406
rect 579613 439922 579679 439925
rect 583520 439922 584960 440012
rect 579613 439920 584960 439922
rect 579613 439864 579618 439920
rect 579674 439864 584960 439920
rect 579613 439862 584960 439864
rect 579613 439859 579679 439862
rect 583520 439772 584960 439862
rect 78489 438834 78555 438837
rect 78489 438832 82156 438834
rect 78489 438776 78494 438832
rect 78550 438776 82156 438832
rect 78489 438774 82156 438776
rect 78489 438771 78555 438774
rect -960 438018 480 438108
rect 3417 438018 3483 438021
rect -960 438016 3483 438018
rect -960 437960 3422 438016
rect 3478 437960 3483 438016
rect -960 437958 3483 437960
rect -960 437868 480 437958
rect 3417 437955 3483 437958
rect 521694 437412 521700 437476
rect 521764 437474 521770 437476
rect 522246 437474 522252 437476
rect 521764 437414 522252 437474
rect 521764 437412 521770 437414
rect 522246 437412 522252 437414
rect 522316 437412 522322 437476
rect 503897 436658 503963 436661
rect 501860 436656 503963 436658
rect 501860 436600 503902 436656
rect 503958 436600 503963 436656
rect 501860 436598 503963 436600
rect 503897 436595 503963 436598
rect 78581 435026 78647 435029
rect 78581 435024 82156 435026
rect 78581 434968 78586 435024
rect 78642 434968 82156 435024
rect 78581 434966 82156 434968
rect 78581 434963 78647 434966
rect 66713 434756 66779 434757
rect 66662 434754 66668 434756
rect 66622 434694 66668 434754
rect 66732 434752 66779 434756
rect 66774 434696 66779 434752
rect 66662 434692 66668 434694
rect 66732 434692 66779 434696
rect 66713 434691 66779 434692
rect 66989 434618 67055 434621
rect 67398 434618 67404 434620
rect 66989 434616 67404 434618
rect 66989 434560 66994 434616
rect 67050 434560 67404 434616
rect 66989 434558 67404 434560
rect 66989 434555 67055 434558
rect 67398 434556 67404 434558
rect 67468 434556 67474 434620
rect 502057 433396 502123 433397
rect 502006 433394 502012 433396
rect 501966 433334 502012 433394
rect 502076 433392 502123 433396
rect 502118 433336 502123 433392
rect 502006 433332 502012 433334
rect 502076 433332 502123 433336
rect 502057 433331 502123 433332
rect 503897 433122 503963 433125
rect 501860 433120 503963 433122
rect 501860 433064 503902 433120
rect 503958 433064 503963 433120
rect 501860 433062 503963 433064
rect 503897 433059 503963 433062
rect 78673 431490 78739 431493
rect 78673 431488 82156 431490
rect 78673 431432 78678 431488
rect 78734 431432 82156 431488
rect 78673 431430 82156 431432
rect 78673 431427 78739 431430
rect 501689 430674 501755 430677
rect 501646 430672 501755 430674
rect 501646 430616 501694 430672
rect 501750 430616 501755 430672
rect 501646 430611 501755 430616
rect 501646 430538 501706 430611
rect 501873 430538 501939 430541
rect 501646 430536 501939 430538
rect 501646 430480 501878 430536
rect 501934 430480 501939 430536
rect 501646 430478 501939 430480
rect 501873 430475 501939 430478
rect 66989 429858 67055 429861
rect 67398 429858 67404 429860
rect 66989 429856 67404 429858
rect 66989 429800 66994 429856
rect 67050 429800 67404 429856
rect 66989 429798 67404 429800
rect 66989 429795 67055 429798
rect 67398 429796 67404 429798
rect 67468 429796 67474 429860
rect 503897 429314 503963 429317
rect 501860 429312 503963 429314
rect 501860 429256 503902 429312
rect 503958 429256 503963 429312
rect 501860 429254 503963 429256
rect 503897 429251 503963 429254
rect 502057 428500 502123 428501
rect 502006 428436 502012 428500
rect 502076 428498 502123 428500
rect 502076 428496 502168 428498
rect 502118 428440 502168 428496
rect 502076 428438 502168 428440
rect 502076 428436 502123 428438
rect 502057 428435 502123 428436
rect 583520 428076 584960 428316
rect 78673 427954 78739 427957
rect 522246 427954 522252 427956
rect 78673 427952 82156 427954
rect 78673 427896 78678 427952
rect 78734 427896 82156 427952
rect 78673 427894 82156 427896
rect 522070 427894 522252 427954
rect 78673 427891 78739 427894
rect 522070 427684 522130 427894
rect 522246 427892 522252 427894
rect 522316 427892 522322 427956
rect 522062 427620 522068 427684
rect 522132 427620 522138 427684
rect 503897 425778 503963 425781
rect 501860 425776 503963 425778
rect 501860 425720 503902 425776
rect 503958 425720 503963 425776
rect 501860 425718 503963 425720
rect 503897 425715 503963 425718
rect 522062 424900 522068 424964
rect 522132 424962 522138 424964
rect 522205 424962 522271 424965
rect 522132 424960 522271 424962
rect 522132 424904 522210 424960
rect 522266 424904 522271 424960
rect 522132 424902 522271 424904
rect 522132 424900 522138 424902
rect 522205 424899 522271 424902
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 74022 423676 74028 423740
rect 74092 423738 74098 423740
rect 82126 423738 82186 424116
rect 74092 423678 82186 423738
rect 74092 423676 74098 423678
rect 503897 422242 503963 422245
rect 501860 422240 503963 422242
rect 501860 422184 503902 422240
rect 503958 422184 503963 422240
rect 501860 422182 503963 422184
rect 503897 422179 503963 422182
rect 78673 420610 78739 420613
rect 78673 420608 82156 420610
rect 78673 420552 78678 420608
rect 78734 420552 82156 420608
rect 78673 420550 82156 420552
rect 78673 420547 78739 420550
rect 509366 418434 509372 418436
rect 501860 418374 509372 418434
rect 509366 418372 509372 418374
rect 509436 418372 509442 418436
rect 78673 416802 78739 416805
rect 78673 416800 82156 416802
rect 78673 416744 78678 416800
rect 78734 416744 82156 416800
rect 78673 416742 82156 416744
rect 78673 416739 78739 416742
rect 580349 416530 580415 416533
rect 583520 416530 584960 416620
rect 580349 416528 584960 416530
rect 580349 416472 580354 416528
rect 580410 416472 584960 416528
rect 580349 416470 584960 416472
rect 580349 416467 580415 416470
rect 583520 416380 584960 416470
rect 501965 415444 502031 415445
rect 501965 415440 502012 415444
rect 502076 415442 502082 415444
rect 501965 415384 501970 415440
rect 501965 415380 502012 415384
rect 502076 415382 502122 415442
rect 502076 415380 502082 415382
rect 521878 415380 521884 415444
rect 521948 415442 521954 415444
rect 522205 415442 522271 415445
rect 521948 415440 522271 415442
rect 521948 415384 522210 415440
rect 522266 415384 522271 415440
rect 521948 415382 522271 415384
rect 521948 415380 521954 415382
rect 501965 415379 502031 415380
rect 522205 415379 522271 415382
rect 502425 414898 502491 414901
rect 501860 414896 502491 414898
rect 501860 414840 502430 414896
rect 502486 414840 502491 414896
rect 501860 414838 502491 414840
rect 502425 414835 502491 414838
rect 502057 413948 502123 413949
rect 502006 413884 502012 413948
rect 502076 413946 502123 413948
rect 502076 413944 502168 413946
rect 502118 413888 502168 413944
rect 502076 413886 502168 413888
rect 502076 413884 502123 413886
rect 502057 413883 502123 413884
rect 78673 413266 78739 413269
rect 78673 413264 82156 413266
rect 78673 413208 78678 413264
rect 78734 413208 82156 413264
rect 78673 413206 82156 413208
rect 78673 413203 78739 413206
rect 502517 411090 502583 411093
rect 501860 411088 502583 411090
rect 501860 411032 502522 411088
rect 502578 411032 502583 411088
rect 501860 411030 502583 411032
rect 502517 411027 502583 411030
rect 81525 409458 81591 409461
rect 81525 409456 82156 409458
rect -960 409172 480 409412
rect 81525 409400 81530 409456
rect 81586 409400 82156 409456
rect 81525 409398 82156 409400
rect 81525 409395 81591 409398
rect 521878 408642 521884 408644
rect 521702 408582 521884 408642
rect 521702 408372 521762 408582
rect 521878 408580 521884 408582
rect 521948 408580 521954 408644
rect 521694 408308 521700 408372
rect 521764 408308 521770 408372
rect 503897 407554 503963 407557
rect 501860 407552 503963 407554
rect 501860 407496 503902 407552
rect 503958 407496 503963 407552
rect 501860 407494 503963 407496
rect 503897 407491 503963 407494
rect 78673 405922 78739 405925
rect 78673 405920 82156 405922
rect 78673 405864 78678 405920
rect 78734 405864 82156 405920
rect 78673 405862 82156 405864
rect 78673 405859 78739 405862
rect 521694 405588 521700 405652
rect 521764 405588 521770 405652
rect 521702 405514 521762 405588
rect 522205 405514 522271 405517
rect 521702 405512 522271 405514
rect 521702 405456 522210 405512
rect 522266 405456 522271 405512
rect 521702 405454 522271 405456
rect 522205 405451 522271 405454
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 502057 404562 502123 404565
rect 502014 404560 502123 404562
rect 502014 404504 502062 404560
rect 502118 404504 502123 404560
rect 502014 404499 502123 404504
rect 502014 404428 502074 404499
rect 502006 404364 502012 404428
rect 502076 404364 502082 404428
rect 503897 403746 503963 403749
rect 501860 403744 503963 403746
rect 501860 403688 503902 403744
rect 503958 403688 503963 403744
rect 501860 403686 503963 403688
rect 503897 403683 503963 403686
rect 78673 402386 78739 402389
rect 78673 402384 82156 402386
rect 78673 402328 78678 402384
rect 78734 402328 82156 402384
rect 78673 402326 82156 402328
rect 78673 402323 78739 402326
rect 503897 400210 503963 400213
rect 501860 400208 503963 400210
rect 501860 400152 503902 400208
rect 503958 400152 503963 400208
rect 501860 400150 503963 400152
rect 503897 400147 503963 400150
rect 66897 398986 66963 398989
rect 67214 398986 67220 398988
rect 66897 398984 67220 398986
rect 66897 398928 66902 398984
rect 66958 398928 67220 398984
rect 66897 398926 67220 398928
rect 66897 398923 66963 398926
rect 67214 398924 67220 398926
rect 67284 398924 67290 398988
rect 78673 398578 78739 398581
rect 78673 398576 82156 398578
rect 78673 398520 78678 398576
rect 78734 398520 82156 398576
rect 78673 398518 82156 398520
rect 78673 398515 78739 398518
rect 505093 396674 505159 396677
rect 501860 396672 505159 396674
rect 501860 396616 505098 396672
rect 505154 396616 505159 396672
rect 501860 396614 505159 396616
rect 505093 396611 505159 396614
rect 66897 396132 66963 396133
rect 66846 396130 66852 396132
rect 66806 396070 66852 396130
rect 66916 396128 66963 396132
rect 66958 396072 66963 396128
rect 66846 396068 66852 396070
rect 66916 396068 66963 396072
rect 66897 396067 66963 396068
rect 504449 396130 504515 396133
rect 504633 396130 504699 396133
rect 504449 396128 504699 396130
rect 504449 396072 504454 396128
rect 504510 396072 504638 396128
rect 504694 396072 504699 396128
rect 504449 396070 504699 396072
rect 504449 396067 504515 396070
rect 504633 396067 504699 396070
rect 521878 396068 521884 396132
rect 521948 396130 521954 396132
rect 522205 396130 522271 396133
rect 521948 396128 522271 396130
rect 521948 396072 522210 396128
rect 522266 396072 522271 396128
rect 521948 396070 522271 396072
rect 521948 396068 521954 396070
rect 522205 396067 522271 396070
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 78397 395042 78463 395045
rect 78397 395040 82156 395042
rect 78397 394984 78402 395040
rect 78458 394984 82156 395040
rect 78397 394982 82156 394984
rect 78397 394979 78463 394982
rect 502057 394636 502123 394637
rect 66846 394572 66852 394636
rect 66916 394572 66922 394636
rect 502006 394572 502012 394636
rect 502076 394634 502123 394636
rect 502076 394632 502168 394634
rect 502118 394576 502168 394632
rect 502076 394574 502168 394576
rect 502076 394572 502123 394574
rect 66854 394498 66914 394572
rect 502057 394571 502123 394572
rect 67030 394498 67036 394500
rect 66854 394438 67036 394498
rect 67030 394436 67036 394438
rect 67100 394436 67106 394500
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 505185 392866 505251 392869
rect 501860 392864 505251 392866
rect 501860 392808 505190 392864
rect 505246 392808 505251 392864
rect 583520 392852 584960 392942
rect 501860 392806 505251 392808
rect 505185 392803 505251 392806
rect 79869 391234 79935 391237
rect 79869 391232 82156 391234
rect 79869 391176 79874 391232
rect 79930 391176 82156 391232
rect 79869 391174 82156 391176
rect 79869 391171 79935 391174
rect 503897 389330 503963 389333
rect 501860 389328 503963 389330
rect 501860 389272 503902 389328
rect 503958 389272 503963 389328
rect 501860 389270 503963 389272
rect 503897 389267 503963 389270
rect 521878 389268 521884 389332
rect 521948 389268 521954 389332
rect 521886 389058 521946 389268
rect 522062 389058 522068 389060
rect 521886 388998 522068 389058
rect 522062 388996 522068 388998
rect 522132 388996 522138 389060
rect 78673 387698 78739 387701
rect 78673 387696 82156 387698
rect 78673 387640 78678 387696
rect 78734 387640 82156 387696
rect 78673 387638 82156 387640
rect 78673 387635 78739 387638
rect 522062 386276 522068 386340
rect 522132 386276 522138 386340
rect 522070 386202 522130 386276
rect 522205 386202 522271 386205
rect 522070 386200 522271 386202
rect 522070 386144 522210 386200
rect 522266 386144 522271 386200
rect 522070 386142 522271 386144
rect 522205 386139 522271 386142
rect 503897 385522 503963 385525
rect 501860 385520 503963 385522
rect 501860 385464 503902 385520
rect 503958 385464 503963 385520
rect 501860 385462 503963 385464
rect 503897 385459 503963 385462
rect 502057 385250 502123 385253
rect 502014 385248 502123 385250
rect 502014 385192 502062 385248
rect 502118 385192 502123 385248
rect 502014 385187 502123 385192
rect 502014 385116 502074 385187
rect 502006 385052 502012 385116
rect 502076 385052 502082 385116
rect 78673 383890 78739 383893
rect 78673 383888 82156 383890
rect 78673 383832 78678 383888
rect 78734 383832 82156 383888
rect 78673 383830 82156 383832
rect 78673 383827 78739 383830
rect 67030 383556 67036 383620
rect 67100 383556 67106 383620
rect 67038 383485 67098 383556
rect 66989 383480 67098 383485
rect 66989 383424 66994 383480
rect 67050 383424 67098 383480
rect 66989 383422 67098 383424
rect 66989 383419 67055 383422
rect 503897 381986 503963 381989
rect 501860 381984 503963 381986
rect 501860 381928 503902 381984
rect 503958 381928 503963 381984
rect 501860 381926 503963 381928
rect 503897 381923 503963 381926
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 81709 380354 81775 380357
rect 81709 380352 82156 380354
rect 81709 380296 81714 380352
rect 81770 380296 82156 380352
rect 81709 380294 82156 380296
rect 81709 380291 81775 380294
rect 503897 378178 503963 378181
rect 501860 378176 503963 378178
rect 501860 378120 503902 378176
rect 503958 378120 503963 378176
rect 501860 378118 503963 378120
rect 503897 378115 503963 378118
rect 82486 377028 82492 377092
rect 82556 377028 82562 377092
rect 82494 376788 82554 377028
rect 522205 376820 522271 376821
rect 522205 376818 522252 376820
rect 522160 376816 522252 376818
rect 522160 376760 522210 376816
rect 522160 376758 522252 376760
rect 522205 376756 522252 376758
rect 522316 376756 522322 376820
rect 522205 376755 522271 376756
rect 503897 374642 503963 374645
rect 501860 374640 503963 374642
rect 501860 374584 503902 374640
rect 503958 374584 503963 374640
rect 501860 374582 503963 374584
rect 503897 374579 503963 374582
rect 66989 374098 67055 374101
rect 67214 374098 67220 374100
rect 66989 374096 67220 374098
rect 66989 374040 66994 374096
rect 67050 374040 67220 374096
rect 66989 374038 67220 374040
rect 66989 374035 67055 374038
rect 67214 374036 67220 374038
rect 67284 374036 67290 374100
rect 66846 373764 66852 373828
rect 66916 373826 66922 373828
rect 67214 373826 67220 373828
rect 66916 373766 67220 373826
rect 66916 373764 66922 373766
rect 67214 373764 67220 373766
rect 67284 373764 67290 373828
rect 81750 372948 81756 373012
rect 81820 373010 81826 373012
rect 81820 372950 82156 373010
rect 81820 372948 81826 372950
rect 503897 371106 503963 371109
rect 501860 371104 503963 371106
rect 501860 371048 503902 371104
rect 503958 371048 503963 371104
rect 501860 371046 503963 371048
rect 503897 371043 503963 371046
rect 522246 370018 522252 370020
rect 522070 369958 522252 370018
rect 522070 369748 522130 369958
rect 522246 369956 522252 369958
rect 522316 369956 522322 370020
rect 522062 369684 522068 369748
rect 522132 369684 522138 369748
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 78673 369474 78739 369477
rect 78673 369472 82156 369474
rect 78673 369416 78678 369472
rect 78734 369416 82156 369472
rect 583520 369460 584960 369550
rect 78673 369414 82156 369416
rect 78673 369411 78739 369414
rect 503989 367298 504055 367301
rect 501860 367296 504055 367298
rect 501860 367240 503994 367296
rect 504050 367240 504055 367296
rect 501860 367238 504055 367240
rect 503989 367235 504055 367238
rect -960 366210 480 366300
rect -960 366150 674 366210
rect -960 366060 480 366150
rect 614 365802 674 366150
rect 71078 365802 71084 365804
rect 614 365742 71084 365802
rect 71078 365740 71084 365742
rect 71148 365740 71154 365804
rect 78070 365604 78076 365668
rect 78140 365666 78146 365668
rect 78140 365606 82156 365666
rect 78140 365604 78146 365606
rect 503989 363762 504055 363765
rect 501860 363760 504055 363762
rect 501860 363704 503994 363760
rect 504050 363704 504055 363760
rect 501860 363702 504055 363704
rect 503989 363699 504055 363702
rect 78673 362130 78739 362133
rect 78673 362128 82156 362130
rect 78673 362072 78678 362128
rect 78734 362072 82156 362128
rect 78673 362070 82156 362072
rect 78673 362067 78739 362070
rect 501822 360844 501828 360908
rect 501892 360906 501898 360908
rect 502057 360906 502123 360909
rect 501892 360904 502123 360906
rect 501892 360848 502062 360904
rect 502118 360848 502123 360904
rect 501892 360846 502123 360848
rect 501892 360844 501898 360846
rect 502057 360843 502123 360846
rect 503989 359954 504055 359957
rect 501860 359952 504055 359954
rect 501860 359896 503994 359952
rect 504050 359896 504055 359952
rect 501860 359894 504055 359896
rect 503989 359891 504055 359894
rect 78673 358322 78739 358325
rect 78673 358320 82156 358322
rect 78673 358264 78678 358320
rect 78734 358264 82156 358320
rect 78673 358262 82156 358264
rect 78673 358259 78739 358262
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect 521878 357308 521884 357372
rect 521948 357370 521954 357372
rect 522205 357370 522271 357373
rect 521948 357368 522271 357370
rect 521948 357312 522210 357368
rect 522266 357312 522271 357368
rect 521948 357310 522271 357312
rect 521948 357308 521954 357310
rect 522205 357307 522271 357310
rect 505277 356418 505343 356421
rect 501860 356416 505343 356418
rect 501860 356360 505282 356416
rect 505338 356360 505343 356416
rect 501860 356358 505343 356360
rect 505277 356355 505343 356358
rect 502057 356146 502123 356149
rect 502190 356146 502196 356148
rect 502057 356144 502196 356146
rect 502057 356088 502062 356144
rect 502118 356088 502196 356144
rect 502057 356086 502196 356088
rect 502057 356083 502123 356086
rect 502190 356084 502196 356086
rect 502260 356084 502266 356148
rect 502241 354652 502307 354653
rect 502190 354588 502196 354652
rect 502260 354650 502307 354652
rect 502260 354648 502352 354650
rect 502302 354592 502352 354648
rect 502260 354590 502352 354592
rect 502260 354588 502307 354590
rect 502241 354587 502307 354588
rect 502609 352610 502675 352613
rect 501860 352608 502675 352610
rect 501860 352552 502614 352608
rect 502670 352552 502675 352608
rect 501860 352550 502675 352552
rect 502609 352547 502675 352550
rect -960 351780 480 352020
rect 78673 351250 78739 351253
rect 78673 351248 82156 351250
rect 78673 351192 78678 351248
rect 78734 351192 82156 351248
rect 78673 351190 82156 351192
rect 78673 351187 78739 351190
rect 67214 350706 67220 350708
rect 66854 350646 67220 350706
rect 66854 350572 66914 350646
rect 67214 350644 67220 350646
rect 67284 350644 67290 350708
rect 66846 350508 66852 350572
rect 66916 350508 66922 350572
rect 521694 350508 521700 350572
rect 521764 350570 521770 350572
rect 522205 350570 522271 350573
rect 521764 350568 522271 350570
rect 521764 350512 522210 350568
rect 522266 350512 522271 350568
rect 521764 350510 522271 350512
rect 521764 350508 521770 350510
rect 522205 350507 522271 350510
rect 501646 348532 501706 349044
rect 501638 348468 501644 348532
rect 501708 348468 501714 348532
rect 521694 347652 521700 347716
rect 521764 347652 521770 347716
rect 521702 347578 521762 347652
rect 522205 347578 522271 347581
rect 521702 347576 522271 347578
rect 521702 347520 522210 347576
rect 522266 347520 522271 347576
rect 521702 347518 522271 347520
rect 522205 347515 522271 347518
rect 78673 347442 78739 347445
rect 78673 347440 82156 347442
rect 78673 347384 78678 347440
rect 78734 347384 82156 347440
rect 78673 347382 82156 347384
rect 78673 347379 78739 347382
rect 580257 346082 580323 346085
rect 583520 346082 584960 346172
rect 580257 346080 584960 346082
rect 580257 346024 580262 346080
rect 580318 346024 584960 346080
rect 580257 346022 584960 346024
rect 580257 346019 580323 346022
rect 583520 345932 584960 346022
rect 504081 345538 504147 345541
rect 501860 345536 504147 345538
rect 501860 345480 504086 345536
rect 504142 345480 504147 345536
rect 501860 345478 504147 345480
rect 504081 345475 504147 345478
rect 502241 345266 502307 345269
rect 502198 345264 502307 345266
rect 502198 345208 502246 345264
rect 502302 345208 502307 345264
rect 502198 345203 502307 345208
rect 502198 345132 502258 345203
rect 502190 345068 502196 345132
rect 502260 345068 502266 345132
rect 79777 343906 79843 343909
rect 79777 343904 82156 343906
rect 79777 343848 79782 343904
rect 79838 343848 82156 343904
rect 79777 343846 82156 343848
rect 79777 343843 79843 343846
rect 504081 341730 504147 341733
rect 501860 341728 504147 341730
rect 501860 341672 504086 341728
rect 504142 341672 504147 341728
rect 501860 341670 504147 341672
rect 504081 341667 504147 341670
rect 66846 340988 66852 341052
rect 66916 340988 66922 341052
rect 66854 340778 66914 340988
rect 67030 340778 67036 340780
rect 66854 340718 67036 340778
rect 67030 340716 67036 340718
rect 67100 340716 67106 340780
rect 80881 340098 80947 340101
rect 80881 340096 82156 340098
rect 80881 340040 80886 340096
rect 80942 340040 82156 340096
rect 80881 340038 82156 340040
rect 80881 340035 80947 340038
rect 502190 339690 502196 339692
rect 502014 339630 502196 339690
rect 502014 339420 502074 339630
rect 502190 339628 502196 339630
rect 502260 339628 502266 339692
rect 502006 339356 502012 339420
rect 502076 339356 502082 339420
rect 504081 338194 504147 338197
rect 501860 338192 504147 338194
rect 501860 338136 504086 338192
rect 504142 338136 504147 338192
rect 501860 338134 504147 338136
rect 504081 338131 504147 338134
rect 521878 338132 521884 338196
rect 521948 338194 521954 338196
rect 522205 338194 522271 338197
rect 521948 338192 522271 338194
rect 521948 338136 522210 338192
rect 522266 338136 522271 338192
rect 521948 338134 522271 338136
rect 521948 338132 521954 338134
rect 522205 338131 522271 338134
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 67030 336636 67036 336700
rect 67100 336636 67106 336700
rect 66713 336562 66779 336565
rect 67038 336562 67098 336636
rect 66713 336560 67098 336562
rect 66713 336504 66718 336560
rect 66774 336504 67098 336560
rect 66713 336502 67098 336504
rect 78673 336562 78739 336565
rect 78673 336560 82156 336562
rect 78673 336504 78678 336560
rect 78734 336504 82156 336560
rect 78673 336502 82156 336504
rect 66713 336499 66779 336502
rect 78673 336499 78739 336502
rect 502057 335340 502123 335341
rect 502006 335338 502012 335340
rect 501966 335278 502012 335338
rect 502076 335336 502123 335340
rect 502118 335280 502123 335336
rect 502006 335276 502012 335278
rect 502076 335276 502123 335280
rect 502057 335275 502123 335276
rect 504081 334386 504147 334389
rect 501860 334384 504147 334386
rect 501860 334328 504086 334384
rect 504142 334328 504147 334384
rect 501860 334326 504147 334328
rect 504081 334323 504147 334326
rect 583520 334236 584960 334476
rect 78673 332754 78739 332757
rect 78673 332752 82156 332754
rect 78673 332696 78678 332752
rect 78734 332696 82156 332752
rect 78673 332694 82156 332696
rect 78673 332691 78739 332694
rect 521878 331332 521884 331396
rect 521948 331332 521954 331396
rect 521886 331122 521946 331332
rect 522062 331122 522068 331124
rect 521886 331062 522068 331122
rect 522062 331060 522068 331062
rect 522132 331060 522138 331124
rect 505369 330850 505435 330853
rect 501860 330848 505435 330850
rect 501860 330792 505374 330848
rect 505430 330792 505435 330848
rect 501860 330790 505435 330792
rect 505369 330787 505435 330790
rect 78673 329218 78739 329221
rect 78673 329216 82156 329218
rect 78673 329160 78678 329216
rect 78734 329160 82156 329216
rect 78673 329158 82156 329160
rect 78673 329155 78739 329158
rect 66897 328402 66963 328405
rect 67398 328402 67404 328404
rect 66897 328400 67404 328402
rect 66897 328344 66902 328400
rect 66958 328344 67404 328400
rect 66897 328342 67404 328344
rect 66897 328339 66963 328342
rect 67398 328340 67404 328342
rect 67468 328340 67474 328404
rect 522062 328340 522068 328404
rect 522132 328402 522138 328404
rect 522205 328402 522271 328405
rect 522132 328400 522271 328402
rect 522132 328344 522210 328400
rect 522266 328344 522271 328400
rect 522132 328342 522271 328344
rect 522132 328340 522138 328342
rect 522205 328339 522271 328342
rect 501689 327586 501755 327589
rect 501646 327584 501755 327586
rect 501646 327528 501694 327584
rect 501750 327528 501755 327584
rect 501646 327523 501755 327528
rect 66713 327314 66779 327317
rect 66670 327312 66779 327314
rect 66670 327256 66718 327312
rect 66774 327256 66779 327312
rect 66670 327251 66779 327256
rect 66670 327180 66730 327251
rect 66662 327116 66668 327180
rect 66732 327116 66738 327180
rect 501646 327012 501706 327523
rect 502057 325818 502123 325821
rect 502190 325818 502196 325820
rect 502057 325816 502196 325818
rect 502057 325760 502062 325816
rect 502118 325760 502196 325816
rect 502057 325758 502196 325760
rect 502057 325755 502123 325758
rect 502190 325756 502196 325758
rect 502260 325756 502266 325820
rect 78673 325682 78739 325685
rect 78673 325680 82156 325682
rect 78673 325624 78678 325680
rect 78734 325624 82156 325680
rect 78673 325622 82156 325624
rect 78673 325619 78739 325622
rect 66897 323642 66963 323645
rect 67398 323642 67404 323644
rect 66897 323640 67404 323642
rect 66897 323584 66902 323640
rect 66958 323584 67404 323640
rect 66897 323582 67404 323584
rect 66897 323579 66963 323582
rect 67398 323580 67404 323582
rect 67468 323580 67474 323644
rect 504081 323506 504147 323509
rect 501860 323504 504147 323506
rect 501860 323448 504086 323504
rect 504142 323448 504147 323504
rect 501860 323446 504147 323448
rect 504081 323443 504147 323446
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 78673 321874 78739 321877
rect 78673 321872 82156 321874
rect 78673 321816 78678 321872
rect 78734 321816 82156 321872
rect 78673 321814 82156 321816
rect 78673 321811 78739 321814
rect 501454 321676 501460 321740
rect 501524 321676 501530 321740
rect 501462 321466 501522 321676
rect 501597 321466 501663 321469
rect 501462 321464 501663 321466
rect 501462 321408 501602 321464
rect 501658 321408 501663 321464
rect 501462 321406 501663 321408
rect 501597 321403 501663 321406
rect 504081 319970 504147 319973
rect 501860 319968 504147 319970
rect 501860 319912 504086 319968
rect 504142 319912 504147 319968
rect 501860 319910 504147 319912
rect 504081 319907 504147 319910
rect 522205 319018 522271 319021
rect 521886 319016 522271 319018
rect 521886 318960 522210 319016
rect 522266 318960 522271 319016
rect 521886 318958 522271 318960
rect 521886 318884 521946 318958
rect 522205 318955 522271 318958
rect 521878 318820 521884 318884
rect 521948 318820 521954 318884
rect 78673 318338 78739 318341
rect 78673 318336 82156 318338
rect 78673 318280 78678 318336
rect 78734 318280 82156 318336
rect 78673 318278 82156 318280
rect 78673 318275 78739 318278
rect 504081 316162 504147 316165
rect 501860 316160 504147 316162
rect 501860 316104 504086 316160
rect 504142 316104 504147 316160
rect 501860 316102 504147 316104
rect 504081 316099 504147 316102
rect 81617 314530 81683 314533
rect 81617 314528 82156 314530
rect 81617 314472 81622 314528
rect 81678 314472 82156 314528
rect 81617 314470 82156 314472
rect 81617 314467 81683 314470
rect 502425 312626 502491 312629
rect 501860 312624 502491 312626
rect 501860 312568 502430 312624
rect 502486 312568 502491 312624
rect 501860 312566 502491 312568
rect 502425 312563 502491 312566
rect 67030 312082 67036 312084
rect 66854 312022 67036 312082
rect 66854 311812 66914 312022
rect 67030 312020 67036 312022
rect 67100 312020 67106 312084
rect 501597 312082 501663 312085
rect 501462 312080 501663 312082
rect 501462 312024 501602 312080
rect 501658 312024 501663 312080
rect 501462 312022 501663 312024
rect 501462 311948 501522 312022
rect 501597 312019 501663 312022
rect 521878 312020 521884 312084
rect 521948 312020 521954 312084
rect 501454 311884 501460 311948
rect 501524 311884 501530 311948
rect 66846 311748 66852 311812
rect 66916 311748 66922 311812
rect 521886 311810 521946 312020
rect 522062 311810 522068 311812
rect 521886 311750 522068 311810
rect 522062 311748 522068 311750
rect 522132 311748 522138 311812
rect 78673 310994 78739 310997
rect 78673 310992 82156 310994
rect 78673 310936 78678 310992
rect 78734 310936 82156 310992
rect 78673 310934 82156 310936
rect 78673 310931 78739 310934
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 522062 309028 522068 309092
rect 522132 309028 522138 309092
rect 522070 308954 522130 309028
rect 522205 308954 522271 308957
rect 522070 308952 522271 308954
rect -960 308818 480 308908
rect 522070 308896 522210 308952
rect 522266 308896 522271 308952
rect 522070 308894 522271 308896
rect 522205 308891 522271 308894
rect 3417 308818 3483 308821
rect -960 308816 3483 308818
rect -960 308760 3422 308816
rect 3478 308760 3483 308816
rect -960 308758 3483 308760
rect -960 308668 480 308758
rect 3417 308755 3483 308758
rect 501646 308277 501706 308788
rect 501597 308272 501706 308277
rect 501597 308216 501602 308272
rect 501658 308216 501706 308272
rect 501597 308214 501706 308216
rect 501597 308211 501663 308214
rect 78213 307186 78279 307189
rect 78213 307184 82156 307186
rect 78213 307128 78218 307184
rect 78274 307128 82156 307184
rect 78213 307126 82156 307128
rect 78213 307123 78279 307126
rect 504081 305282 504147 305285
rect 501860 305280 504147 305282
rect 501860 305224 504086 305280
rect 504142 305224 504147 305280
rect 501860 305222 504147 305224
rect 504081 305219 504147 305222
rect 78121 303650 78187 303653
rect 78121 303648 82156 303650
rect 78121 303592 78126 303648
rect 78182 303592 82156 303648
rect 78121 303590 82156 303592
rect 78121 303587 78187 303590
rect 66662 302228 66668 302292
rect 66732 302228 66738 302292
rect 66670 302154 66730 302228
rect 66846 302154 66852 302156
rect 66670 302094 66852 302154
rect 66846 302092 66852 302094
rect 66916 302092 66922 302156
rect 521878 302092 521884 302156
rect 521948 302154 521954 302156
rect 522205 302154 522271 302157
rect 521948 302152 522271 302154
rect 521948 302096 522210 302152
rect 522266 302096 522271 302152
rect 521948 302094 522271 302096
rect 521948 302092 521954 302094
rect 522205 302091 522271 302094
rect 505461 301474 505527 301477
rect 501860 301472 505527 301474
rect 501860 301416 505466 301472
rect 505522 301416 505527 301472
rect 501860 301414 505527 301416
rect 505461 301411 505527 301414
rect 79225 300114 79291 300117
rect 79225 300112 82156 300114
rect 79225 300056 79230 300112
rect 79286 300056 82156 300112
rect 79225 300054 82156 300056
rect 79225 300051 79291 300054
rect 67030 299372 67036 299436
rect 67100 299372 67106 299436
rect 67038 299301 67098 299372
rect 66989 299296 67098 299301
rect 66989 299240 66994 299296
rect 67050 299240 67098 299296
rect 66989 299238 67098 299240
rect 66989 299235 67055 299238
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 504030 297938 504036 297940
rect 501860 297878 504036 297938
rect 504030 297876 504036 297878
rect 504100 297876 504106 297940
rect 78673 296306 78739 296309
rect 78673 296304 82156 296306
rect 78673 296248 78678 296304
rect 78734 296248 82156 296304
rect 78673 296246 82156 296248
rect 78673 296243 78739 296246
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect 504081 294402 504147 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect 501860 294400 504147 294402
rect 501860 294344 504086 294400
rect 504142 294344 504147 294400
rect 501860 294342 504147 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 504081 294339 504147 294342
rect 78673 292770 78739 292773
rect 78673 292768 82156 292770
rect 78673 292712 78678 292768
rect 78734 292712 82156 292768
rect 78673 292710 82156 292712
rect 78673 292707 78739 292710
rect 504081 290594 504147 290597
rect 501860 290592 504147 290594
rect 501860 290536 504086 290592
rect 504142 290536 504147 290592
rect 501860 290534 504147 290536
rect 504081 290531 504147 290534
rect 66989 290050 67055 290053
rect 66989 290048 67098 290050
rect 66989 289992 66994 290048
rect 67050 289992 67098 290048
rect 66989 289987 67098 289992
rect 67038 289916 67098 289987
rect 67030 289852 67036 289916
rect 67100 289852 67106 289916
rect 522062 289716 522068 289780
rect 522132 289716 522138 289780
rect 522070 289642 522130 289716
rect 522205 289642 522271 289645
rect 522070 289640 522271 289642
rect 522070 289584 522210 289640
rect 522266 289584 522271 289640
rect 522070 289582 522271 289584
rect 522205 289579 522271 289582
rect 69974 288492 69980 288556
rect 70044 288554 70050 288556
rect 82126 288554 82186 288932
rect 70044 288494 82186 288554
rect 70044 288492 70050 288494
rect 583520 287316 584960 287556
rect 504081 287058 504147 287061
rect 501860 287056 504147 287058
rect 501860 287000 504086 287056
rect 504142 287000 504147 287056
rect 501860 286998 504147 287000
rect 504081 286995 504147 286998
rect 82494 284884 82554 285396
rect 82486 284820 82492 284884
rect 82556 284820 82562 284884
rect 504030 283324 504036 283388
rect 504100 283386 504106 283388
rect 504173 283386 504239 283389
rect 504100 283384 504239 283386
rect 504100 283328 504178 283384
rect 504234 283328 504239 283384
rect 504100 283326 504239 283328
rect 504100 283324 504106 283326
rect 504173 283323 504239 283326
rect 504081 283250 504147 283253
rect 501860 283248 504147 283250
rect 501860 283192 504086 283248
rect 504142 283192 504147 283248
rect 501860 283190 504147 283192
rect 504081 283187 504147 283190
rect 78673 281618 78739 281621
rect 78673 281616 82156 281618
rect 78673 281560 78678 281616
rect 78734 281560 82156 281616
rect 78673 281558 82156 281560
rect 78673 281555 78739 281558
rect 504173 280394 504239 280397
rect 522205 280394 522271 280397
rect 504038 280392 504239 280394
rect 504038 280336 504178 280392
rect 504234 280336 504239 280392
rect 504038 280334 504239 280336
rect 504038 280260 504098 280334
rect 504173 280331 504239 280334
rect 521886 280392 522271 280394
rect 521886 280336 522210 280392
rect 522266 280336 522271 280392
rect 521886 280334 522271 280336
rect 521886 280260 521946 280334
rect 522205 280331 522271 280334
rect -960 280122 480 280212
rect 504030 280196 504036 280260
rect 504100 280196 504106 280260
rect 521878 280196 521884 280260
rect 521948 280196 521954 280260
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 66897 280122 66963 280125
rect 67030 280122 67036 280124
rect 66897 280120 67036 280122
rect 66897 280064 66902 280120
rect 66958 280064 67036 280120
rect 66897 280062 67036 280064
rect 66897 280059 66963 280062
rect 67030 280060 67036 280062
rect 67100 280060 67106 280124
rect 501830 279173 501890 279684
rect 501781 279168 501890 279173
rect 501781 279112 501786 279168
rect 501842 279112 501890 279168
rect 501781 279110 501890 279112
rect 501781 279107 501847 279110
rect 3417 278898 3483 278901
rect 21214 278898 21220 278900
rect 3417 278896 21220 278898
rect 3417 278840 3422 278896
rect 3478 278840 21220 278896
rect 3417 278838 21220 278840
rect 3417 278835 3483 278838
rect 21214 278836 21220 278838
rect 21284 278836 21290 278900
rect 512821 278762 512887 278765
rect 513005 278762 513071 278765
rect 512821 278760 513071 278762
rect 512821 278704 512826 278760
rect 512882 278704 513010 278760
rect 513066 278704 513071 278760
rect 512821 278702 513071 278704
rect 512821 278699 512887 278702
rect 513005 278699 513071 278702
rect 78673 278082 78739 278085
rect 78673 278080 82156 278082
rect 78673 278024 78678 278080
rect 78734 278024 82156 278080
rect 78673 278022 82156 278024
rect 78673 278019 78739 278022
rect 504081 275906 504147 275909
rect 501860 275904 504147 275906
rect 501860 275848 504086 275904
rect 504142 275848 504147 275904
rect 501860 275846 504147 275848
rect 504081 275843 504147 275846
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 78673 274546 78739 274549
rect 78673 274544 82156 274546
rect 78673 274488 78678 274544
rect 78734 274488 82156 274544
rect 78673 274486 82156 274488
rect 78673 274483 78739 274486
rect 521878 273396 521884 273460
rect 521948 273396 521954 273460
rect 521886 273050 521946 273396
rect 522062 273050 522068 273052
rect 521886 272990 522068 273050
rect 522062 272988 522068 272990
rect 522132 272988 522138 273052
rect 501646 271965 501706 272340
rect 501646 271960 501755 271965
rect 501646 271904 501694 271960
rect 501750 271904 501755 271960
rect 501646 271902 501755 271904
rect 501689 271899 501755 271902
rect 66897 270738 66963 270741
rect 66854 270736 66963 270738
rect 66854 270680 66902 270736
rect 66958 270680 66963 270736
rect 66854 270675 66963 270680
rect 81617 270738 81683 270741
rect 81617 270736 82156 270738
rect 81617 270680 81622 270736
rect 81678 270680 82156 270736
rect 81617 270678 82156 270680
rect 81617 270675 81683 270678
rect 66854 270604 66914 270675
rect 66846 270540 66852 270604
rect 66916 270540 66922 270604
rect 522062 270404 522068 270468
rect 522132 270466 522138 270468
rect 522205 270466 522271 270469
rect 522132 270464 522271 270466
rect 522132 270408 522210 270464
rect 522266 270408 522271 270464
rect 522132 270406 522271 270408
rect 522132 270404 522138 270406
rect 522205 270403 522271 270406
rect 501822 269180 501828 269244
rect 501892 269242 501898 269244
rect 502006 269242 502012 269244
rect 501892 269182 502012 269242
rect 501892 269180 501898 269182
rect 502006 269180 502012 269182
rect 502076 269180 502082 269244
rect 504081 268834 504147 268837
rect 501860 268832 504147 268834
rect 501860 268776 504086 268832
rect 504142 268776 504147 268832
rect 501860 268774 504147 268776
rect 504081 268771 504147 268774
rect 78673 267202 78739 267205
rect 78673 267200 82156 267202
rect 78673 267144 78678 267200
rect 78734 267144 82156 267200
rect 78673 267142 82156 267144
rect 78673 267139 78739 267142
rect -960 265706 480 265796
rect 3417 265706 3483 265709
rect -960 265704 3483 265706
rect -960 265648 3422 265704
rect 3478 265648 3483 265704
rect -960 265646 3483 265648
rect -960 265556 480 265646
rect 3417 265643 3483 265646
rect 502701 265026 502767 265029
rect 501860 265024 502767 265026
rect 501860 264968 502706 265024
rect 502762 264968 502767 265024
rect 501860 264966 502767 264968
rect 502701 264963 502767 264966
rect 583520 263938 584960 264028
rect 538262 263878 547890 263938
rect 529054 263604 529060 263668
rect 529124 263666 529130 263668
rect 538262 263666 538322 263878
rect 547830 263802 547890 263878
rect 557582 263878 567210 263938
rect 547830 263742 557458 263802
rect 529124 263606 538322 263666
rect 557398 263666 557458 263742
rect 557582 263666 557642 263878
rect 567150 263802 567210 263878
rect 583342 263878 584960 263938
rect 567150 263742 576778 263802
rect 557398 263606 557642 263666
rect 576718 263666 576778 263742
rect 583342 263666 583402 263878
rect 583520 263788 584960 263878
rect 576718 263606 583402 263666
rect 529124 263604 529130 263606
rect 78673 263394 78739 263397
rect 78673 263392 82156 263394
rect 78673 263336 78678 263392
rect 78734 263336 82156 263392
rect 78673 263334 82156 263336
rect 78673 263331 78739 263334
rect 504081 261490 504147 261493
rect 501860 261488 504147 261490
rect 501860 261432 504086 261488
rect 504142 261432 504147 261488
rect 501860 261430 504147 261432
rect 504081 261427 504147 261430
rect 522205 261082 522271 261085
rect 521886 261080 522271 261082
rect 521886 261024 522210 261080
rect 522266 261024 522271 261080
rect 521886 261022 522271 261024
rect 521886 260948 521946 261022
rect 522205 261019 522271 261022
rect 521878 260884 521884 260948
rect 521948 260884 521954 260948
rect 66662 260748 66668 260812
rect 66732 260810 66738 260812
rect 67030 260810 67036 260812
rect 66732 260750 67036 260810
rect 66732 260748 66738 260750
rect 67030 260748 67036 260750
rect 67100 260748 67106 260812
rect 79685 259858 79751 259861
rect 79685 259856 82156 259858
rect 79685 259800 79690 259856
rect 79746 259800 82156 259856
rect 79685 259798 82156 259800
rect 79685 259795 79751 259798
rect 512821 259450 512887 259453
rect 513005 259450 513071 259453
rect 512821 259448 513071 259450
rect 512821 259392 512826 259448
rect 512882 259392 513010 259448
rect 513066 259392 513071 259448
rect 512821 259390 513071 259392
rect 512821 259387 512887 259390
rect 513005 259387 513071 259390
rect 504081 257682 504147 257685
rect 501860 257680 504147 257682
rect 501860 257624 504086 257680
rect 504142 257624 504147 257680
rect 501860 257622 504147 257624
rect 504081 257619 504147 257622
rect 81014 255988 81020 256052
rect 81084 256050 81090 256052
rect 81084 255990 82156 256050
rect 81084 255988 81090 255990
rect 501270 255988 501276 256052
rect 501340 256050 501346 256052
rect 501454 256050 501460 256052
rect 501340 255990 501460 256050
rect 501340 255988 501346 255990
rect 501454 255988 501460 255990
rect 501524 255988 501530 256052
rect 503621 254418 503687 254421
rect 504030 254418 504036 254420
rect 503621 254416 504036 254418
rect 503621 254360 503626 254416
rect 503682 254360 504036 254416
rect 503621 254358 504036 254360
rect 503621 254355 503687 254358
rect 504030 254356 504036 254358
rect 504100 254356 504106 254420
rect 505553 254146 505619 254149
rect 501860 254144 505619 254146
rect 501860 254088 505558 254144
rect 505614 254088 505619 254144
rect 501860 254086 505619 254088
rect 505553 254083 505619 254086
rect 521878 253948 521884 254012
rect 521948 253948 521954 254012
rect 503621 253876 503687 253877
rect 503621 253872 503668 253876
rect 503732 253874 503738 253876
rect 503621 253816 503626 253872
rect 503621 253812 503668 253816
rect 503732 253814 503778 253874
rect 503732 253812 503738 253814
rect 503621 253811 503687 253812
rect 521886 253738 521946 253948
rect 522062 253738 522068 253740
rect 521886 253678 522068 253738
rect 522062 253676 522068 253678
rect 522132 253676 522138 253740
rect 78673 252514 78739 252517
rect 78673 252512 82156 252514
rect 78673 252456 78678 252512
rect 78734 252456 82156 252512
rect 78673 252454 82156 252456
rect 78673 252451 78739 252454
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 67214 251092 67220 251156
rect 67284 251092 67290 251156
rect 522062 251092 522068 251156
rect 522132 251154 522138 251156
rect 522205 251154 522271 251157
rect 522132 251152 522271 251154
rect 522132 251096 522210 251152
rect 522266 251096 522271 251152
rect 522132 251094 522271 251096
rect 522132 251092 522138 251094
rect 67030 250956 67036 251020
rect 67100 251018 67106 251020
rect 67222 251018 67282 251092
rect 522205 251091 522271 251094
rect 67100 250958 67282 251018
rect 67100 250956 67106 250958
rect 504081 250338 504147 250341
rect 501860 250336 504147 250338
rect 501860 250280 504086 250336
rect 504142 250280 504147 250336
rect 501860 250278 504147 250280
rect 504081 250275 504147 250278
rect 78673 248978 78739 248981
rect 78673 248976 82156 248978
rect 78673 248920 78678 248976
rect 78734 248920 82156 248976
rect 78673 248918 82156 248920
rect 78673 248915 78739 248918
rect 504081 246802 504147 246805
rect 501860 246800 504147 246802
rect 501860 246744 504086 246800
rect 504142 246744 504147 246800
rect 501860 246742 504147 246744
rect 504081 246739 504147 246742
rect 79358 245108 79364 245172
rect 79428 245170 79434 245172
rect 79428 245110 82156 245170
rect 79428 245108 79434 245110
rect 504081 243266 504147 243269
rect 501860 243264 504147 243266
rect 501860 243208 504086 243264
rect 504142 243208 504147 243264
rect 501860 243206 504147 243208
rect 504081 243203 504147 243206
rect 67398 242042 67404 242044
rect 67222 241982 67404 242042
rect 67222 241634 67282 241982
rect 67398 241980 67404 241982
rect 67468 241980 67474 242044
rect 522205 241770 522271 241773
rect 521886 241768 522271 241770
rect 521886 241712 522210 241768
rect 522266 241712 522271 241768
rect 521886 241710 522271 241712
rect 67398 241634 67404 241636
rect 67222 241574 67404 241634
rect 67398 241572 67404 241574
rect 67468 241572 67474 241636
rect 78673 241634 78739 241637
rect 521886 241636 521946 241710
rect 522205 241707 522271 241710
rect 78673 241632 82156 241634
rect 78673 241576 78678 241632
rect 78734 241576 82156 241632
rect 78673 241574 82156 241576
rect 78673 241571 78739 241574
rect 521878 241572 521884 241636
rect 521948 241572 521954 241636
rect 583520 240396 584960 240636
rect 67081 240138 67147 240141
rect 67214 240138 67220 240140
rect 67081 240136 67220 240138
rect 67081 240080 67086 240136
rect 67142 240080 67220 240136
rect 67081 240078 67220 240080
rect 67081 240075 67147 240078
rect 67214 240076 67220 240078
rect 67284 240076 67290 240140
rect 512821 240138 512887 240141
rect 513005 240138 513071 240141
rect 512821 240136 513071 240138
rect 512821 240080 512826 240136
rect 512882 240080 513010 240136
rect 513066 240080 513071 240136
rect 512821 240078 513071 240080
rect 512821 240075 512887 240078
rect 513005 240075 513071 240078
rect 501830 238914 501890 239428
rect 502006 238914 502012 238916
rect 501830 238854 502012 238914
rect 502006 238852 502012 238854
rect 502076 238852 502082 238916
rect 78673 237826 78739 237829
rect 78673 237824 82156 237826
rect 78673 237768 78678 237824
rect 78734 237768 82156 237824
rect 78673 237766 82156 237768
rect 78673 237763 78739 237766
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 504081 235922 504147 235925
rect 501860 235920 504147 235922
rect 501860 235864 504086 235920
rect 504142 235864 504147 235920
rect 501860 235862 504147 235864
rect 504081 235859 504147 235862
rect 521878 234636 521884 234700
rect 521948 234636 521954 234700
rect 521886 234426 521946 234636
rect 522062 234426 522068 234428
rect 521886 234366 522068 234426
rect 522062 234364 522068 234366
rect 522132 234364 522138 234428
rect 78673 234290 78739 234293
rect 78673 234288 82156 234290
rect 78673 234232 78678 234288
rect 78734 234232 82156 234288
rect 78673 234230 82156 234232
rect 78673 234227 78739 234230
rect 503662 232188 503668 232252
rect 503732 232250 503738 232252
rect 503732 232190 504282 232250
rect 503732 232188 503738 232190
rect 504081 232114 504147 232117
rect 501860 232112 504147 232114
rect 501860 232056 504086 232112
rect 504142 232056 504147 232112
rect 501860 232054 504147 232056
rect 504081 232051 504147 232054
rect 503846 231814 503852 231878
rect 503916 231876 503922 231878
rect 504222 231876 504282 232190
rect 503916 231816 504282 231876
rect 503916 231814 503922 231816
rect 78673 230482 78739 230485
rect 78673 230480 82156 230482
rect 78673 230424 78678 230480
rect 78734 230424 82156 230480
rect 78673 230422 82156 230424
rect 78673 230419 78739 230422
rect 501454 229196 501460 229260
rect 501524 229196 501530 229260
rect 501462 228988 501522 229196
rect 501454 228924 501460 228988
rect 501524 228924 501530 228988
rect 501638 228788 501644 228852
rect 501708 228850 501714 228852
rect 501965 228850 502031 228853
rect 501708 228848 502031 228850
rect 501708 228792 501970 228848
rect 502026 228792 502031 228848
rect 501708 228790 502031 228792
rect 501708 228788 501714 228790
rect 501965 228787 502031 228790
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 504081 228578 504147 228581
rect 501860 228576 504147 228578
rect 501860 228520 504086 228576
rect 504142 228520 504147 228576
rect 501860 228518 504147 228520
rect 504081 228515 504147 228518
rect 501822 228108 501828 228172
rect 501892 228170 501898 228172
rect 507158 228170 507164 228172
rect 501892 228110 507164 228170
rect 501892 228108 501898 228110
rect 507158 228108 507164 228110
rect 507228 228108 507234 228172
rect 82486 227428 82492 227492
rect 82556 227428 82562 227492
rect 511574 227428 511580 227492
rect 511644 227490 511650 227492
rect 522246 227490 522252 227492
rect 511644 227430 522252 227490
rect 511644 227428 511650 227430
rect 522246 227428 522252 227430
rect 522316 227428 522322 227492
rect 82494 226916 82554 227428
rect 504081 224770 504147 224773
rect 501860 224768 504147 224770
rect 501860 224712 504086 224768
rect 504142 224712 504147 224768
rect 501860 224710 504147 224712
rect 504081 224707 504147 224710
rect 78673 223410 78739 223413
rect 78673 223408 82156 223410
rect 78673 223352 78678 223408
rect 78734 223352 82156 223408
rect 78673 223350 82156 223352
rect 78673 223347 78739 223350
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 67081 222458 67147 222461
rect 67038 222456 67147 222458
rect 67038 222400 67086 222456
rect 67142 222400 67147 222456
rect 67038 222395 67147 222400
rect 67038 222324 67098 222395
rect 67030 222260 67036 222324
rect 67100 222260 67106 222324
rect 521878 222124 521884 222188
rect 521948 222186 521954 222188
rect 522205 222186 522271 222189
rect 521948 222184 522271 222186
rect 521948 222128 522210 222184
rect 522266 222128 522271 222184
rect 521948 222126 522271 222128
rect 521948 222124 521954 222126
rect 522205 222123 522271 222126
rect 504081 221234 504147 221237
rect 501860 221232 504147 221234
rect 501860 221176 504086 221232
rect 504142 221176 504147 221232
rect 501860 221174 504147 221176
rect 504081 221171 504147 221174
rect 501965 220962 502031 220965
rect 501965 220960 502074 220962
rect 501822 220866 501828 220930
rect 501892 220928 501898 220930
rect 501965 220928 501970 220960
rect 501892 220904 501970 220928
rect 502026 220904 502074 220960
rect 501892 220868 502074 220904
rect 501892 220866 501898 220868
rect 512821 220826 512887 220829
rect 513005 220826 513071 220829
rect 512821 220824 513071 220826
rect 512821 220768 512826 220824
rect 512882 220768 513010 220824
rect 513066 220768 513071 220824
rect 512821 220766 513071 220768
rect 512821 220763 512887 220766
rect 513005 220763 513071 220766
rect 79593 219602 79659 219605
rect 79593 219600 82156 219602
rect 79593 219544 79598 219600
rect 79654 219544 82156 219600
rect 79593 219542 82156 219544
rect 79593 219539 79659 219542
rect 501270 219540 501276 219604
rect 501340 219602 501346 219604
rect 501340 219542 501522 219602
rect 501340 219540 501346 219542
rect 501462 219468 501522 219542
rect 501454 219404 501460 219468
rect 501524 219404 501530 219468
rect 502885 217698 502951 217701
rect 501860 217696 502951 217698
rect 501860 217640 502890 217696
rect 502946 217640 502951 217696
rect 501860 217638 502951 217640
rect 502885 217635 502951 217638
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 81709 216066 81775 216069
rect 81709 216064 82156 216066
rect 81709 216008 81714 216064
rect 81770 216008 82156 216064
rect 81709 216006 82156 216008
rect 81709 216003 81775 216006
rect 67030 215522 67036 215524
rect 66854 215462 67036 215522
rect 66854 215252 66914 215462
rect 67030 215460 67036 215462
rect 67100 215460 67106 215524
rect 66846 215188 66852 215252
rect 66916 215188 66922 215252
rect 504081 213890 504147 213893
rect 501860 213888 504147 213890
rect 501860 213832 504086 213888
rect 504142 213832 504147 213888
rect 501860 213830 504147 213832
rect 504081 213827 504147 213830
rect 522062 212604 522068 212668
rect 522132 212666 522138 212668
rect 522205 212666 522271 212669
rect 522132 212664 522271 212666
rect 522132 212608 522210 212664
rect 522266 212608 522271 212664
rect 522132 212606 522271 212608
rect 522132 212604 522138 212606
rect 522205 212603 522271 212606
rect 522062 212468 522068 212532
rect 522132 212530 522138 212532
rect 522205 212530 522271 212533
rect 522132 212528 522271 212530
rect 522132 212472 522210 212528
rect 522266 212472 522271 212528
rect 522132 212470 522271 212472
rect 522132 212468 522138 212470
rect 522205 212467 522271 212470
rect 78673 212258 78739 212261
rect 78673 212256 82156 212258
rect 78673 212200 78678 212256
rect 78734 212200 82156 212256
rect 78673 212198 82156 212200
rect 78673 212195 78739 212198
rect 512821 211170 512887 211173
rect 513005 211170 513071 211173
rect 512821 211168 513071 211170
rect 512821 211112 512826 211168
rect 512882 211112 513010 211168
rect 513066 211112 513071 211168
rect 512821 211110 513071 211112
rect 512821 211107 512887 211110
rect 513005 211107 513071 211110
rect 504081 210354 504147 210357
rect 501860 210352 504147 210354
rect 501860 210296 504086 210352
rect 504142 210296 504147 210352
rect 501860 210294 504147 210296
rect 504081 210291 504147 210294
rect 78673 208722 78739 208725
rect 78673 208720 82156 208722
rect 78673 208664 78678 208720
rect 78734 208664 82156 208720
rect 78673 208662 82156 208664
rect 78673 208659 78739 208662
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 501822 206892 501828 206956
rect 501892 206892 501898 206956
rect 501830 206818 501890 206892
rect 502006 206818 502012 206820
rect 501830 206758 502012 206818
rect 502006 206756 502012 206758
rect 502076 206756 502082 206820
rect 67081 206002 67147 206005
rect 67398 206002 67404 206004
rect 67081 206000 67404 206002
rect 67081 205944 67086 206000
rect 67142 205944 67404 206000
rect 67081 205942 67404 205944
rect 67081 205939 67147 205942
rect 67398 205940 67404 205942
rect 67468 205940 67474 206004
rect 76465 206002 76531 206005
rect 77150 206002 77156 206004
rect 76465 206000 77156 206002
rect 76465 205944 76470 206000
rect 76526 205944 77156 206000
rect 76465 205942 77156 205944
rect 76465 205939 76531 205942
rect 77150 205940 77156 205942
rect 77220 205940 77226 206004
rect 501462 205732 501522 206516
rect 521878 206212 521884 206276
rect 521948 206274 521954 206276
rect 522205 206274 522271 206277
rect 521948 206272 522271 206274
rect 521948 206216 522210 206272
rect 522266 206216 522271 206272
rect 521948 206214 522271 206216
rect 521948 206212 521954 206214
rect 522205 206211 522271 206214
rect 61326 205668 61332 205732
rect 61396 205730 61402 205732
rect 75862 205730 75868 205732
rect 61396 205670 75868 205730
rect 61396 205668 61402 205670
rect 75862 205668 75868 205670
rect 75932 205668 75938 205732
rect 501454 205668 501460 205732
rect 501524 205668 501530 205732
rect 70158 205532 70164 205596
rect 70228 205594 70234 205596
rect 70228 205534 82186 205594
rect 70228 205532 70234 205534
rect 67081 205458 67147 205461
rect 67398 205458 67404 205460
rect 67081 205456 67404 205458
rect 67081 205400 67086 205456
rect 67142 205400 67404 205456
rect 67081 205398 67404 205400
rect 67081 205395 67147 205398
rect 67398 205396 67404 205398
rect 67468 205396 67474 205460
rect 76465 205458 76531 205461
rect 77150 205458 77156 205460
rect 76465 205456 77156 205458
rect 76465 205400 76470 205456
rect 76526 205400 77156 205456
rect 76465 205398 77156 205400
rect 76465 205395 76531 205398
rect 77150 205396 77156 205398
rect 77220 205396 77226 205460
rect 75862 204988 75868 205052
rect 75932 205050 75938 205052
rect 78990 205050 78996 205052
rect 75932 204990 78996 205050
rect 75932 204988 75938 204990
rect 78990 204988 78996 204990
rect 79060 204988 79066 205052
rect 82126 204884 82186 205534
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect 504081 203010 504147 203013
rect 501860 203008 504147 203010
rect 501860 202952 504086 203008
rect 504142 202952 504147 203008
rect 501860 202950 504147 202952
rect 504081 202947 504147 202950
rect 66713 201380 66779 201381
rect 66662 201316 66668 201380
rect 66732 201378 66779 201380
rect 80789 201378 80855 201381
rect 66732 201376 66824 201378
rect 66774 201320 66824 201376
rect 66732 201318 66824 201320
rect 80789 201376 82156 201378
rect 80789 201320 80794 201376
rect 80850 201320 82156 201376
rect 80789 201318 82156 201320
rect 66732 201316 66779 201318
rect 66713 201315 66779 201316
rect 80789 201315 80855 201318
rect 521561 200018 521627 200021
rect 521878 200018 521884 200020
rect 521561 200016 521884 200018
rect 521561 199960 521566 200016
rect 521622 199960 521884 200016
rect 521561 199958 521884 199960
rect 521561 199955 521627 199958
rect 521878 199956 521884 199958
rect 521948 199956 521954 200020
rect 501462 198932 501522 199172
rect 501454 198868 501460 198932
rect 501524 198868 501530 198932
rect 77937 197842 78003 197845
rect 77937 197840 82156 197842
rect 77937 197784 77942 197840
rect 77998 197784 82156 197840
rect 77937 197782 82156 197784
rect 77937 197779 78003 197782
rect 504173 195666 504239 195669
rect 501860 195664 504239 195666
rect 501860 195608 504178 195664
rect 504234 195608 504239 195664
rect 501860 195606 504239 195608
rect 504173 195603 504239 195606
rect 66478 195468 66484 195532
rect 66548 195530 66554 195532
rect 66713 195530 66779 195533
rect 66548 195528 66779 195530
rect 66548 195472 66718 195528
rect 66774 195472 66779 195528
rect 66548 195470 66779 195472
rect 66548 195468 66554 195470
rect 66713 195467 66779 195470
rect 503846 194516 503852 194580
rect 503916 194516 503922 194580
rect 503854 194442 503914 194516
rect 504265 194442 504331 194445
rect 503854 194440 504331 194442
rect 503854 194384 504270 194440
rect 504326 194384 504331 194440
rect 503854 194382 504331 194384
rect 504265 194379 504331 194382
rect 78673 194034 78739 194037
rect 78673 194032 82156 194034
rect -960 193898 480 193988
rect 78673 193976 78678 194032
rect 78734 193976 82156 194032
rect 78673 193974 82156 193976
rect 78673 193971 78739 193974
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 504030 192130 504036 192132
rect 501860 192070 504036 192130
rect 504030 192068 504036 192070
rect 504100 192068 504106 192132
rect 512821 191858 512887 191861
rect 513005 191858 513071 191861
rect 512821 191856 513071 191858
rect 512821 191800 512826 191856
rect 512882 191800 513010 191856
rect 513066 191800 513071 191856
rect 512821 191798 513071 191800
rect 512821 191795 512887 191798
rect 513005 191795 513071 191798
rect 66478 191660 66484 191724
rect 66548 191660 66554 191724
rect 66486 191586 66546 191660
rect 67081 191586 67147 191589
rect 66486 191584 67147 191586
rect 66486 191528 67086 191584
rect 67142 191528 67147 191584
rect 66486 191526 67147 191528
rect 67081 191523 67147 191526
rect 72325 190498 72391 190501
rect 73061 190498 73127 190501
rect 72325 190496 73127 190498
rect 72325 190440 72330 190496
rect 72386 190440 73066 190496
rect 73122 190440 73127 190496
rect 72325 190438 73127 190440
rect 72325 190435 72391 190438
rect 73061 190435 73127 190438
rect 78673 190498 78739 190501
rect 521561 190498 521627 190501
rect 521694 190498 521700 190500
rect 78673 190496 82156 190498
rect 78673 190440 78678 190496
rect 78734 190440 82156 190496
rect 78673 190438 82156 190440
rect 521561 190496 521700 190498
rect 521561 190440 521566 190496
rect 521622 190440 521700 190496
rect 521561 190438 521700 190440
rect 78673 190435 78739 190438
rect 521561 190435 521627 190438
rect 521694 190436 521700 190438
rect 521764 190436 521770 190500
rect 504173 188322 504239 188325
rect 501860 188320 504239 188322
rect 501860 188264 504178 188320
rect 504234 188264 504239 188320
rect 501860 188262 504239 188264
rect 504173 188259 504239 188262
rect 75494 187716 75500 187780
rect 75564 187778 75570 187780
rect 79409 187778 79475 187781
rect 75564 187776 79475 187778
rect 75564 187720 79414 187776
rect 79470 187720 79475 187776
rect 75564 187718 79475 187720
rect 75564 187716 75570 187718
rect 79409 187715 79475 187718
rect 502006 187716 502012 187780
rect 502076 187716 502082 187780
rect 502014 187506 502074 187716
rect 502190 187506 502196 187508
rect 502014 187446 502196 187506
rect 502190 187444 502196 187446
rect 502260 187444 502266 187508
rect 79225 186690 79291 186693
rect 79225 186688 82156 186690
rect 79225 186632 79230 186688
rect 79286 186632 82156 186688
rect 79225 186630 82156 186632
rect 79225 186627 79291 186630
rect 504265 186284 504331 186285
rect 504214 186220 504220 186284
rect 504284 186282 504331 186284
rect 504284 186280 504376 186282
rect 504326 186224 504376 186280
rect 504284 186222 504376 186224
rect 504284 186220 504331 186222
rect 504265 186219 504331 186220
rect 504265 185332 504331 185333
rect 504214 185330 504220 185332
rect 504174 185270 504220 185330
rect 504284 185328 504331 185332
rect 504326 185272 504331 185328
rect 504214 185268 504220 185270
rect 504284 185268 504331 185272
rect 504265 185267 504331 185268
rect 504173 185194 504239 185197
rect 503854 185192 504239 185194
rect 503854 185136 504178 185192
rect 504234 185136 504239 185192
rect 503854 185134 504239 185136
rect 503854 185060 503914 185134
rect 504173 185131 504239 185134
rect 503846 184996 503852 185060
rect 503916 184996 503922 185060
rect 504265 184786 504331 184789
rect 501860 184784 504331 184786
rect 501860 184728 504270 184784
rect 504326 184728 504331 184784
rect 501860 184726 504331 184728
rect 504265 184723 504331 184726
rect 501454 183908 501460 183972
rect 501524 183970 501530 183972
rect 501873 183970 501939 183973
rect 501524 183968 501939 183970
rect 501524 183912 501878 183968
rect 501934 183912 501939 183968
rect 501524 183910 501939 183912
rect 501524 183908 501530 183910
rect 501873 183907 501939 183910
rect 78673 183154 78739 183157
rect 78673 183152 82156 183154
rect 78673 183096 78678 183152
rect 78734 183096 82156 183152
rect 78673 183094 82156 183096
rect 78673 183091 78739 183094
rect 501822 182820 501828 182884
rect 501892 182882 501898 182884
rect 502190 182882 502196 182884
rect 501892 182822 502196 182882
rect 501892 182820 501898 182822
rect 502190 182820 502196 182822
rect 502260 182820 502266 182884
rect 583520 181930 584960 182020
rect 583342 181870 584960 181930
rect 531262 181324 531268 181388
rect 531332 181386 531338 181388
rect 540881 181386 540947 181389
rect 531332 181384 540947 181386
rect 531332 181328 540886 181384
rect 540942 181328 540947 181384
rect 531332 181326 540947 181328
rect 531332 181324 531338 181326
rect 540881 181323 540947 181326
rect 503294 181188 503300 181252
rect 503364 181250 503370 181252
rect 503805 181250 503871 181253
rect 503364 181248 503871 181250
rect 503364 181192 503810 181248
rect 503866 181192 503871 181248
rect 503364 181190 503871 181192
rect 503364 181188 503370 181190
rect 503805 181187 503871 181190
rect 522246 181052 522252 181116
rect 522316 181114 522322 181116
rect 540881 181114 540947 181117
rect 583342 181114 583402 181870
rect 583520 181780 584960 181870
rect 522316 181054 524522 181114
rect 522316 181052 522322 181054
rect 505645 180978 505711 180981
rect 501860 180976 505711 180978
rect 501860 180920 505650 180976
rect 505706 180920 505711 180976
rect 501860 180918 505711 180920
rect 524462 180978 524522 181054
rect 540881 181112 553410 181114
rect 540881 181056 540886 181112
rect 540942 181056 553410 181112
rect 540881 181054 553410 181056
rect 540881 181051 540947 181054
rect 531262 180978 531268 180980
rect 524462 180918 531268 180978
rect 505645 180915 505711 180918
rect 531262 180916 531268 180918
rect 531332 180916 531338 180980
rect 553350 180978 553410 181054
rect 572670 181054 583402 181114
rect 553350 180918 562978 180978
rect 562918 180842 562978 180918
rect 572670 180842 572730 181054
rect 562918 180782 572730 180842
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 78673 179346 78739 179349
rect 78673 179344 82156 179346
rect 78673 179288 78678 179344
rect 78734 179288 82156 179344
rect 78673 179286 82156 179288
rect 78673 179283 78739 179286
rect 503805 177442 503871 177445
rect 501860 177440 503871 177442
rect 501860 177384 503810 177440
rect 503866 177384 503871 177440
rect 501860 177382 503871 177384
rect 503805 177379 503871 177382
rect 521878 176762 521884 176764
rect 521702 176702 521884 176762
rect 504173 176628 504239 176629
rect 504173 176626 504220 176628
rect 504128 176624 504220 176626
rect 504128 176568 504178 176624
rect 504128 176566 504220 176568
rect 504173 176564 504220 176566
rect 504284 176564 504290 176628
rect 504173 176563 504239 176564
rect 521702 176492 521762 176702
rect 521878 176700 521884 176702
rect 521948 176700 521954 176764
rect 521694 176428 521700 176492
rect 521764 176428 521770 176492
rect 82678 175405 82738 175780
rect 82629 175400 82738 175405
rect 504173 175404 504239 175405
rect 504173 175402 504220 175404
rect 82629 175344 82634 175400
rect 82690 175344 82738 175400
rect 82629 175342 82738 175344
rect 504128 175400 504220 175402
rect 504128 175344 504178 175400
rect 504128 175342 504220 175344
rect 82629 175339 82695 175342
rect 504173 175340 504220 175342
rect 504284 175340 504290 175404
rect 504173 175339 504239 175340
rect 503846 175204 503852 175268
rect 503916 175204 503922 175268
rect 503854 175130 503914 175204
rect 504357 175130 504423 175133
rect 503854 175128 504423 175130
rect 503854 175072 504362 175128
rect 504418 175072 504423 175128
rect 503854 175070 504423 175072
rect 504357 175067 504423 175070
rect 67081 174178 67147 174181
rect 67081 174176 67282 174178
rect 67081 174120 67086 174176
rect 67142 174120 67282 174176
rect 67081 174118 67282 174120
rect 67081 174115 67147 174118
rect 67222 174044 67282 174118
rect 503713 174044 503779 174045
rect 67214 173980 67220 174044
rect 67284 173980 67290 174044
rect 503662 174042 503668 174044
rect 503622 173982 503668 174042
rect 503732 174040 503779 174044
rect 503774 173984 503779 174040
rect 503662 173980 503668 173982
rect 503732 173980 503779 173984
rect 503713 173979 503779 173980
rect 521694 173844 521700 173908
rect 521764 173906 521770 173908
rect 522205 173906 522271 173909
rect 521764 173904 522271 173906
rect 521764 173848 522210 173904
rect 522266 173848 522271 173904
rect 521764 173846 522271 173848
rect 521764 173844 521770 173846
rect 522205 173843 522271 173846
rect 504173 173634 504239 173637
rect 501860 173632 504239 173634
rect 501860 173576 504178 173632
rect 504234 173576 504239 173632
rect 501860 173574 504239 173576
rect 504173 173571 504239 173574
rect 512821 172546 512887 172549
rect 513005 172546 513071 172549
rect 512821 172544 513071 172546
rect 512821 172488 512826 172544
rect 512882 172488 513010 172544
rect 513066 172488 513071 172544
rect 512821 172486 513071 172488
rect 512821 172483 512887 172486
rect 513005 172483 513071 172486
rect 78673 172274 78739 172277
rect 78673 172272 82156 172274
rect 78673 172216 78678 172272
rect 78734 172216 82156 172272
rect 78673 172214 82156 172216
rect 78673 172211 78739 172214
rect 503713 170098 503779 170101
rect 501860 170096 503779 170098
rect 501860 170040 503718 170096
rect 503774 170040 503779 170096
rect 501860 170038 503779 170040
rect 503713 170035 503779 170038
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 81801 168466 81867 168469
rect 81801 168464 82156 168466
rect 81801 168408 81806 168464
rect 81862 168408 82156 168464
rect 81801 168406 82156 168408
rect 81801 168403 81867 168406
rect 503713 166562 503779 166565
rect 501860 166560 503779 166562
rect 501860 166504 503718 166560
rect 503774 166504 503779 166560
rect 501860 166502 503779 166504
rect 503713 166499 503779 166502
rect 504357 165882 504423 165885
rect 503716 165880 504423 165882
rect 503716 165824 504362 165880
rect 504418 165824 504423 165880
rect 503716 165822 504423 165824
rect 503716 165644 503776 165822
rect 504357 165819 504423 165822
rect 503846 165644 503852 165646
rect 503716 165584 503852 165644
rect 503846 165582 503852 165584
rect 503916 165582 503922 165646
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 78673 164930 78739 164933
rect 78673 164928 82156 164930
rect 78673 164872 78678 164928
rect 78734 164872 82156 164928
rect 78673 164870 82156 164872
rect 78673 164867 78739 164870
rect 521878 164188 521884 164252
rect 521948 164250 521954 164252
rect 522205 164250 522271 164253
rect 521948 164248 522271 164250
rect 521948 164192 522210 164248
rect 522266 164192 522271 164248
rect 521948 164190 522271 164192
rect 521948 164188 521954 164190
rect 522205 164187 522271 164190
rect 504449 162754 504515 162757
rect 501860 162752 504515 162754
rect 501860 162696 504454 162752
rect 504510 162696 504515 162752
rect 501860 162694 504515 162696
rect 504449 162691 504515 162694
rect 78029 161122 78095 161125
rect 78029 161120 82156 161122
rect 78029 161064 78034 161120
rect 78090 161064 82156 161120
rect 78029 161062 82156 161064
rect 78029 161059 78095 161062
rect 502793 159218 502859 159221
rect 501860 159216 502859 159218
rect 501860 159160 502798 159216
rect 502854 159160 502859 159216
rect 501860 159158 502859 159160
rect 502793 159155 502859 159158
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 78673 157586 78739 157589
rect 78673 157584 82156 157586
rect 78673 157528 78678 157584
rect 78734 157528 82156 157584
rect 78673 157526 82156 157528
rect 78673 157523 78739 157526
rect 521878 157450 521884 157452
rect 521702 157390 521884 157450
rect 521702 157180 521762 157390
rect 521878 157388 521884 157390
rect 521948 157388 521954 157452
rect 521694 157116 521700 157180
rect 521764 157116 521770 157180
rect 72182 155212 72188 155276
rect 72252 155274 72258 155276
rect 82077 155274 82143 155277
rect 72252 155272 82143 155274
rect 72252 155216 82082 155272
rect 82138 155216 82143 155272
rect 72252 155214 82143 155216
rect 72252 155212 72258 155214
rect 82077 155211 82143 155214
rect 501462 154868 501522 155380
rect 501454 154804 501460 154868
rect 501524 154804 501530 154868
rect 78673 153778 78739 153781
rect 78673 153776 82156 153778
rect 78673 153720 78678 153776
rect 78734 153720 82156 153776
rect 78673 153718 82156 153720
rect 78673 153715 78739 153718
rect 503713 151874 503779 151877
rect 501860 151872 503779 151874
rect 501860 151816 503718 151872
rect 503774 151816 503779 151872
rect 501860 151814 503779 151816
rect 503713 151811 503779 151814
rect 501454 151132 501460 151196
rect 501524 151194 501530 151196
rect 503989 151194 504055 151197
rect 501524 151192 504055 151194
rect 501524 151136 503994 151192
rect 504050 151136 504055 151192
rect 501524 151134 504055 151136
rect 501524 151132 501530 151134
rect 503989 151131 504055 151134
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 78673 150242 78739 150245
rect 78673 150240 82156 150242
rect 78673 150184 78678 150240
rect 78734 150184 82156 150240
rect 78673 150182 82156 150184
rect 78673 150179 78739 150182
rect 503713 148066 503779 148069
rect 501860 148064 503779 148066
rect 501860 148008 503718 148064
rect 503774 148008 503779 148064
rect 501860 148006 503779 148008
rect 503713 148003 503779 148006
rect 521694 147596 521700 147660
rect 521764 147658 521770 147660
rect 522430 147658 522436 147660
rect 521764 147598 522436 147658
rect 521764 147596 521770 147598
rect 522430 147596 522436 147598
rect 522500 147596 522506 147660
rect 78673 146706 78739 146709
rect 78673 146704 82156 146706
rect 78673 146648 78678 146704
rect 78734 146648 82156 146704
rect 78673 146646 82156 146648
rect 78673 146643 78739 146646
rect 583520 146556 584960 146796
rect 66662 144876 66668 144940
rect 66732 144938 66738 144940
rect 66846 144938 66852 144940
rect 66732 144878 66852 144938
rect 66732 144876 66738 144878
rect 66846 144876 66852 144878
rect 66916 144876 66922 144940
rect 504541 144530 504607 144533
rect 501860 144528 504607 144530
rect 501860 144472 504546 144528
rect 504602 144472 504607 144528
rect 501860 144470 504607 144472
rect 504541 144467 504607 144470
rect 79501 142898 79567 142901
rect 79501 142896 82156 142898
rect 79501 142840 79506 142896
rect 79562 142840 82156 142896
rect 79501 142838 82156 142840
rect 79501 142835 79567 142838
rect 504541 140994 504607 140997
rect 501860 140992 504607 140994
rect 501860 140936 504546 140992
rect 504602 140936 504607 140992
rect 501860 140934 504607 140936
rect 504541 140931 504607 140934
rect 82494 138821 82554 139332
rect 82494 138816 82603 138821
rect 82494 138760 82542 138816
rect 82598 138760 82603 138816
rect 82494 138758 82603 138760
rect 82537 138755 82603 138758
rect 522430 138138 522436 138140
rect 522254 138078 522436 138138
rect 66662 137804 66668 137868
rect 66732 137866 66738 137868
rect 67214 137866 67220 137868
rect 66732 137806 67220 137866
rect 66732 137804 66738 137806
rect 67214 137804 67220 137806
rect 67284 137804 67290 137868
rect 501505 137866 501571 137869
rect 522254 137868 522314 138078
rect 522430 138076 522436 138078
rect 522500 138076 522506 138140
rect 501638 137866 501644 137868
rect 501505 137864 501644 137866
rect 501505 137808 501510 137864
rect 501566 137808 501644 137864
rect 501505 137806 501644 137808
rect 501505 137803 501571 137806
rect 501638 137804 501644 137806
rect 501708 137804 501714 137868
rect 522246 137804 522252 137868
rect 522316 137804 522322 137868
rect 501462 136645 501522 137156
rect 501462 136640 501571 136645
rect 501462 136584 501510 136640
rect 501566 136584 501571 136640
rect 501462 136582 501571 136584
rect 501505 136579 501571 136582
rect -960 136370 480 136460
rect 3509 136370 3575 136373
rect -960 136368 3575 136370
rect -960 136312 3514 136368
rect 3570 136312 3575 136368
rect -960 136310 3575 136312
rect -960 136220 480 136310
rect 3509 136307 3575 136310
rect 82678 135013 82738 135524
rect 522297 135148 522363 135149
rect 522246 135084 522252 135148
rect 522316 135146 522363 135148
rect 522316 135144 522408 135146
rect 522358 135088 522408 135144
rect 522316 135086 522408 135088
rect 522316 135084 522363 135086
rect 522297 135083 522363 135084
rect 82629 135008 82738 135013
rect 82629 134952 82634 135008
rect 82690 134952 82738 135008
rect 82629 134950 82738 134952
rect 82629 134947 82695 134950
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 503069 133650 503135 133653
rect 501860 133648 503135 133650
rect 501860 133592 503074 133648
rect 503130 133592 503135 133648
rect 501860 133590 503135 133592
rect 503069 133587 503135 133590
rect 78673 132018 78739 132021
rect 78673 132016 82156 132018
rect 78673 131960 78678 132016
rect 78734 131960 82156 132016
rect 78673 131958 82156 131960
rect 78673 131955 78739 131958
rect 505737 129842 505803 129845
rect 501860 129840 505803 129842
rect 501860 129784 505742 129840
rect 505798 129784 505803 129840
rect 501860 129782 505803 129784
rect 505737 129779 505803 129782
rect 78673 128210 78739 128213
rect 78673 128208 82156 128210
rect 78673 128152 78678 128208
rect 78734 128152 82156 128208
rect 78673 128150 82156 128152
rect 78673 128147 78739 128150
rect 501454 126924 501460 126988
rect 501524 126986 501530 126988
rect 501965 126986 502031 126989
rect 501524 126984 502031 126986
rect 501524 126928 501970 126984
rect 502026 126928 502031 126984
rect 501524 126926 502031 126928
rect 501524 126924 501530 126926
rect 501965 126923 502031 126926
rect 504541 126306 504607 126309
rect 501860 126304 504607 126306
rect 501860 126248 504546 126304
rect 504602 126248 504607 126304
rect 501860 126246 504607 126248
rect 504541 126243 504607 126246
rect 521878 125564 521884 125628
rect 521948 125626 521954 125628
rect 522297 125626 522363 125629
rect 521948 125624 522363 125626
rect 521948 125568 522302 125624
rect 522358 125568 522363 125624
rect 521948 125566 522363 125568
rect 521948 125564 521954 125566
rect 522297 125563 522363 125566
rect 79409 124674 79475 124677
rect 79409 124672 82156 124674
rect 79409 124616 79414 124672
rect 79470 124616 82156 124672
rect 79409 124614 82156 124616
rect 79409 124611 79475 124614
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect 501873 122770 501939 122773
rect 502006 122770 502012 122772
rect 501873 122768 502012 122770
rect 501873 122712 501878 122768
rect 501934 122712 502012 122768
rect 501873 122710 502012 122712
rect 501873 122707 501939 122710
rect 502006 122708 502012 122710
rect 502076 122708 502082 122772
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 501830 121957 501890 122468
rect 501830 121952 501939 121957
rect 501830 121896 501878 121952
rect 501934 121896 501939 121952
rect 501830 121894 501939 121896
rect 501873 121891 501939 121894
rect 501454 121484 501460 121548
rect 501524 121546 501530 121548
rect 501524 121486 501706 121546
rect 501524 121484 501530 121486
rect 501646 121276 501706 121486
rect 501638 121212 501644 121276
rect 501708 121212 501714 121276
rect 82126 120597 82186 121108
rect 82126 120592 82235 120597
rect 82126 120536 82174 120592
rect 82230 120536 82235 120592
rect 82126 120534 82235 120536
rect 82169 120531 82235 120534
rect 501454 119308 501460 119372
rect 501524 119370 501530 119372
rect 501965 119370 502031 119373
rect 501524 119368 502031 119370
rect 501524 119312 501970 119368
rect 502026 119312 502031 119368
rect 501524 119310 502031 119312
rect 501524 119308 501530 119310
rect 501965 119307 502031 119310
rect 503989 118962 504055 118965
rect 501860 118960 504055 118962
rect 501860 118904 503994 118960
rect 504050 118904 504055 118960
rect 501860 118902 504055 118904
rect 503989 118899 504055 118902
rect 521878 118764 521884 118828
rect 521948 118764 521954 118828
rect 521886 118554 521946 118764
rect 522062 118554 522068 118556
rect 521886 118494 522068 118554
rect 522062 118492 522068 118494
rect 522132 118492 522138 118556
rect 81985 117058 82051 117061
rect 82126 117058 82186 117300
rect 81985 117056 82186 117058
rect 81985 117000 81990 117056
rect 82046 117000 82186 117056
rect 81985 116998 82186 117000
rect 81985 116995 82051 116998
rect 522062 115772 522068 115836
rect 522132 115834 522138 115836
rect 522205 115834 522271 115837
rect 522132 115832 522271 115834
rect 522132 115776 522210 115832
rect 522266 115776 522271 115832
rect 522132 115774 522271 115776
rect 522132 115772 522138 115774
rect 522205 115771 522271 115774
rect 501830 114882 501890 115396
rect 501830 114822 502074 114882
rect 502014 114610 502074 114822
rect 512678 114610 512684 114612
rect 502014 114550 512684 114610
rect 512678 114548 512684 114550
rect 512748 114548 512754 114612
rect 67081 114476 67147 114477
rect 67030 114412 67036 114476
rect 67100 114474 67147 114476
rect 67100 114472 67192 114474
rect 67142 114416 67192 114472
rect 67100 114414 67192 114416
rect 67100 114412 67147 114414
rect 67081 114411 67147 114412
rect 79133 113794 79199 113797
rect 79133 113792 82156 113794
rect 79133 113736 79138 113792
rect 79194 113736 82156 113792
rect 79133 113734 82156 113736
rect 79133 113731 79199 113734
rect 67081 113386 67147 113389
rect 67038 113384 67147 113386
rect 67038 113328 67086 113384
rect 67142 113328 67147 113384
rect 67038 113323 67147 113328
rect 67038 113252 67098 113323
rect 67030 113188 67036 113252
rect 67100 113188 67106 113252
rect 503253 111618 503319 111621
rect 501860 111616 503319 111618
rect 501860 111560 503258 111616
rect 503314 111560 503319 111616
rect 501860 111558 503319 111560
rect 503253 111555 503319 111558
rect 580257 111482 580323 111485
rect 583520 111482 584960 111572
rect 580257 111480 584960 111482
rect 580257 111424 580262 111480
rect 580318 111424 584960 111480
rect 580257 111422 584960 111424
rect 580257 111419 580323 111422
rect 583520 111332 584960 111422
rect 78673 109986 78739 109989
rect 78673 109984 82156 109986
rect 78673 109928 78678 109984
rect 78734 109928 82156 109984
rect 78673 109926 82156 109928
rect 78673 109923 78739 109926
rect 503345 108082 503411 108085
rect 501860 108080 503411 108082
rect 501860 108024 503350 108080
rect 503406 108024 503411 108080
rect 501860 108022 503411 108024
rect 503345 108019 503411 108022
rect -960 107674 480 107764
rect 4061 107674 4127 107677
rect -960 107672 4127 107674
rect -960 107616 4066 107672
rect 4122 107616 4127 107672
rect -960 107614 4127 107616
rect -960 107524 480 107614
rect 4061 107611 4127 107614
rect 82629 106722 82695 106725
rect 82629 106720 82738 106722
rect 82629 106664 82634 106720
rect 82690 106664 82738 106720
rect 82629 106659 82738 106664
rect 82678 106420 82738 106659
rect 521878 106252 521884 106316
rect 521948 106314 521954 106316
rect 522205 106314 522271 106317
rect 521948 106312 522271 106314
rect 521948 106256 522210 106312
rect 522266 106256 522271 106312
rect 521948 106254 522271 106256
rect 521948 106252 521954 106254
rect 522205 106251 522271 106254
rect 504541 104274 504607 104277
rect 501860 104272 504607 104274
rect 501860 104216 504546 104272
rect 504602 104216 504607 104272
rect 501860 104214 504607 104216
rect 504541 104211 504607 104214
rect 67030 103396 67036 103460
rect 67100 103396 67106 103460
rect 67038 103325 67098 103396
rect 67038 103320 67147 103325
rect 67038 103264 67086 103320
rect 67142 103264 67147 103320
rect 67038 103262 67147 103264
rect 67081 103259 67147 103262
rect 75177 102778 75243 102781
rect 502374 102778 502380 102780
rect 75177 102776 108314 102778
rect 75177 102720 75182 102776
rect 75238 102720 108314 102776
rect 75177 102718 108314 102720
rect 75177 102715 75243 102718
rect 108254 102642 108314 102718
rect 118742 102718 124322 102778
rect 108941 102642 109007 102645
rect 108254 102640 109007 102642
rect 108254 102584 108946 102640
rect 109002 102584 109007 102640
rect 108254 102582 109007 102584
rect 108941 102579 109007 102582
rect 109125 102642 109191 102645
rect 118417 102642 118483 102645
rect 109125 102640 118483 102642
rect 109125 102584 109130 102640
rect 109186 102584 118422 102640
rect 118478 102584 118483 102640
rect 109125 102582 118483 102584
rect 109125 102579 109191 102582
rect 118417 102579 118483 102582
rect 118601 102642 118667 102645
rect 118742 102642 118802 102718
rect 118601 102640 118802 102642
rect 118601 102584 118606 102640
rect 118662 102584 118802 102640
rect 118601 102582 118802 102584
rect 124262 102642 124322 102718
rect 138614 102718 144930 102778
rect 125501 102642 125567 102645
rect 124262 102640 125567 102642
rect 124262 102584 125506 102640
rect 125562 102584 125567 102640
rect 124262 102582 125567 102584
rect 118601 102579 118667 102582
rect 125501 102579 125567 102582
rect 133689 102642 133755 102645
rect 133873 102642 133939 102645
rect 133689 102640 133939 102642
rect 133689 102584 133694 102640
rect 133750 102584 133878 102640
rect 133934 102584 133939 102640
rect 133689 102582 133939 102584
rect 133689 102579 133755 102582
rect 133873 102579 133939 102582
rect 82854 102444 82860 102508
rect 82924 102506 82930 102508
rect 84009 102506 84075 102509
rect 82924 102504 84075 102506
rect 82924 102448 84014 102504
rect 84070 102448 84075 102504
rect 82924 102446 84075 102448
rect 82924 102444 82930 102446
rect 84009 102443 84075 102446
rect 133965 102506 134031 102509
rect 138614 102506 138674 102718
rect 144870 102644 144930 102718
rect 154622 102718 166826 102778
rect 144862 102580 144868 102644
rect 144932 102580 144938 102644
rect 154622 102642 154682 102718
rect 154438 102582 154682 102642
rect 166766 102608 166826 102718
rect 274590 102718 502380 102778
rect 176745 102642 176811 102645
rect 167134 102640 176811 102642
rect 167134 102608 176750 102640
rect 166766 102584 176750 102608
rect 176806 102584 176811 102640
rect 166766 102582 176811 102584
rect 133965 102504 138674 102506
rect 133965 102448 133970 102504
rect 134026 102448 138674 102504
rect 133965 102446 138674 102448
rect 133965 102443 134031 102446
rect 144862 102308 144868 102372
rect 144932 102370 144938 102372
rect 154438 102370 154498 102582
rect 166766 102548 167194 102582
rect 176745 102579 176811 102582
rect 274590 102509 274650 102718
rect 502374 102716 502380 102718
rect 502444 102716 502450 102780
rect 307661 102642 307727 102645
rect 497774 102642 497780 102644
rect 307661 102640 497780 102642
rect 307661 102584 307666 102640
rect 307722 102584 497780 102640
rect 307661 102582 497780 102584
rect 307661 102579 307727 102582
rect 497774 102580 497780 102582
rect 497844 102580 497850 102644
rect 500902 102580 500908 102644
rect 500972 102642 500978 102644
rect 501270 102642 501276 102644
rect 500972 102582 501276 102642
rect 500972 102580 500978 102582
rect 501270 102580 501276 102582
rect 501340 102580 501346 102644
rect 274541 102504 274650 102509
rect 274541 102448 274546 102504
rect 274602 102448 274650 102504
rect 274541 102446 274650 102448
rect 274541 102443 274607 102446
rect 492806 102444 492812 102508
rect 492876 102444 492882 102508
rect 493726 102506 493732 102508
rect 492998 102446 493732 102506
rect 144932 102310 154498 102370
rect 144932 102308 144938 102310
rect 483013 102234 483079 102237
rect 492814 102236 492874 102444
rect 492998 102372 493058 102446
rect 493726 102444 493732 102446
rect 493796 102444 493802 102508
rect 492990 102308 492996 102372
rect 493060 102308 493066 102372
rect 499982 102308 499988 102372
rect 500052 102370 500058 102372
rect 500052 102310 500234 102370
rect 500052 102308 500058 102310
rect 500174 102236 500234 102310
rect 487102 102234 487108 102236
rect 483013 102232 487108 102234
rect 483013 102176 483018 102232
rect 483074 102176 487108 102232
rect 483013 102174 487108 102176
rect 483013 102171 483079 102174
rect 487102 102172 487108 102174
rect 487172 102172 487178 102236
rect 492806 102172 492812 102236
rect 492876 102172 492882 102236
rect 495198 102234 495204 102236
rect 494102 102174 495204 102234
rect 24761 102098 24827 102101
rect 88333 102098 88399 102101
rect 24761 102096 88399 102098
rect 24761 102040 24766 102096
rect 24822 102040 88338 102096
rect 88394 102040 88399 102096
rect 24761 102038 88399 102040
rect 24761 102035 24827 102038
rect 88333 102035 88399 102038
rect 492857 102098 492923 102101
rect 492990 102098 492996 102100
rect 492857 102096 492996 102098
rect 492857 102040 492862 102096
rect 492918 102040 492996 102096
rect 492857 102038 492996 102040
rect 492857 102035 492923 102038
rect 492990 102036 492996 102038
rect 493060 102036 493066 102100
rect 494102 101965 494162 102174
rect 495198 102172 495204 102174
rect 495268 102172 495274 102236
rect 500166 102172 500172 102236
rect 500236 102172 500242 102236
rect 495249 102098 495315 102101
rect 580257 102098 580323 102101
rect 495249 102096 580323 102098
rect 495249 102040 495254 102096
rect 495310 102040 580262 102096
rect 580318 102040 580323 102096
rect 495249 102038 580323 102040
rect 495249 102035 495315 102038
rect 580257 102035 580323 102038
rect 76925 101962 76991 101965
rect 85573 101962 85639 101965
rect 76925 101960 85639 101962
rect 76925 101904 76930 101960
rect 76986 101904 85578 101960
rect 85634 101904 85639 101960
rect 76925 101902 85639 101904
rect 494102 101960 494211 101965
rect 494102 101904 494150 101960
rect 494206 101904 494211 101960
rect 494102 101902 494211 101904
rect 76925 101899 76991 101902
rect 85573 101899 85639 101902
rect 494145 101899 494211 101902
rect 324221 101826 324287 101829
rect 489126 101826 489132 101828
rect 324221 101824 489132 101826
rect 324221 101768 324226 101824
rect 324282 101768 489132 101824
rect 324221 101766 489132 101768
rect 324221 101763 324287 101766
rect 489126 101764 489132 101766
rect 489196 101764 489202 101828
rect 59169 101690 59235 101693
rect 89989 101690 90055 101693
rect 59169 101688 90055 101690
rect 59169 101632 59174 101688
rect 59230 101632 89994 101688
rect 90050 101632 90055 101688
rect 59169 101630 90055 101632
rect 59169 101627 59235 101630
rect 89989 101627 90055 101630
rect 241462 101628 241468 101692
rect 241532 101690 241538 101692
rect 251030 101690 251036 101692
rect 241532 101630 251036 101690
rect 241532 101628 241538 101630
rect 251030 101628 251036 101630
rect 251100 101628 251106 101692
rect 322841 101690 322907 101693
rect 517881 101690 517947 101693
rect 322841 101688 517947 101690
rect 322841 101632 322846 101688
rect 322902 101632 517886 101688
rect 517942 101632 517947 101688
rect 322841 101630 517947 101632
rect 322841 101627 322907 101630
rect 517881 101627 517947 101630
rect 73797 101554 73863 101557
rect 116117 101554 116183 101557
rect 73797 101552 116183 101554
rect 73797 101496 73802 101552
rect 73858 101496 116122 101552
rect 116178 101496 116183 101552
rect 73797 101494 116183 101496
rect 73797 101491 73863 101494
rect 116117 101491 116183 101494
rect 212257 101554 212323 101557
rect 516593 101554 516659 101557
rect 212257 101552 516659 101554
rect 212257 101496 212262 101552
rect 212318 101496 516598 101552
rect 516654 101496 516659 101552
rect 212257 101494 516659 101496
rect 212257 101491 212323 101494
rect 516593 101491 516659 101494
rect 72877 101418 72943 101421
rect 131205 101418 131271 101421
rect 72877 101416 131271 101418
rect 72877 101360 72882 101416
rect 72938 101360 131210 101416
rect 131266 101360 131271 101416
rect 72877 101358 131271 101360
rect 72877 101355 72943 101358
rect 131205 101355 131271 101358
rect 176561 101418 176627 101421
rect 493726 101418 493732 101420
rect 176561 101416 493732 101418
rect 176561 101360 176566 101416
rect 176622 101360 493732 101416
rect 176561 101358 493732 101360
rect 176561 101355 176627 101358
rect 493726 101356 493732 101358
rect 493796 101356 493802 101420
rect 395838 100948 395844 101012
rect 395908 101010 395914 101012
rect 402830 101010 402836 101012
rect 395908 100950 402836 101010
rect 395908 100948 395914 100950
rect 402830 100948 402836 100950
rect 402900 100948 402906 101012
rect 403750 100948 403756 101012
rect 403820 101010 403826 101012
rect 412398 101010 412404 101012
rect 403820 100950 412404 101010
rect 403820 100948 403826 100950
rect 412398 100948 412404 100950
rect 412468 100948 412474 101012
rect 481582 100948 481588 101012
rect 481652 101010 481658 101012
rect 495198 101010 495204 101012
rect 481652 100950 495204 101010
rect 481652 100948 481658 100950
rect 495198 100948 495204 100950
rect 495268 100948 495274 101012
rect 504582 100948 504588 101012
rect 504652 101010 504658 101012
rect 507158 101010 507164 101012
rect 504652 100950 507164 101010
rect 504652 100948 504658 100950
rect 507158 100948 507164 100950
rect 507228 100948 507234 101012
rect 193673 100874 193739 100877
rect 569217 100874 569283 100877
rect 193673 100872 569283 100874
rect 193673 100816 193678 100872
rect 193734 100816 569222 100872
rect 569278 100816 569283 100872
rect 193673 100814 569283 100816
rect 193673 100811 193739 100814
rect 569217 100811 569283 100814
rect 68870 100676 68876 100740
rect 68940 100738 68946 100740
rect 141785 100738 141851 100741
rect 68940 100736 141851 100738
rect 68940 100680 141790 100736
rect 141846 100680 141851 100736
rect 68940 100678 141851 100680
rect 68940 100676 68946 100678
rect 141785 100675 141851 100678
rect 171409 100738 171475 100741
rect 486366 100738 486372 100740
rect 171409 100736 486372 100738
rect 171409 100680 171414 100736
rect 171470 100680 486372 100736
rect 171409 100678 486372 100680
rect 171409 100675 171475 100678
rect 486366 100676 486372 100678
rect 486436 100676 486442 100740
rect 498878 100676 498884 100740
rect 498948 100738 498954 100740
rect 499113 100738 499179 100741
rect 498948 100736 499179 100738
rect 498948 100680 499118 100736
rect 499174 100680 499179 100736
rect 498948 100678 499179 100680
rect 498948 100676 498954 100678
rect 499113 100675 499179 100678
rect 77201 100602 77267 100605
rect 124489 100602 124555 100605
rect 77201 100600 124555 100602
rect 77201 100544 77206 100600
rect 77262 100544 124494 100600
rect 124550 100544 124555 100600
rect 77201 100542 124555 100544
rect 77201 100539 77267 100542
rect 124489 100539 124555 100542
rect 67449 100466 67515 100469
rect 87321 100466 87387 100469
rect 67449 100464 87387 100466
rect 67449 100408 67454 100464
rect 67510 100408 87326 100464
rect 87382 100408 87387 100464
rect 67449 100406 87387 100408
rect 67449 100403 67515 100406
rect 87321 100403 87387 100406
rect 231894 100268 231900 100332
rect 231964 100330 231970 100332
rect 241278 100330 241284 100332
rect 231964 100270 241284 100330
rect 231964 100268 231970 100270
rect 241278 100268 241284 100270
rect 241348 100268 241354 100332
rect 270534 100268 270540 100332
rect 270604 100330 270610 100332
rect 273846 100330 273852 100332
rect 270604 100270 273852 100330
rect 270604 100268 270610 100270
rect 273846 100268 273852 100270
rect 273916 100268 273922 100332
rect 347814 100268 347820 100332
rect 347884 100330 347890 100332
rect 351126 100330 351132 100332
rect 347884 100270 351132 100330
rect 347884 100268 347890 100270
rect 351126 100268 351132 100270
rect 351196 100268 351202 100332
rect 583520 99636 584960 99876
rect 406377 99106 406443 99109
rect 504214 99106 504220 99108
rect 406377 99104 504220 99106
rect 406377 99048 406382 99104
rect 406438 99048 504220 99104
rect 406377 99046 504220 99048
rect 406377 99043 406443 99046
rect 504214 99044 504220 99046
rect 504284 99044 504290 99108
rect 83222 98908 83228 98972
rect 83292 98970 83298 98972
rect 120073 98970 120139 98973
rect 83292 98968 120139 98970
rect 83292 98912 120078 98968
rect 120134 98912 120139 98968
rect 83292 98910 120139 98912
rect 83292 98908 83298 98910
rect 120073 98907 120139 98910
rect 289721 98970 289787 98973
rect 509325 98970 509391 98973
rect 289721 98968 509391 98970
rect 289721 98912 289726 98968
rect 289782 98912 509330 98968
rect 509386 98912 509391 98968
rect 289721 98910 509391 98912
rect 289721 98907 289787 98910
rect 509325 98907 509391 98910
rect 81566 98772 81572 98836
rect 81636 98834 81642 98836
rect 331213 98834 331279 98837
rect 81636 98832 331279 98834
rect 81636 98776 331218 98832
rect 331274 98776 331279 98832
rect 81636 98774 331279 98776
rect 81636 98772 81642 98774
rect 331213 98771 331279 98774
rect 344921 98834 344987 98837
rect 521878 98834 521884 98836
rect 344921 98832 521884 98834
rect 344921 98776 344926 98832
rect 344982 98776 521884 98832
rect 344921 98774 521884 98776
rect 344921 98771 344987 98774
rect 521878 98772 521884 98774
rect 521948 98772 521954 98836
rect 72366 98636 72372 98700
rect 72436 98698 72442 98700
rect 129733 98698 129799 98701
rect 72436 98696 129799 98698
rect 72436 98640 129738 98696
rect 129794 98640 129799 98696
rect 72436 98638 129799 98640
rect 72436 98636 72442 98638
rect 129733 98635 129799 98638
rect 237281 98698 237347 98701
rect 517973 98698 518039 98701
rect 237281 98696 518039 98698
rect 237281 98640 237286 98696
rect 237342 98640 517978 98696
rect 518034 98640 518039 98696
rect 237281 98638 518039 98640
rect 237281 98635 237347 98638
rect 517973 98635 518039 98638
rect 161473 97882 161539 97885
rect 519486 97882 519492 97884
rect 161473 97880 519492 97882
rect 161473 97824 161478 97880
rect 161534 97824 519492 97880
rect 161473 97822 519492 97824
rect 161473 97819 161539 97822
rect 519486 97820 519492 97822
rect 519556 97820 519562 97884
rect 304901 97338 304967 97341
rect 483013 97338 483079 97341
rect 304901 97336 483079 97338
rect 304901 97280 304906 97336
rect 304962 97280 483018 97336
rect 483074 97280 483079 97336
rect 304901 97278 483079 97280
rect 304901 97275 304967 97278
rect 483013 97275 483079 97278
rect 242801 97202 242867 97205
rect 499798 97202 499804 97204
rect 242801 97200 499804 97202
rect 242801 97144 242806 97200
rect 242862 97144 499804 97200
rect 242801 97142 499804 97144
rect 242801 97139 242867 97142
rect 499798 97140 499804 97142
rect 499868 97140 499874 97204
rect 198365 96658 198431 96661
rect 198733 96658 198799 96661
rect 198365 96656 198799 96658
rect 198365 96600 198370 96656
rect 198426 96600 198738 96656
rect 198794 96600 198799 96656
rect 198365 96598 198799 96600
rect 198365 96595 198431 96598
rect 198733 96595 198799 96598
rect 423397 96658 423463 96661
rect 423581 96658 423647 96661
rect 423397 96656 423647 96658
rect 423397 96600 423402 96656
rect 423458 96600 423586 96656
rect 423642 96600 423647 96656
rect 423397 96598 423647 96600
rect 423397 96595 423463 96598
rect 423581 96595 423647 96598
rect 445477 96658 445543 96661
rect 445661 96658 445727 96661
rect 445477 96656 445727 96658
rect 445477 96600 445482 96656
rect 445538 96600 445666 96656
rect 445722 96600 445727 96656
rect 445477 96598 445727 96600
rect 445477 96595 445543 96598
rect 445661 96595 445727 96598
rect 484485 96658 484551 96661
rect 487838 96658 487844 96660
rect 484485 96656 487844 96658
rect 484485 96600 484490 96656
rect 484546 96600 487844 96656
rect 484485 96598 487844 96600
rect 484485 96595 484551 96598
rect 487838 96596 487844 96598
rect 487908 96596 487914 96660
rect 488625 96658 488691 96661
rect 489862 96658 489868 96660
rect 488625 96656 489868 96658
rect 488625 96600 488630 96656
rect 488686 96600 489868 96656
rect 488625 96598 489868 96600
rect 488625 96595 488691 96598
rect 489862 96596 489868 96598
rect 489932 96596 489938 96660
rect 71078 96460 71084 96524
rect 71148 96522 71154 96524
rect 480161 96522 480227 96525
rect 71148 96520 480227 96522
rect 71148 96464 480166 96520
rect 480222 96464 480227 96520
rect 71148 96462 480227 96464
rect 71148 96460 71154 96462
rect 480161 96459 480227 96462
rect 357341 96114 357407 96117
rect 492857 96114 492923 96117
rect 357341 96112 492923 96114
rect 357341 96056 357346 96112
rect 357402 96056 492862 96112
rect 492918 96056 492923 96112
rect 357341 96054 492923 96056
rect 357341 96051 357407 96054
rect 492857 96051 492923 96054
rect 319989 95978 320055 95981
rect 492806 95978 492812 95980
rect 319989 95976 492812 95978
rect 319989 95920 319994 95976
rect 320050 95920 492812 95976
rect 319989 95918 492812 95920
rect 319989 95915 320055 95918
rect 492806 95916 492812 95918
rect 492876 95916 492882 95980
rect 164141 95842 164207 95845
rect 514937 95842 515003 95845
rect 164141 95840 515003 95842
rect 164141 95784 164146 95840
rect 164202 95784 514942 95840
rect 514998 95784 515003 95840
rect 164141 95782 515003 95784
rect 164141 95779 164207 95782
rect 514937 95779 515003 95782
rect 78254 94420 78260 94484
rect 78324 94482 78330 94484
rect 309133 94482 309199 94485
rect 78324 94480 309199 94482
rect 78324 94424 309138 94480
rect 309194 94424 309199 94480
rect 78324 94422 309199 94424
rect 78324 94420 78330 94422
rect 309133 94419 309199 94422
rect 496486 93876 496492 93940
rect 496556 93876 496562 93940
rect 496494 93668 496554 93876
rect 496486 93604 496492 93668
rect 496556 93604 496562 93668
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 81014 93060 81020 93124
rect 81084 93122 81090 93124
rect 563053 93122 563119 93125
rect 81084 93120 563119 93122
rect 81084 93064 563058 93120
rect 563114 93064 563119 93120
rect 81084 93062 563119 93064
rect 81084 93060 81090 93062
rect 563053 93059 563119 93062
rect 501270 92442 501276 92444
rect 501094 92382 501276 92442
rect 501094 92308 501154 92382
rect 501270 92380 501276 92382
rect 501340 92380 501346 92444
rect 501086 92244 501092 92308
rect 501156 92244 501162 92308
rect 79358 90476 79364 90540
rect 79428 90538 79434 90540
rect 454033 90538 454099 90541
rect 79428 90536 454099 90538
rect 79428 90480 454038 90536
rect 454094 90480 454099 90536
rect 79428 90478 454099 90480
rect 79428 90476 79434 90478
rect 454033 90475 454099 90478
rect 77201 90402 77267 90405
rect 509182 90402 509188 90404
rect 77201 90400 509188 90402
rect 77201 90344 77206 90400
rect 77262 90344 509188 90400
rect 77201 90342 509188 90344
rect 77201 90339 77267 90342
rect 509182 90340 509188 90342
rect 509252 90340 509258 90404
rect 67081 89724 67147 89725
rect 67030 89722 67036 89724
rect 66990 89662 67036 89722
rect 67100 89720 67147 89724
rect 67142 89664 67147 89720
rect 67030 89660 67036 89662
rect 67100 89660 67147 89664
rect 67081 89659 67147 89660
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 506422 87818 506428 87820
rect 500174 87758 506428 87818
rect 209681 87682 209747 87685
rect 500174 87682 500234 87758
rect 506422 87756 506428 87758
rect 506492 87756 506498 87820
rect 500493 87684 500559 87685
rect 500493 87682 500540 87684
rect 209681 87680 500234 87682
rect 209681 87624 209686 87680
rect 209742 87624 500234 87680
rect 209681 87622 500234 87624
rect 500448 87680 500540 87682
rect 500448 87624 500498 87680
rect 500448 87622 500540 87624
rect 209681 87619 209747 87622
rect 500493 87620 500540 87622
rect 500604 87620 500610 87684
rect 500493 87619 500559 87620
rect 79726 87484 79732 87548
rect 79796 87546 79802 87548
rect 511441 87546 511507 87549
rect 79796 87544 511507 87546
rect 79796 87488 511446 87544
rect 511502 87488 511507 87544
rect 79796 87486 511507 87488
rect 79796 87484 79802 87486
rect 511441 87483 511507 87486
rect 500166 87348 500172 87412
rect 500236 87410 500242 87412
rect 500718 87410 500724 87412
rect 500236 87350 500724 87410
rect 500236 87348 500242 87350
rect 500718 87348 500724 87350
rect 500788 87348 500794 87412
rect 514710 87214 534090 87274
rect 138013 87002 138079 87005
rect 140773 87002 140839 87005
rect 138013 87000 140839 87002
rect 138013 86944 138018 87000
rect 138074 86944 140778 87000
rect 140834 86944 140839 87000
rect 138013 86942 140839 86944
rect 138013 86939 138079 86942
rect 140773 86939 140839 86942
rect 511206 86940 511212 87004
rect 511276 87002 511282 87004
rect 514710 87002 514770 87214
rect 534030 87138 534090 87214
rect 557582 87214 567210 87274
rect 534030 87078 543658 87138
rect 511276 86942 514770 87002
rect 543598 87002 543658 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 543598 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 511276 86940 511282 86942
rect 83406 86260 83412 86324
rect 83476 86322 83482 86324
rect 213913 86322 213979 86325
rect 83476 86320 213979 86322
rect 83476 86264 213918 86320
rect 213974 86264 213979 86320
rect 83476 86262 213979 86264
rect 83476 86260 83482 86262
rect 213913 86259 213979 86262
rect 263409 86322 263475 86325
rect 505686 86322 505692 86324
rect 263409 86320 505692 86322
rect 263409 86264 263414 86320
rect 263470 86264 505692 86320
rect 263409 86262 505692 86264
rect 263409 86259 263475 86262
rect 505686 86260 505692 86262
rect 505756 86260 505762 86324
rect 81382 86124 81388 86188
rect 81452 86186 81458 86188
rect 448513 86186 448579 86189
rect 81452 86184 448579 86186
rect 81452 86128 448518 86184
rect 448574 86128 448579 86184
rect 81452 86126 448579 86128
rect 81452 86124 81458 86126
rect 448513 86123 448579 86126
rect 496486 85642 496492 85644
rect 496310 85582 496492 85642
rect 496310 85370 496370 85582
rect 496486 85580 496492 85582
rect 496556 85580 496562 85644
rect 496486 85370 496492 85372
rect 496310 85310 496492 85370
rect 496486 85308 496492 85310
rect 496556 85308 496562 85372
rect 422201 82106 422267 82109
rect 500493 82106 500559 82109
rect 422201 82104 500559 82106
rect 422201 82048 422206 82104
rect 422262 82048 500498 82104
rect 500554 82048 500559 82104
rect 422201 82046 500559 82048
rect 422201 82043 422267 82046
rect 500493 82043 500559 82046
rect 3417 80066 3483 80069
rect 510654 80066 510660 80068
rect 3417 80064 510660 80066
rect 3417 80008 3422 80064
rect 3478 80008 510660 80064
rect 3417 80006 510660 80008
rect 3417 80003 3483 80006
rect 510654 80004 510660 80006
rect 510724 80004 510730 80068
rect 135161 79386 135227 79389
rect 503846 79386 503852 79388
rect 135161 79384 503852 79386
rect 135161 79328 135166 79384
rect 135222 79328 503852 79384
rect 135161 79326 503852 79328
rect 135161 79323 135227 79326
rect 503846 79324 503852 79326
rect 503916 79324 503922 79388
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 74022 77828 74028 77892
rect 74092 77890 74098 77892
rect 481633 77890 481699 77893
rect 74092 77888 481699 77890
rect 74092 77832 481638 77888
rect 481694 77832 481699 77888
rect 74092 77830 481699 77832
rect 74092 77828 74098 77830
rect 481633 77827 481699 77830
rect 499614 77482 499620 77484
rect 499438 77422 499620 77482
rect 89897 77346 89963 77349
rect 90081 77346 90147 77349
rect 499438 77348 499498 77422
rect 499614 77420 499620 77422
rect 499684 77420 499690 77484
rect 89897 77344 90147 77346
rect 89897 77288 89902 77344
rect 89958 77288 90086 77344
rect 90142 77288 90147 77344
rect 89897 77286 90147 77288
rect 89897 77283 89963 77286
rect 90081 77283 90147 77286
rect 499430 77284 499436 77348
rect 499500 77284 499506 77348
rect 140497 77210 140563 77213
rect 140773 77210 140839 77213
rect 140497 77208 140839 77210
rect 140497 77152 140502 77208
rect 140558 77152 140778 77208
rect 140834 77152 140839 77208
rect 140497 77150 140839 77152
rect 140497 77147 140563 77150
rect 140773 77147 140839 77150
rect 280245 77210 280311 77213
rect 280429 77210 280495 77213
rect 280245 77208 280495 77210
rect 280245 77152 280250 77208
rect 280306 77152 280434 77208
rect 280490 77152 280495 77208
rect 280245 77150 280495 77152
rect 280245 77147 280311 77150
rect 280429 77147 280495 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 84101 75170 84167 75173
rect 499430 75170 499436 75172
rect 84101 75168 499436 75170
rect 84101 75112 84106 75168
rect 84162 75112 499436 75168
rect 84101 75110 499436 75112
rect 84101 75107 84167 75110
rect 499430 75108 499436 75110
rect 499500 75108 499506 75172
rect 67265 72452 67331 72453
rect 67214 72388 67220 72452
rect 67284 72450 67331 72452
rect 248321 72450 248387 72453
rect 505870 72450 505876 72452
rect 67284 72448 67376 72450
rect 67326 72392 67376 72448
rect 67284 72390 67376 72392
rect 248321 72448 505876 72450
rect 248321 72392 248326 72448
rect 248382 72392 505876 72448
rect 248321 72390 505876 72392
rect 67284 72388 67331 72390
rect 67265 72387 67331 72388
rect 248321 72387 248387 72390
rect 505870 72388 505876 72390
rect 505940 72388 505946 72452
rect 78438 71300 78444 71364
rect 78508 71362 78514 71364
rect 266353 71362 266419 71365
rect 78508 71360 266419 71362
rect 78508 71304 266358 71360
rect 266414 71304 266419 71360
rect 78508 71302 266419 71304
rect 78508 71300 78514 71302
rect 266353 71299 266419 71302
rect 266169 71226 266235 71229
rect 501638 71226 501644 71228
rect 266169 71224 501644 71226
rect 266169 71168 266174 71224
rect 266230 71168 501644 71224
rect 266169 71166 501644 71168
rect 266169 71163 266235 71166
rect 501638 71164 501644 71166
rect 501708 71164 501714 71228
rect 79542 71028 79548 71092
rect 79612 71090 79618 71092
rect 437565 71090 437631 71093
rect 79612 71088 437631 71090
rect 79612 71032 437570 71088
rect 437626 71032 437631 71088
rect 79612 71030 437631 71032
rect 79612 71028 79618 71030
rect 437565 71027 437631 71030
rect 76230 69532 76236 69596
rect 76300 69594 76306 69596
rect 509233 69594 509299 69597
rect 76300 69592 509299 69594
rect 76300 69536 509238 69592
rect 509294 69536 509299 69592
rect 76300 69534 509299 69536
rect 76300 69532 76306 69534
rect 509233 69531 509299 69534
rect 67265 67692 67331 67693
rect 67214 67690 67220 67692
rect 67174 67630 67220 67690
rect 67284 67688 67331 67692
rect 67326 67632 67331 67688
rect 67214 67628 67220 67630
rect 67284 67628 67331 67632
rect 67265 67627 67331 67628
rect 140497 67690 140563 67693
rect 140773 67690 140839 67693
rect 499113 67692 499179 67693
rect 499062 67690 499068 67692
rect 140497 67688 140839 67690
rect 140497 67632 140502 67688
rect 140558 67632 140778 67688
rect 140834 67632 140839 67688
rect 140497 67630 140839 67632
rect 499022 67630 499068 67690
rect 499132 67688 499179 67692
rect 499174 67632 499179 67688
rect 140497 67627 140563 67630
rect 140773 67627 140839 67630
rect 499062 67628 499068 67630
rect 499132 67628 499179 67632
rect 499113 67627 499179 67628
rect 499062 66948 499068 67012
rect 499132 67010 499138 67012
rect 499205 67010 499271 67013
rect 499132 67008 499271 67010
rect 499132 66952 499210 67008
rect 499266 66952 499271 67008
rect 499132 66950 499271 66952
rect 499132 66948 499138 66950
rect 499205 66947 499271 66950
rect 78070 66812 78076 66876
rect 78140 66874 78146 66876
rect 426433 66874 426499 66877
rect 78140 66872 426499 66874
rect 78140 66816 426438 66872
rect 426494 66816 426499 66872
rect 78140 66814 426499 66816
rect 78140 66812 78146 66814
rect 426433 66811 426499 66814
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 67214 60890 67220 60892
rect 67038 60830 67220 60890
rect 67038 60620 67098 60830
rect 67214 60828 67220 60830
rect 67284 60828 67290 60892
rect 500902 60828 500908 60892
rect 500972 60828 500978 60892
rect 67030 60556 67036 60620
rect 67100 60556 67106 60620
rect 500910 60618 500970 60828
rect 501086 60618 501092 60620
rect 500910 60558 501092 60618
rect 501086 60556 501092 60558
rect 501156 60556 501162 60620
rect 499205 60076 499271 60077
rect 499205 60074 499252 60076
rect 499160 60072 499252 60074
rect 499160 60016 499210 60072
rect 499160 60014 499252 60016
rect 499205 60012 499252 60014
rect 499316 60012 499322 60076
rect 499205 60011 499271 60012
rect 81750 59876 81756 59940
rect 81820 59938 81826 59940
rect 458173 59938 458239 59941
rect 81820 59936 458239 59938
rect 81820 59880 458178 59936
rect 458234 59880 458239 59936
rect 81820 59878 458239 59880
rect 81820 59876 81826 59878
rect 458173 59875 458239 59878
rect 67081 57900 67147 57901
rect 67030 57836 67036 57900
rect 67100 57898 67147 57900
rect 67100 57896 67192 57898
rect 67142 57840 67192 57896
rect 67100 57838 67192 57840
rect 67100 57836 67147 57838
rect 67081 57835 67147 57836
rect 340781 57218 340847 57221
rect 500350 57218 500356 57220
rect 340781 57216 500356 57218
rect 340781 57160 340786 57216
rect 340842 57160 500356 57216
rect 340781 57158 500356 57160
rect 340781 57155 340847 57158
rect 500350 57156 500356 57158
rect 500420 57156 500426 57220
rect 499205 55180 499271 55181
rect 499205 55178 499252 55180
rect 499160 55176 499252 55178
rect 499160 55120 499210 55176
rect 499160 55118 499252 55120
rect 499205 55116 499252 55118
rect 499316 55116 499322 55180
rect 499205 55115 499271 55116
rect 74206 53076 74212 53140
rect 74276 53138 74282 53140
rect 389173 53138 389239 53141
rect 74276 53136 389239 53138
rect 74276 53080 389178 53136
rect 389234 53080 389239 53136
rect 74276 53078 389239 53080
rect 74276 53076 74282 53078
rect 389173 53075 389239 53078
rect 583520 52716 584960 52956
rect 317321 51778 317387 51781
rect 502742 51778 502748 51780
rect 317321 51776 502748 51778
rect 317321 51720 317326 51776
rect 317382 51720 502748 51776
rect 317321 51718 502748 51720
rect 317321 51715 317387 51718
rect 502742 51716 502748 51718
rect 502812 51716 502818 51780
rect 67081 50964 67147 50965
rect 67030 50962 67036 50964
rect 66990 50902 67036 50962
rect 67100 50960 67147 50964
rect 67142 50904 67147 50960
rect 67030 50900 67036 50902
rect 67100 50900 67147 50904
rect 67081 50899 67147 50900
rect 400121 50418 400187 50421
rect 486182 50418 486188 50420
rect 400121 50416 486188 50418
rect 400121 50360 400126 50416
rect 400182 50360 486188 50416
rect 400121 50358 486188 50360
rect 400121 50355 400187 50358
rect 486182 50356 486188 50358
rect 486252 50356 486258 50420
rect 115749 50282 115815 50285
rect 502558 50282 502564 50284
rect 115749 50280 502564 50282
rect -960 50146 480 50236
rect 115749 50224 115754 50280
rect 115810 50224 502564 50280
rect 115749 50222 502564 50224
rect 115749 50219 115815 50222
rect 502558 50220 502564 50222
rect 502628 50220 502634 50284
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 81198 47500 81204 47564
rect 81268 47562 81274 47564
rect 433425 47562 433491 47565
rect 81268 47560 433491 47562
rect 81268 47504 433430 47560
rect 433486 47504 433491 47560
rect 81268 47502 433491 47504
rect 81268 47500 81274 47502
rect 433425 47499 433491 47502
rect 190361 46202 190427 46205
rect 506606 46202 506612 46204
rect 190361 46200 506612 46202
rect 190361 46144 190366 46200
rect 190422 46144 506612 46200
rect 190361 46142 506612 46144
rect 190361 46139 190427 46142
rect 506606 46140 506612 46142
rect 506676 46140 506682 46204
rect 499205 45796 499271 45797
rect 499205 45792 499252 45796
rect 499316 45794 499322 45796
rect 499205 45736 499210 45792
rect 499205 45732 499252 45736
rect 499316 45734 499362 45794
rect 499316 45732 499322 45734
rect 499205 45731 499271 45732
rect 496353 45522 496419 45525
rect 499205 45524 499271 45525
rect 496486 45522 496492 45524
rect 496353 45520 496492 45522
rect 496353 45464 496358 45520
rect 496414 45464 496492 45520
rect 496353 45462 496492 45464
rect 496353 45459 496419 45462
rect 496486 45460 496492 45462
rect 496556 45460 496562 45524
rect 499205 45522 499252 45524
rect 499160 45520 499252 45522
rect 499160 45464 499210 45520
rect 499160 45462 499252 45464
rect 499205 45460 499252 45462
rect 499316 45460 499322 45524
rect 500033 45522 500099 45525
rect 501086 45522 501092 45524
rect 500033 45520 501092 45522
rect 500033 45464 500038 45520
rect 500094 45464 501092 45520
rect 500033 45462 501092 45464
rect 499205 45459 499271 45460
rect 500033 45459 500099 45462
rect 501086 45460 501092 45462
rect 501156 45460 501162 45524
rect 140681 44842 140747 44845
rect 506790 44842 506796 44844
rect 140681 44840 506796 44842
rect 140681 44784 140686 44840
rect 140742 44784 506796 44840
rect 140681 44782 506796 44784
rect 140681 44779 140747 44782
rect 506790 44780 506796 44782
rect 506860 44780 506866 44844
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 496353 40764 496419 40765
rect 496302 40762 496308 40764
rect 496262 40702 496308 40762
rect 496372 40760 496419 40764
rect 496414 40704 496419 40760
rect 496302 40700 496308 40702
rect 496372 40700 496419 40704
rect 496353 40699 496419 40700
rect 499205 40764 499271 40765
rect 499205 40760 499252 40764
rect 499316 40762 499322 40764
rect 499205 40704 499210 40760
rect 499205 40700 499252 40704
rect 499316 40702 499362 40762
rect 499316 40700 499322 40702
rect 499205 40699 499271 40700
rect 64229 39266 64295 39269
rect 500033 39266 500099 39269
rect 64229 39264 500099 39266
rect 64229 39208 64234 39264
rect 64290 39208 500038 39264
rect 500094 39208 500099 39264
rect 64229 39206 500099 39208
rect 64229 39203 64295 39206
rect 500033 39203 500099 39206
rect 148961 36546 149027 36549
rect 505502 36546 505508 36548
rect 148961 36544 505508 36546
rect 148961 36488 148966 36544
rect 149022 36488 505508 36544
rect 148961 36486 505508 36488
rect 148961 36483 149027 36486
rect 505502 36484 505508 36486
rect 505572 36484 505578 36548
rect -960 35866 480 35956
rect 64086 35866 64092 35868
rect -960 35806 64092 35866
rect -960 35716 480 35806
rect 64086 35804 64092 35806
rect 64156 35804 64162 35868
rect 74390 35124 74396 35188
rect 74460 35186 74466 35188
rect 409873 35186 409939 35189
rect 74460 35184 409939 35186
rect 74460 35128 409878 35184
rect 409934 35128 409939 35184
rect 74460 35126 409939 35128
rect 74460 35124 74466 35126
rect 409873 35123 409939 35126
rect 13629 30970 13695 30973
rect 509366 30970 509372 30972
rect 13629 30968 509372 30970
rect 13629 30912 13634 30968
rect 13690 30912 509372 30968
rect 13629 30910 509372 30912
rect 13629 30907 13695 30910
rect 509366 30908 509372 30910
rect 509436 30908 509442 30972
rect 560201 29338 560267 29341
rect 583520 29338 584960 29428
rect 534030 29278 543842 29338
rect 409873 29202 409939 29205
rect 409873 29200 414076 29202
rect 409873 29144 409878 29200
rect 409934 29144 414076 29200
rect 409873 29142 414076 29144
rect 409873 29139 409939 29142
rect 414016 29069 414076 29142
rect 414013 29064 414079 29069
rect 414013 29008 414018 29064
rect 414074 29008 414079 29064
rect 414013 29003 414079 29008
rect 516726 29004 516732 29068
rect 516796 29066 516802 29068
rect 534030 29066 534090 29278
rect 543782 29202 543842 29278
rect 560201 29336 572730 29338
rect 560201 29280 560206 29336
rect 560262 29280 572730 29336
rect 560201 29278 572730 29280
rect 560201 29275 560267 29278
rect 553117 29202 553183 29205
rect 543782 29200 553183 29202
rect 543782 29144 553122 29200
rect 553178 29144 553183 29200
rect 543782 29142 553183 29144
rect 553117 29139 553183 29142
rect 516796 29006 534090 29066
rect 572670 29066 572730 29278
rect 583342 29278 584960 29338
rect 583342 29066 583402 29278
rect 583520 29188 584960 29278
rect 572670 29006 583402 29066
rect 516796 29004 516802 29006
rect 498326 28868 498332 28932
rect 498396 28868 498402 28932
rect 498334 28797 498394 28868
rect 498334 28792 498443 28797
rect 498334 28736 498382 28792
rect 498438 28736 498443 28792
rect 498334 28734 498443 28736
rect 498377 28731 498443 28734
rect 99189 26890 99255 26893
rect 504030 26890 504036 26892
rect 99189 26888 504036 26890
rect 99189 26832 99194 26888
rect 99250 26832 504036 26888
rect 99189 26830 504036 26832
rect 99189 26827 99255 26830
rect 504030 26828 504036 26830
rect 504100 26828 504106 26892
rect 33041 24170 33107 24173
rect 70894 24170 70900 24172
rect 33041 24168 70900 24170
rect 33041 24112 33046 24168
rect 33102 24112 70900 24168
rect 33041 24110 70900 24112
rect 33041 24107 33107 24110
rect 70894 24108 70900 24110
rect 70964 24108 70970 24172
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 498377 21178 498443 21181
rect 498510 21178 498516 21180
rect 498377 21176 498516 21178
rect 498377 21120 498382 21176
rect 498438 21120 498516 21176
rect 498377 21118 498516 21120
rect 498377 21115 498443 21118
rect 498510 21116 498516 21118
rect 498580 21116 498586 21180
rect 411161 19410 411227 19413
rect 411345 19410 411411 19413
rect 411161 19408 411411 19410
rect 411161 19352 411166 19408
rect 411222 19352 411350 19408
rect 411406 19352 411411 19408
rect 411161 19350 411411 19352
rect 411161 19347 411227 19350
rect 411345 19347 411411 19350
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 496302 12610 496308 12612
rect 496126 12550 496308 12610
rect 496126 12340 496186 12550
rect 496302 12548 496308 12550
rect 496372 12548 496378 12612
rect 496118 12276 496124 12340
rect 496188 12276 496194 12340
rect 75494 11732 75500 11796
rect 75564 11794 75570 11796
rect 386413 11794 386479 11797
rect 75564 11792 386479 11794
rect 75564 11736 386418 11792
rect 386474 11736 386479 11792
rect 75564 11734 386479 11736
rect 75564 11732 75570 11734
rect 386413 11731 386479 11734
rect 64597 11658 64663 11661
rect 495934 11658 495940 11660
rect 64597 11656 495940 11658
rect 64597 11600 64602 11656
rect 64658 11600 495940 11656
rect 64597 11598 495940 11600
rect 64597 11595 64663 11598
rect 495934 11596 495940 11598
rect 496004 11596 496010 11660
rect 66662 9284 66668 9348
rect 66732 9346 66738 9348
rect 253749 9346 253815 9349
rect 66732 9344 253815 9346
rect 66732 9288 253754 9344
rect 253810 9288 253815 9344
rect 66732 9286 253815 9288
rect 66732 9284 66738 9286
rect 253749 9283 253815 9286
rect 346669 9346 346735 9349
rect 491334 9346 491340 9348
rect 346669 9344 491340 9346
rect 346669 9288 346674 9344
rect 346730 9288 491340 9344
rect 346669 9286 491340 9288
rect 346669 9283 346735 9286
rect 491334 9284 491340 9286
rect 491404 9284 491410 9348
rect 73061 9210 73127 9213
rect 390645 9210 390711 9213
rect 73061 9208 390711 9210
rect 73061 9152 73066 9208
rect 73122 9152 390650 9208
rect 390706 9152 390711 9208
rect 73061 9150 390711 9152
rect 73061 9147 73127 9150
rect 390645 9147 390711 9150
rect 46841 9074 46907 9077
rect 369209 9074 369275 9077
rect 46841 9072 369275 9074
rect 46841 9016 46846 9072
rect 46902 9016 369214 9072
rect 369270 9016 369275 9072
rect 46841 9014 369275 9016
rect 46841 9011 46907 9014
rect 369209 9011 369275 9014
rect 395429 9074 395495 9077
rect 497406 9074 497412 9076
rect 395429 9072 497412 9074
rect 395429 9016 395434 9072
rect 395490 9016 497412 9072
rect 395429 9014 497412 9016
rect 395429 9011 395495 9014
rect 497406 9012 497412 9014
rect 497476 9012 497482 9076
rect 16021 8938 16087 8941
rect 498510 8938 498516 8940
rect 16021 8936 498516 8938
rect 16021 8880 16026 8936
rect 16082 8880 498516 8936
rect 16021 8878 498516 8880
rect 16021 8875 16087 8878
rect 498510 8876 498516 8878
rect 498580 8876 498586 8940
rect 295517 7578 295583 7581
rect 494830 7578 494836 7580
rect 295517 7576 494836 7578
rect 295517 7520 295522 7576
rect 295578 7520 494836 7576
rect 295517 7518 494836 7520
rect 295517 7515 295583 7518
rect 494830 7516 494836 7518
rect 494900 7516 494906 7580
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 471513 6762 471579 6765
rect 495566 6762 495572 6764
rect 471513 6760 495572 6762
rect 471513 6704 471518 6760
rect 471574 6704 495572 6760
rect 471513 6702 495572 6704
rect 471513 6699 471579 6702
rect 495566 6700 495572 6702
rect 495636 6700 495642 6764
rect 415393 6626 415459 6629
rect 424961 6626 425027 6629
rect 415393 6624 425027 6626
rect 415393 6568 415398 6624
rect 415454 6568 424966 6624
rect 425022 6568 425027 6624
rect 415393 6566 425027 6568
rect 415393 6563 415459 6566
rect 424961 6563 425027 6566
rect 425145 6626 425211 6629
rect 507894 6626 507900 6628
rect 425145 6624 507900 6626
rect 425145 6568 425150 6624
rect 425206 6568 507900 6624
rect 425145 6566 507900 6568
rect 425145 6563 425211 6566
rect 507894 6564 507900 6566
rect 507964 6564 507970 6628
rect 403709 6490 403775 6493
rect 492622 6490 492628 6492
rect 403709 6488 492628 6490
rect 403709 6432 403714 6488
rect 403770 6432 492628 6488
rect 403709 6430 492628 6432
rect 403709 6427 403775 6430
rect 492622 6428 492628 6430
rect 492692 6428 492698 6492
rect 72182 6292 72188 6356
rect 72252 6354 72258 6356
rect 325233 6354 325299 6357
rect 72252 6352 325299 6354
rect 72252 6296 325238 6352
rect 325294 6296 325299 6352
rect 72252 6294 325299 6296
rect 72252 6292 72258 6294
rect 325233 6291 325299 6294
rect 407297 6354 407363 6357
rect 496854 6354 496860 6356
rect 407297 6352 496860 6354
rect 407297 6296 407302 6352
rect 407358 6296 496860 6352
rect 407297 6294 496860 6296
rect 407297 6291 407363 6294
rect 496854 6292 496860 6294
rect 496924 6292 496930 6356
rect 69974 6156 69980 6220
rect 70044 6218 70050 6220
rect 536925 6218 536991 6221
rect 70044 6216 536991 6218
rect 70044 6160 536930 6216
rect 536986 6160 536991 6216
rect 70044 6158 536991 6160
rect 70044 6156 70050 6158
rect 536925 6155 536991 6158
rect 220629 6082 220695 6085
rect 222142 6082 222148 6084
rect 220629 6080 222148 6082
rect 220629 6024 220634 6080
rect 220690 6024 222148 6080
rect 220629 6022 222148 6024
rect 220629 6019 220695 6022
rect 222142 6020 222148 6022
rect 222212 6020 222218 6084
rect 230422 6020 230428 6084
rect 230492 6082 230498 6084
rect 239990 6082 239996 6084
rect 230492 6022 239996 6082
rect 230492 6020 230498 6022
rect 239990 6020 239996 6022
rect 240060 6020 240066 6084
rect 249742 6020 249748 6084
rect 249812 6082 249818 6084
rect 259361 6082 259427 6085
rect 249812 6080 259427 6082
rect 249812 6024 259366 6080
rect 259422 6024 259427 6080
rect 249812 6022 259427 6024
rect 249812 6020 249818 6022
rect 259361 6019 259427 6022
rect 288382 6020 288388 6084
rect 288452 6082 288458 6084
rect 297950 6082 297956 6084
rect 288452 6022 297956 6082
rect 288452 6020 288458 6022
rect 297950 6020 297956 6022
rect 298020 6020 298026 6084
rect 384982 6020 384988 6084
rect 385052 6082 385058 6084
rect 394601 6082 394667 6085
rect 385052 6080 394667 6082
rect 385052 6024 394606 6080
rect 394662 6024 394667 6080
rect 385052 6022 394667 6024
rect 385052 6020 385058 6022
rect 394601 6019 394667 6022
rect 405774 6020 405780 6084
rect 405844 6082 405850 6084
rect 415393 6082 415459 6085
rect 405844 6080 415459 6082
rect 405844 6024 415398 6080
rect 415454 6024 415459 6080
rect 405844 6022 415459 6024
rect 405844 6020 405850 6022
rect 415393 6019 415459 6022
rect 424961 6082 425027 6085
rect 424961 6080 433258 6082
rect 424961 6024 424966 6080
rect 425022 6024 433258 6080
rect 424961 6022 433258 6024
rect 424961 6019 425027 6022
rect 153142 5884 153148 5948
rect 153212 5946 153218 5948
rect 162761 5946 162827 5949
rect 201585 5946 201651 5949
rect 211061 5948 211127 5949
rect 211061 5946 211108 5948
rect 153212 5944 162827 5946
rect 153212 5888 162766 5944
rect 162822 5888 162827 5944
rect 153212 5886 162827 5888
rect 153212 5884 153218 5886
rect 162761 5883 162827 5886
rect 201542 5944 201651 5946
rect 201542 5888 201590 5944
rect 201646 5888 201651 5944
rect 201542 5883 201651 5888
rect 211020 5944 211108 5946
rect 211020 5888 211066 5944
rect 211020 5886 211108 5888
rect 211061 5884 211108 5886
rect 211172 5884 211178 5948
rect 433198 5946 433258 6022
rect 468477 5946 468543 5949
rect 481817 5946 481883 5949
rect 278638 5886 280170 5946
rect 433198 5886 433442 5946
rect 211061 5883 211127 5884
rect 77150 5748 77156 5812
rect 77220 5810 77226 5812
rect 135253 5810 135319 5813
rect 77220 5808 135319 5810
rect 77220 5752 135258 5808
rect 135314 5752 135319 5808
rect 77220 5750 135319 5752
rect 77220 5748 77226 5750
rect 135253 5747 135319 5750
rect 199929 5810 199995 5813
rect 201542 5810 201602 5883
rect 199929 5808 201602 5810
rect 199929 5752 199934 5808
rect 199990 5752 201602 5808
rect 199929 5750 201602 5752
rect 199929 5747 199995 5750
rect 239990 5748 239996 5812
rect 240060 5810 240066 5812
rect 249742 5810 249748 5812
rect 240060 5750 249748 5810
rect 240060 5748 240066 5750
rect 249742 5748 249748 5750
rect 249812 5748 249818 5812
rect 260966 5748 260972 5812
rect 261036 5810 261042 5812
rect 269062 5810 269068 5812
rect 261036 5750 269068 5810
rect 261036 5748 261042 5750
rect 269062 5748 269068 5750
rect 269132 5748 269138 5812
rect 273897 5810 273963 5813
rect 278638 5810 278698 5886
rect 273897 5808 278698 5810
rect 273897 5752 273902 5808
rect 273958 5752 278698 5808
rect 273897 5750 278698 5752
rect 280110 5810 280170 5886
rect 282821 5810 282887 5813
rect 280110 5808 282887 5810
rect 280110 5752 282826 5808
rect 282882 5752 282887 5808
rect 280110 5750 282887 5752
rect 273897 5747 273963 5750
rect 282821 5747 282887 5750
rect 283005 5810 283071 5813
rect 288382 5810 288388 5812
rect 283005 5808 288388 5810
rect 283005 5752 283010 5808
rect 283066 5752 288388 5808
rect 283005 5750 288388 5752
rect 283005 5747 283071 5750
rect 288382 5748 288388 5750
rect 288452 5748 288458 5812
rect 297950 5748 297956 5812
rect 298020 5810 298026 5812
rect 307702 5810 307708 5812
rect 298020 5750 307708 5810
rect 298020 5748 298026 5750
rect 307702 5748 307708 5750
rect 307772 5748 307778 5812
rect 317270 5748 317276 5812
rect 317340 5810 317346 5812
rect 330845 5810 330911 5813
rect 360142 5810 360148 5812
rect 317340 5808 330911 5810
rect 317340 5752 330850 5808
rect 330906 5752 330911 5808
rect 317340 5750 330911 5752
rect 317340 5748 317346 5750
rect 330845 5747 330911 5750
rect 341566 5750 346410 5810
rect 145005 5674 145071 5677
rect 153142 5674 153148 5676
rect 145005 5672 153148 5674
rect 145005 5616 145010 5672
rect 145066 5616 153148 5672
rect 145005 5614 153148 5616
rect 145005 5611 145071 5614
rect 153142 5612 153148 5614
rect 153212 5612 153218 5676
rect 182173 5674 182239 5677
rect 172470 5672 182239 5674
rect 172470 5616 182178 5672
rect 182234 5616 182239 5672
rect 172470 5614 182239 5616
rect 162761 5538 162827 5541
rect 163037 5538 163103 5541
rect 172470 5538 172530 5614
rect 182173 5611 182239 5614
rect 259361 5674 259427 5677
rect 260782 5674 260788 5676
rect 259361 5672 260788 5674
rect 259361 5616 259366 5672
rect 259422 5616 260788 5672
rect 259361 5614 260788 5616
rect 259361 5611 259427 5614
rect 260782 5612 260788 5614
rect 260852 5612 260858 5676
rect 330937 5674 331003 5677
rect 341566 5674 341626 5750
rect 330937 5672 341626 5674
rect 330937 5616 330942 5672
rect 330998 5616 341626 5672
rect 330937 5614 341626 5616
rect 346350 5674 346410 5750
rect 357390 5750 360148 5810
rect 350441 5674 350507 5677
rect 346350 5672 350507 5674
rect 346350 5616 350446 5672
rect 350502 5616 350507 5672
rect 346350 5614 350507 5616
rect 330937 5611 331003 5614
rect 350441 5611 350507 5614
rect 350625 5674 350691 5677
rect 357390 5674 357450 5750
rect 360142 5748 360148 5750
rect 360212 5748 360218 5812
rect 360326 5748 360332 5812
rect 360396 5810 360402 5812
rect 365662 5810 365668 5812
rect 360396 5750 365668 5810
rect 360396 5748 360402 5750
rect 365662 5748 365668 5750
rect 365732 5748 365738 5812
rect 375281 5810 375347 5813
rect 384982 5810 384988 5812
rect 375281 5808 384988 5810
rect 375281 5752 375286 5808
rect 375342 5752 384988 5808
rect 375281 5750 384988 5752
rect 375281 5747 375347 5750
rect 384982 5748 384988 5750
rect 385052 5748 385058 5812
rect 433382 5810 433442 5886
rect 468477 5944 481883 5946
rect 468477 5888 468482 5944
rect 468538 5888 481822 5944
rect 481878 5888 481883 5944
rect 468477 5886 481883 5888
rect 468477 5883 468543 5886
rect 481817 5883 481883 5886
rect 491201 5946 491267 5949
rect 491201 5944 502442 5946
rect 491201 5888 491206 5944
rect 491262 5888 502442 5944
rect 491201 5886 502442 5888
rect 491201 5883 491267 5886
rect 438117 5810 438183 5813
rect 433382 5808 438183 5810
rect 433382 5752 438122 5808
rect 438178 5752 438183 5808
rect 433382 5750 438183 5752
rect 438117 5747 438183 5750
rect 442901 5810 442967 5813
rect 447041 5810 447107 5813
rect 456742 5810 456748 5812
rect 442901 5808 447107 5810
rect 442901 5752 442906 5808
rect 442962 5752 447046 5808
rect 447102 5752 447107 5808
rect 442901 5750 447107 5752
rect 442901 5747 442967 5750
rect 447041 5747 447107 5750
rect 453990 5750 456748 5810
rect 350625 5672 357450 5674
rect 350625 5616 350630 5672
rect 350686 5616 357450 5672
rect 350625 5614 357450 5616
rect 394601 5674 394667 5677
rect 405774 5674 405780 5676
rect 394601 5672 405780 5674
rect 394601 5616 394606 5672
rect 394662 5616 405780 5672
rect 394601 5614 405780 5616
rect 350625 5611 350691 5614
rect 394601 5611 394667 5614
rect 405774 5612 405780 5614
rect 405844 5612 405850 5676
rect 447225 5674 447291 5677
rect 453990 5674 454050 5750
rect 456742 5748 456748 5750
rect 456812 5748 456818 5812
rect 456926 5748 456932 5812
rect 456996 5810 457002 5812
rect 502382 5810 502442 5886
rect 514661 5810 514727 5813
rect 456996 5750 463802 5810
rect 502382 5808 514727 5810
rect 502382 5752 514666 5808
rect 514722 5752 514727 5808
rect 502382 5750 514727 5752
rect 456996 5748 457002 5750
rect 447225 5672 454050 5674
rect 447225 5616 447230 5672
rect 447286 5616 454050 5672
rect 447225 5614 454050 5616
rect 447225 5611 447291 5614
rect 162761 5536 162962 5538
rect 162761 5480 162766 5536
rect 162822 5480 162962 5536
rect 162761 5478 162962 5480
rect 162761 5475 162827 5478
rect 162902 5405 162962 5478
rect 163037 5536 172530 5538
rect 163037 5480 163042 5536
rect 163098 5480 172530 5536
rect 163037 5478 172530 5480
rect 163037 5475 163103 5478
rect 222142 5476 222148 5540
rect 222212 5538 222218 5540
rect 230422 5538 230428 5540
rect 222212 5478 230428 5538
rect 222212 5476 222218 5478
rect 230422 5476 230428 5478
rect 230492 5476 230498 5540
rect 269062 5476 269068 5540
rect 269132 5538 269138 5540
rect 273897 5538 273963 5541
rect 269132 5536 273963 5538
rect 269132 5480 273902 5536
rect 273958 5480 273963 5536
rect 269132 5478 273963 5480
rect 269132 5476 269138 5478
rect 273897 5475 273963 5478
rect 307702 5476 307708 5540
rect 307772 5538 307778 5540
rect 317270 5538 317276 5540
rect 307772 5478 317276 5538
rect 307772 5476 307778 5478
rect 317270 5476 317276 5478
rect 317340 5476 317346 5540
rect 365662 5476 365668 5540
rect 365732 5538 365738 5540
rect 375281 5538 375347 5541
rect 365732 5536 375347 5538
rect 365732 5480 375286 5536
rect 375342 5480 375347 5536
rect 365732 5478 375347 5480
rect 463742 5538 463802 5750
rect 514661 5747 514727 5750
rect 514845 5810 514911 5813
rect 526437 5810 526503 5813
rect 535494 5810 535500 5812
rect 514845 5808 521762 5810
rect 514845 5752 514850 5808
rect 514906 5752 521762 5808
rect 514845 5750 521762 5752
rect 514845 5747 514911 5750
rect 468477 5538 468543 5541
rect 463742 5536 468543 5538
rect 463742 5480 468482 5536
rect 468538 5480 468543 5536
rect 463742 5478 468543 5480
rect 521702 5538 521762 5750
rect 526437 5808 535500 5810
rect 526437 5752 526442 5808
rect 526498 5752 535500 5808
rect 526437 5750 535500 5752
rect 526437 5747 526503 5750
rect 535494 5748 535500 5750
rect 535564 5748 535570 5812
rect 583520 5796 584960 6036
rect 526437 5538 526503 5541
rect 521702 5536 526503 5538
rect 521702 5480 526442 5536
rect 526498 5480 526503 5536
rect 521702 5478 526503 5480
rect 365732 5476 365738 5478
rect 375281 5475 375347 5478
rect 468477 5475 468543 5478
rect 526437 5475 526503 5478
rect 162902 5400 163011 5405
rect 162902 5344 162950 5400
rect 163006 5344 163011 5400
rect 162902 5342 163011 5344
rect 162945 5339 163011 5342
rect 211102 5340 211108 5404
rect 211172 5402 211178 5404
rect 220629 5402 220695 5405
rect 211172 5400 220695 5402
rect 211172 5344 220634 5400
rect 220690 5344 220695 5400
rect 211172 5342 220695 5344
rect 211172 5340 211178 5342
rect 220629 5339 220695 5342
rect 55213 4858 55279 4861
rect 499246 4858 499252 4860
rect 55213 4856 499252 4858
rect 55213 4800 55218 4856
rect 55274 4800 499252 4856
rect 55213 4798 499252 4800
rect 55213 4795 55279 4798
rect 499246 4796 499252 4798
rect 499316 4796 499322 4860
rect 169385 4042 169451 4045
rect 169518 4042 169524 4044
rect 169385 4040 169524 4042
rect 169385 3984 169390 4040
rect 169446 3984 169524 4040
rect 169385 3982 169524 3984
rect 169385 3979 169451 3982
rect 169518 3980 169524 3982
rect 169588 3980 169594 4044
rect 488574 3980 488580 4044
rect 488644 4042 488650 4044
rect 489361 4042 489427 4045
rect 488644 4040 489427 4042
rect 488644 3984 489366 4040
rect 489422 3984 489427 4040
rect 488644 3982 489427 3984
rect 488644 3980 488650 3982
rect 489361 3979 489427 3982
rect 535494 3980 535500 4044
rect 535564 4042 535570 4044
rect 535729 4042 535795 4045
rect 535564 4040 535795 4042
rect 535564 3984 535734 4040
rect 535790 3984 535795 4040
rect 535564 3982 535795 3984
rect 535564 3980 535570 3982
rect 535729 3979 535795 3982
rect 69657 3906 69723 3909
rect 73245 3906 73311 3909
rect 69657 3904 73311 3906
rect 69657 3848 69662 3904
rect 69718 3848 73250 3904
rect 73306 3848 73311 3904
rect 69657 3846 73311 3848
rect 69657 3843 69723 3846
rect 73245 3843 73311 3846
rect 464429 3906 464495 3909
rect 490230 3906 490236 3908
rect 464429 3904 490236 3906
rect 464429 3848 464434 3904
rect 464490 3848 490236 3904
rect 464429 3846 490236 3848
rect 464429 3843 464495 3846
rect 490230 3844 490236 3846
rect 490300 3844 490306 3908
rect 23105 3770 23171 3773
rect 75126 3770 75132 3772
rect 23105 3768 75132 3770
rect 23105 3712 23110 3768
rect 23166 3712 75132 3768
rect 23105 3710 75132 3712
rect 23105 3707 23171 3710
rect 75126 3708 75132 3710
rect 75196 3708 75202 3772
rect 75453 3770 75519 3773
rect 75678 3770 75684 3772
rect 75453 3768 75684 3770
rect 75453 3712 75458 3768
rect 75514 3712 75684 3768
rect 75453 3710 75684 3712
rect 75453 3707 75519 3710
rect 75678 3708 75684 3710
rect 75748 3708 75754 3772
rect 451365 3770 451431 3773
rect 485998 3770 486004 3772
rect 451365 3768 486004 3770
rect 451365 3712 451370 3768
rect 451426 3712 486004 3768
rect 451365 3710 486004 3712
rect 451365 3707 451431 3710
rect 485998 3708 486004 3710
rect 486068 3708 486074 3772
rect 490557 3770 490623 3773
rect 516133 3770 516199 3773
rect 490557 3768 516199 3770
rect 490557 3712 490562 3768
rect 490618 3712 516138 3768
rect 516194 3712 516199 3768
rect 490557 3710 516199 3712
rect 490557 3707 490623 3710
rect 516133 3707 516199 3710
rect 71681 3634 71747 3637
rect 263317 3634 263383 3637
rect 71681 3632 263383 3634
rect 71681 3576 71686 3632
rect 71742 3576 263322 3632
rect 263378 3576 263383 3632
rect 71681 3574 263383 3576
rect 71681 3571 71747 3574
rect 263317 3571 263383 3574
rect 450169 3634 450235 3637
rect 491886 3634 491892 3636
rect 450169 3632 491892 3634
rect 450169 3576 450174 3632
rect 450230 3576 491892 3632
rect 450169 3574 491892 3576
rect 450169 3571 450235 3574
rect 491886 3572 491892 3574
rect 491956 3572 491962 3636
rect 67173 3498 67239 3501
rect 67398 3498 67404 3500
rect 67173 3496 67404 3498
rect 67173 3440 67178 3496
rect 67234 3440 67404 3496
rect 67173 3438 67404 3440
rect 67173 3435 67239 3438
rect 67398 3436 67404 3438
rect 67468 3436 67474 3500
rect 72550 3436 72556 3500
rect 72620 3498 72626 3500
rect 73061 3498 73127 3501
rect 72620 3496 73127 3498
rect 72620 3440 73066 3496
rect 73122 3440 73127 3496
rect 72620 3438 73127 3440
rect 72620 3436 72626 3438
rect 73061 3435 73127 3438
rect 73245 3498 73311 3501
rect 299105 3498 299171 3501
rect 73245 3496 299171 3498
rect 73245 3440 73250 3496
rect 73306 3440 299110 3496
rect 299166 3440 299171 3496
rect 73245 3438 299171 3440
rect 73245 3435 73311 3438
rect 299105 3435 299171 3438
rect 381169 3498 381235 3501
rect 501454 3498 501460 3500
rect 381169 3496 501460 3498
rect 381169 3440 381174 3496
rect 381230 3440 501460 3496
rect 381169 3438 501460 3440
rect 381169 3435 381235 3438
rect 501454 3436 501460 3438
rect 501524 3436 501530 3500
rect 71313 3362 71379 3365
rect 504817 3362 504883 3365
rect 71313 3360 504883 3362
rect 71313 3304 71318 3360
rect 71374 3304 504822 3360
rect 504878 3304 504883 3360
rect 71313 3302 504883 3304
rect 71313 3299 71379 3302
rect 504817 3299 504883 3302
rect 5257 2818 5323 2821
rect 133689 2818 133755 2821
rect 5257 2816 133755 2818
rect 5257 2760 5262 2816
rect 5318 2760 133694 2816
rect 133750 2760 133755 2816
rect 5257 2758 133755 2760
rect 5257 2755 5323 2758
rect 133689 2755 133755 2758
rect 465625 2818 465691 2821
rect 466126 2818 466132 2820
rect 465625 2816 466132 2818
rect 465625 2760 465630 2816
rect 465686 2760 466132 2816
rect 465625 2758 466132 2760
rect 465625 2755 465691 2758
rect 466126 2756 466132 2758
rect 466196 2756 466202 2820
<< via3 >>
rect 68876 700300 68940 700364
rect 486372 700300 486436 700364
rect 519492 697172 519556 697236
rect 512684 681804 512748 681868
rect 183508 674052 183572 674116
rect 70164 673508 70228 673572
rect 183508 673780 183572 673844
rect 489868 607548 489932 607612
rect 487844 607412 487908 607476
rect 491156 607276 491220 607340
rect 428228 606596 428292 606660
rect 437796 606596 437860 606660
rect 458772 606596 458836 606660
rect 500908 606460 500972 606524
rect 235948 606188 236012 606252
rect 244412 606188 244476 606252
rect 253980 606188 254044 606252
rect 272932 606188 272996 606252
rect 273300 606188 273364 606252
rect 502380 606324 502444 606388
rect 507900 606188 507964 606252
rect 118924 606052 118988 606116
rect 128676 606052 128740 606116
rect 138428 606052 138492 606116
rect 157196 606052 157260 606116
rect 176884 606052 176948 606116
rect 195836 606052 195900 606116
rect 196572 606052 196636 606116
rect 207060 606052 207124 606116
rect 499436 606052 499500 606116
rect 516732 605916 516796 605980
rect 89116 605508 89180 605572
rect 90220 605508 90284 605572
rect 109724 605508 109788 605572
rect 118556 605508 118620 605572
rect 157748 605508 157812 605572
rect 176516 605508 176580 605572
rect 492812 604964 492876 605028
rect 67404 604828 67468 604892
rect 491892 604828 491956 604892
rect 496860 604692 496924 604756
rect 108436 604148 108500 604212
rect 109724 604148 109788 604212
rect 147444 604148 147508 604212
rect 157932 604148 157996 604212
rect 223620 604148 223684 604212
rect 224908 604148 224972 604212
rect 263364 604148 263428 604212
rect 264468 604148 264532 604212
rect 281212 604148 281276 604212
rect 283052 604148 283116 604212
rect 378548 604148 378612 604212
rect 389036 604148 389100 604212
rect 414428 604148 414492 604212
rect 421604 604148 421668 604212
rect 437244 604148 437308 604212
rect 453988 604148 454052 604212
rect 86908 604012 86972 604076
rect 86908 603740 86972 603804
rect 153148 604012 153212 604076
rect 153148 603740 153212 603804
rect 488580 604012 488644 604076
rect 384988 603876 385052 603940
rect 70900 603604 70964 603668
rect 384988 603604 385052 603668
rect 453988 603740 454052 603804
rect 89668 603468 89732 603532
rect 72372 603332 72436 603396
rect 486004 603332 486068 603396
rect 82860 603196 82924 603260
rect 495940 603060 496004 603124
rect 496860 602924 496924 602988
rect 497228 602788 497292 602852
rect 482876 602380 482940 602444
rect 492628 602244 492692 602308
rect 72556 602108 72620 602172
rect 488580 602108 488644 602172
rect 75132 601972 75196 602036
rect 501644 601700 501708 601764
rect 75868 601292 75932 601356
rect 162900 601352 162964 601356
rect 162900 601296 162914 601352
rect 162914 601296 162964 601352
rect 162900 601292 162964 601296
rect 200620 601292 200684 601356
rect 200804 601292 200868 601356
rect 258764 601292 258828 601356
rect 260788 601292 260852 601356
rect 270356 601292 270420 601356
rect 270540 601292 270604 601356
rect 86908 601156 86972 601220
rect 75868 601020 75932 601084
rect 135116 601156 135180 601220
rect 86908 600884 86972 600948
rect 124260 601020 124324 601084
rect 153148 601156 153212 601220
rect 167684 601156 167748 601220
rect 172284 601156 172348 601220
rect 124076 600884 124140 600948
rect 135116 600884 135180 600948
rect 153148 600884 153212 600948
rect 172284 600884 172348 600948
rect 195836 600884 195900 600948
rect 202828 600884 202892 600948
rect 215340 601020 215404 601084
rect 215156 600884 215220 600948
rect 234660 601020 234724 601084
rect 234476 600884 234540 600948
rect 253980 601020 254044 601084
rect 260788 601020 260852 601084
rect 270356 601020 270420 601084
rect 253796 600884 253860 600948
rect 270540 600884 270604 600948
rect 167684 600748 167748 600812
rect 301452 601292 301516 601356
rect 405044 601292 405108 601356
rect 409092 601292 409156 601356
rect 476988 601352 477052 601356
rect 476988 601296 477002 601352
rect 477002 601296 477052 601352
rect 476988 601292 477052 601296
rect 486188 601292 486252 601356
rect 494836 601292 494900 601356
rect 497596 600884 497660 600948
rect 498332 600748 498396 600812
rect 167684 600612 167748 600676
rect 172284 600612 172348 600676
rect 200804 600612 200868 600676
rect 258764 600612 258828 600676
rect 495388 600612 495452 600676
rect 301452 600476 301516 600540
rect 409092 600476 409156 600540
rect 494284 600476 494348 600540
rect 200620 600340 200684 600404
rect 511212 600340 511276 600404
rect 75684 600068 75748 600132
rect 82860 600204 82924 600268
rect 167684 600204 167748 600268
rect 172284 600204 172348 600268
rect 195836 600204 195900 600268
rect 202644 600204 202708 600268
rect 499804 600204 499868 600268
rect 80836 600068 80900 600132
rect 89668 600068 89732 600132
rect 487844 600068 487908 600132
rect 488212 600068 488276 600132
rect 162900 599932 162964 599996
rect 405044 599932 405108 599996
rect 482876 599932 482940 599996
rect 489868 599932 489932 599996
rect 491156 599932 491220 599996
rect 493180 599932 493244 599996
rect 405044 599388 405108 599452
rect 511580 598028 511644 598092
rect 515260 598028 515324 598092
rect 513420 596260 513484 596324
rect 82492 595444 82556 595508
rect 522068 592044 522132 592108
rect 521884 591772 521948 591836
rect 501644 589324 501708 589388
rect 501828 589052 501892 589116
rect 78444 588372 78508 588436
rect 66852 582388 66916 582452
rect 521884 582388 521948 582452
rect 67036 582116 67100 582180
rect 522068 582116 522132 582180
rect 81388 581300 81452 581364
rect 501644 579668 501708 579732
rect 501644 579532 501708 579596
rect 522068 579532 522132 579596
rect 505508 579124 505572 579188
rect 67036 578232 67100 578236
rect 67036 578176 67050 578232
rect 67050 578176 67100 578232
rect 67036 578172 67100 578176
rect 67036 572656 67100 572660
rect 67036 572600 67050 572656
rect 67050 572600 67100 572656
rect 67036 572596 67100 572600
rect 521884 570012 521948 570076
rect 521884 563076 521948 563140
rect 522068 562804 522132 562868
rect 522068 560280 522132 560284
rect 522068 560224 522118 560280
rect 522118 560224 522132 560280
rect 522068 560220 522132 560224
rect 506428 557092 506492 557156
rect 501644 554916 501708 554980
rect 501828 554780 501892 554844
rect 66852 553420 66916 553484
rect 67036 553148 67100 553212
rect 77156 551924 77220 551988
rect 522252 550700 522316 550764
rect 78260 548388 78324 548452
rect 67036 543900 67100 543964
rect 74212 543764 74276 543828
rect 522252 543900 522316 543964
rect 522068 543628 522132 543692
rect 67036 543492 67100 543556
rect 74396 541044 74460 541108
rect 522068 540968 522132 540972
rect 522068 540912 522082 540968
rect 522082 540912 522132 540968
rect 522068 540908 522132 540912
rect 76236 537236 76300 537300
rect 67036 534304 67100 534308
rect 67036 534248 67050 534304
rect 67050 534248 67100 534304
rect 67036 534244 67100 534248
rect 81204 533700 81268 533764
rect 504220 531524 504284 531588
rect 67036 531388 67100 531452
rect 521884 531388 521948 531452
rect 501276 526356 501340 526420
rect 67036 524724 67100 524788
rect 502012 524724 502076 524788
rect 521884 524452 521948 524516
rect 66668 524180 66732 524244
rect 522068 524180 522132 524244
rect 79732 522820 79796 522884
rect 501276 522820 501340 522884
rect 501828 522336 501892 522340
rect 501828 522280 501878 522336
rect 501878 522280 501892 522336
rect 501828 522276 501892 522280
rect 66668 521596 66732 521660
rect 522068 521656 522132 521660
rect 522068 521600 522082 521656
rect 522082 521600 522132 521656
rect 522068 521596 522132 521600
rect 502564 517108 502628 517172
rect 81572 515476 81636 515540
rect 505692 513300 505756 513364
rect 66484 512076 66548 512140
rect 521884 512076 521948 512140
rect 66484 510444 66548 510508
rect 502748 509764 502812 509828
rect 502012 507784 502076 507788
rect 502012 507728 502062 507784
rect 502062 507728 502076 507784
rect 502012 507724 502076 507728
rect 501460 505548 501524 505612
rect 521884 505140 521948 505204
rect 521700 504868 521764 504932
rect 510660 502420 510724 502484
rect 521700 502284 521764 502348
rect 67036 500924 67100 500988
rect 502012 498204 502076 498268
rect 521884 492628 521948 492692
rect 67036 491192 67100 491196
rect 67036 491136 67050 491192
rect 67050 491136 67100 491192
rect 67036 491132 67100 491136
rect 501460 490996 501524 491060
rect 79548 489908 79612 489972
rect 501644 487460 501708 487524
rect 502012 487460 502076 487524
rect 33732 487188 33796 487252
rect 46796 487188 46860 487252
rect 17908 485828 17972 485892
rect 27476 485828 27540 485892
rect 521884 485828 521948 485892
rect 521700 485556 521764 485620
rect 67036 483712 67100 483716
rect 67036 483656 67050 483712
rect 67050 483656 67100 483712
rect 67036 483652 67100 483656
rect 502012 481536 502076 481540
rect 502012 481480 502026 481536
rect 502026 481480 502076 481536
rect 502012 481476 502076 481480
rect 505876 480388 505940 480452
rect 67036 478816 67100 478820
rect 67036 478760 67050 478816
rect 67050 478760 67100 478816
rect 67036 478756 67100 478760
rect 521700 476036 521764 476100
rect 522436 476036 522500 476100
rect 82492 474948 82556 475012
rect 502012 472016 502076 472020
rect 502012 471960 502026 472016
rect 502026 471960 502076 472016
rect 502012 471956 502076 471960
rect 502012 471880 502076 471884
rect 502012 471824 502062 471880
rect 502062 471824 502076 471880
rect 502012 471820 502076 471824
rect 67036 469432 67100 469436
rect 67036 469376 67050 469432
rect 67050 469376 67100 469432
rect 67036 469372 67100 469376
rect 67036 469100 67100 469164
rect 82492 467604 82556 467668
rect 522436 466516 522500 466580
rect 522252 466244 522316 466308
rect 506612 465972 506676 466036
rect 522252 463524 522316 463588
rect 502012 462632 502076 462636
rect 502012 462576 502062 462632
rect 502062 462576 502076 462632
rect 502012 462572 502076 462576
rect 66852 459580 66916 459644
rect 501644 458900 501708 458964
rect 501644 458220 501708 458284
rect 506796 454820 506860 454884
rect 521884 454004 521948 454068
rect 502012 452704 502076 452708
rect 502012 452648 502026 452704
rect 502026 452648 502076 452704
rect 502012 452644 502076 452648
rect 10180 452508 10244 452572
rect 521884 447204 521948 447268
rect 522068 446932 522132 446996
rect 67036 446388 67100 446452
rect 502012 442912 502076 442916
rect 502012 442856 502062 442912
rect 502062 442856 502076 442912
rect 502012 442852 502076 442856
rect 521700 437412 521764 437476
rect 522252 437412 522316 437476
rect 66668 434752 66732 434756
rect 66668 434696 66718 434752
rect 66718 434696 66732 434752
rect 66668 434692 66732 434696
rect 67404 434556 67468 434620
rect 502012 433392 502076 433396
rect 502012 433336 502062 433392
rect 502062 433336 502076 433392
rect 502012 433332 502076 433336
rect 67404 429796 67468 429860
rect 502012 428496 502076 428500
rect 502012 428440 502062 428496
rect 502062 428440 502076 428496
rect 502012 428436 502076 428440
rect 522252 427892 522316 427956
rect 522068 427620 522132 427684
rect 522068 424900 522132 424964
rect 74028 423676 74092 423740
rect 509372 418372 509436 418436
rect 502012 415440 502076 415444
rect 502012 415384 502026 415440
rect 502026 415384 502076 415440
rect 502012 415380 502076 415384
rect 521884 415380 521948 415444
rect 502012 413944 502076 413948
rect 502012 413888 502062 413944
rect 502062 413888 502076 413944
rect 502012 413884 502076 413888
rect 521884 408580 521948 408644
rect 521700 408308 521764 408372
rect 521700 405588 521764 405652
rect 502012 404364 502076 404428
rect 67220 398924 67284 398988
rect 66852 396128 66916 396132
rect 66852 396072 66902 396128
rect 66902 396072 66916 396128
rect 66852 396068 66916 396072
rect 521884 396068 521948 396132
rect 66852 394572 66916 394636
rect 502012 394632 502076 394636
rect 502012 394576 502062 394632
rect 502062 394576 502076 394632
rect 502012 394572 502076 394576
rect 67036 394436 67100 394500
rect 521884 389268 521948 389332
rect 522068 388996 522132 389060
rect 522068 386276 522132 386340
rect 502012 385052 502076 385116
rect 67036 383556 67100 383620
rect 82492 377028 82556 377092
rect 522252 376816 522316 376820
rect 522252 376760 522266 376816
rect 522266 376760 522316 376816
rect 522252 376756 522316 376760
rect 67220 374036 67284 374100
rect 66852 373764 66916 373828
rect 67220 373764 67284 373828
rect 81756 372948 81820 373012
rect 522252 369956 522316 370020
rect 522068 369684 522132 369748
rect 71084 365740 71148 365804
rect 78076 365604 78140 365668
rect 501828 360844 501892 360908
rect 521884 357308 521948 357372
rect 502196 356084 502260 356148
rect 502196 354648 502260 354652
rect 502196 354592 502246 354648
rect 502246 354592 502260 354648
rect 502196 354588 502260 354592
rect 67220 350644 67284 350708
rect 66852 350508 66916 350572
rect 521700 350508 521764 350572
rect 501644 348468 501708 348532
rect 521700 347652 521764 347716
rect 502196 345068 502260 345132
rect 66852 340988 66916 341052
rect 67036 340716 67100 340780
rect 502196 339628 502260 339692
rect 502012 339356 502076 339420
rect 521884 338132 521948 338196
rect 67036 336636 67100 336700
rect 502012 335336 502076 335340
rect 502012 335280 502062 335336
rect 502062 335280 502076 335336
rect 502012 335276 502076 335280
rect 521884 331332 521948 331396
rect 522068 331060 522132 331124
rect 67404 328340 67468 328404
rect 522068 328340 522132 328404
rect 66668 327116 66732 327180
rect 502196 325756 502260 325820
rect 67404 323580 67468 323644
rect 501460 321676 501524 321740
rect 521884 318820 521948 318884
rect 67036 312020 67100 312084
rect 521884 312020 521948 312084
rect 501460 311884 501524 311948
rect 66852 311748 66916 311812
rect 522068 311748 522132 311812
rect 522068 309028 522132 309092
rect 66668 302228 66732 302292
rect 66852 302092 66916 302156
rect 521884 302092 521948 302156
rect 67036 299372 67100 299436
rect 504036 297876 504100 297940
rect 67036 289852 67100 289916
rect 522068 289716 522132 289780
rect 69980 288492 70044 288556
rect 82492 284820 82556 284884
rect 504036 283324 504100 283388
rect 504036 280196 504100 280260
rect 521884 280196 521948 280260
rect 67036 280060 67100 280124
rect 21220 278836 21284 278900
rect 521884 273396 521948 273460
rect 522068 272988 522132 273052
rect 66852 270540 66916 270604
rect 522068 270404 522132 270468
rect 501828 269180 501892 269244
rect 502012 269180 502076 269244
rect 529060 263604 529124 263668
rect 521884 260884 521948 260948
rect 66668 260748 66732 260812
rect 67036 260748 67100 260812
rect 81020 255988 81084 256052
rect 501276 255988 501340 256052
rect 501460 255988 501524 256052
rect 504036 254356 504100 254420
rect 521884 253948 521948 254012
rect 503668 253872 503732 253876
rect 503668 253816 503682 253872
rect 503682 253816 503732 253872
rect 503668 253812 503732 253816
rect 522068 253676 522132 253740
rect 67220 251092 67284 251156
rect 522068 251092 522132 251156
rect 67036 250956 67100 251020
rect 79364 245108 79428 245172
rect 67404 241980 67468 242044
rect 67404 241572 67468 241636
rect 521884 241572 521948 241636
rect 67220 240076 67284 240140
rect 502012 238852 502076 238916
rect 521884 234636 521948 234700
rect 522068 234364 522132 234428
rect 503668 232188 503732 232252
rect 503852 231814 503916 231878
rect 501460 229196 501524 229260
rect 501460 228924 501524 228988
rect 501644 228788 501708 228852
rect 501828 228108 501892 228172
rect 507164 228108 507228 228172
rect 82492 227428 82556 227492
rect 511580 227428 511644 227492
rect 522252 227428 522316 227492
rect 67036 222260 67100 222324
rect 521884 222124 521948 222188
rect 501828 220866 501892 220930
rect 501276 219540 501340 219604
rect 501460 219404 501524 219468
rect 67036 215460 67100 215524
rect 66852 215188 66916 215252
rect 522068 212604 522132 212668
rect 522068 212468 522132 212532
rect 501828 206892 501892 206956
rect 502012 206756 502076 206820
rect 67404 205940 67468 206004
rect 77156 205940 77220 206004
rect 521884 206212 521948 206276
rect 61332 205668 61396 205732
rect 75868 205668 75932 205732
rect 501460 205668 501524 205732
rect 70164 205532 70228 205596
rect 67404 205396 67468 205460
rect 77156 205396 77220 205460
rect 75868 204988 75932 205052
rect 78996 204988 79060 205052
rect 66668 201376 66732 201380
rect 66668 201320 66718 201376
rect 66718 201320 66732 201376
rect 66668 201316 66732 201320
rect 521884 199956 521948 200020
rect 501460 198868 501524 198932
rect 66484 195468 66548 195532
rect 503852 194516 503916 194580
rect 504036 192068 504100 192132
rect 66484 191660 66548 191724
rect 521700 190436 521764 190500
rect 75500 187716 75564 187780
rect 502012 187716 502076 187780
rect 502196 187444 502260 187508
rect 504220 186280 504284 186284
rect 504220 186224 504270 186280
rect 504270 186224 504284 186280
rect 504220 186220 504284 186224
rect 504220 185328 504284 185332
rect 504220 185272 504270 185328
rect 504270 185272 504284 185328
rect 504220 185268 504284 185272
rect 503852 184996 503916 185060
rect 501460 183908 501524 183972
rect 501828 182820 501892 182884
rect 502196 182820 502260 182884
rect 531268 181324 531332 181388
rect 503300 181188 503364 181252
rect 522252 181052 522316 181116
rect 531268 180916 531332 180980
rect 504220 176624 504284 176628
rect 504220 176568 504234 176624
rect 504234 176568 504284 176624
rect 504220 176564 504284 176568
rect 521884 176700 521948 176764
rect 521700 176428 521764 176492
rect 504220 175400 504284 175404
rect 504220 175344 504234 175400
rect 504234 175344 504284 175400
rect 504220 175340 504284 175344
rect 503852 175204 503916 175268
rect 67220 173980 67284 174044
rect 503668 174040 503732 174044
rect 503668 173984 503718 174040
rect 503718 173984 503732 174040
rect 503668 173980 503732 173984
rect 521700 173844 521764 173908
rect 503852 165582 503916 165646
rect 521884 164188 521948 164252
rect 521884 157388 521948 157452
rect 521700 157116 521764 157180
rect 72188 155212 72252 155276
rect 501460 154804 501524 154868
rect 501460 151132 501524 151196
rect 521700 147596 521764 147660
rect 522436 147596 522500 147660
rect 66668 144876 66732 144940
rect 66852 144876 66916 144940
rect 66668 137804 66732 137868
rect 67220 137804 67284 137868
rect 522436 138076 522500 138140
rect 501644 137804 501708 137868
rect 522252 137804 522316 137868
rect 522252 135144 522316 135148
rect 522252 135088 522302 135144
rect 522302 135088 522316 135144
rect 522252 135084 522316 135088
rect 501460 126924 501524 126988
rect 521884 125564 521948 125628
rect 502012 122708 502076 122772
rect 501460 121484 501524 121548
rect 501644 121212 501708 121276
rect 501460 119308 501524 119372
rect 521884 118764 521948 118828
rect 522068 118492 522132 118556
rect 522068 115772 522132 115836
rect 512684 114548 512748 114612
rect 67036 114472 67100 114476
rect 67036 114416 67086 114472
rect 67086 114416 67100 114472
rect 67036 114412 67100 114416
rect 67036 113188 67100 113252
rect 521884 106252 521948 106316
rect 67036 103396 67100 103460
rect 82860 102444 82924 102508
rect 144868 102580 144932 102644
rect 144868 102308 144932 102372
rect 502380 102716 502444 102780
rect 497780 102580 497844 102644
rect 500908 102580 500972 102644
rect 501276 102580 501340 102644
rect 492812 102444 492876 102508
rect 493732 102444 493796 102508
rect 492996 102308 493060 102372
rect 499988 102308 500052 102372
rect 487108 102172 487172 102236
rect 492812 102172 492876 102236
rect 492996 102036 493060 102100
rect 495204 102172 495268 102236
rect 500172 102172 500236 102236
rect 489132 101764 489196 101828
rect 241468 101628 241532 101692
rect 251036 101628 251100 101692
rect 493732 101356 493796 101420
rect 395844 100948 395908 101012
rect 402836 100948 402900 101012
rect 403756 100948 403820 101012
rect 412404 100948 412468 101012
rect 481588 100948 481652 101012
rect 495204 100948 495268 101012
rect 504588 100948 504652 101012
rect 507164 100948 507228 101012
rect 68876 100676 68940 100740
rect 486372 100676 486436 100740
rect 498884 100676 498948 100740
rect 231900 100268 231964 100332
rect 241284 100268 241348 100332
rect 270540 100268 270604 100332
rect 273852 100268 273916 100332
rect 347820 100268 347884 100332
rect 351132 100268 351196 100332
rect 504220 99044 504284 99108
rect 83228 98908 83292 98972
rect 81572 98772 81636 98836
rect 521884 98772 521948 98836
rect 72372 98636 72436 98700
rect 519492 97820 519556 97884
rect 499804 97140 499868 97204
rect 487844 96596 487908 96660
rect 489868 96596 489932 96660
rect 71084 96460 71148 96524
rect 492812 95916 492876 95980
rect 78260 94420 78324 94484
rect 496492 93876 496556 93940
rect 496492 93604 496556 93668
rect 81020 93060 81084 93124
rect 501276 92380 501340 92444
rect 501092 92244 501156 92308
rect 79364 90476 79428 90540
rect 509188 90340 509252 90404
rect 67036 89720 67100 89724
rect 67036 89664 67086 89720
rect 67086 89664 67100 89720
rect 67036 89660 67100 89664
rect 506428 87756 506492 87820
rect 500540 87680 500604 87684
rect 500540 87624 500554 87680
rect 500554 87624 500604 87680
rect 500540 87620 500604 87624
rect 79732 87484 79796 87548
rect 500172 87348 500236 87412
rect 500724 87348 500788 87412
rect 511212 86940 511276 87004
rect 83412 86260 83476 86324
rect 505692 86260 505756 86324
rect 81388 86124 81452 86188
rect 496492 85580 496556 85644
rect 496492 85308 496556 85372
rect 510660 80004 510724 80068
rect 503852 79324 503916 79388
rect 74028 77828 74092 77892
rect 499620 77420 499684 77484
rect 499436 77284 499500 77348
rect 499436 75108 499500 75172
rect 67220 72448 67284 72452
rect 67220 72392 67270 72448
rect 67270 72392 67284 72448
rect 67220 72388 67284 72392
rect 505876 72388 505940 72452
rect 78444 71300 78508 71364
rect 501644 71164 501708 71228
rect 79548 71028 79612 71092
rect 76236 69532 76300 69596
rect 67220 67688 67284 67692
rect 67220 67632 67270 67688
rect 67270 67632 67284 67688
rect 67220 67628 67284 67632
rect 499068 67688 499132 67692
rect 499068 67632 499118 67688
rect 499118 67632 499132 67688
rect 499068 67628 499132 67632
rect 499068 66948 499132 67012
rect 78076 66812 78140 66876
rect 67220 60828 67284 60892
rect 500908 60828 500972 60892
rect 67036 60556 67100 60620
rect 501092 60556 501156 60620
rect 499252 60072 499316 60076
rect 499252 60016 499266 60072
rect 499266 60016 499316 60072
rect 499252 60012 499316 60016
rect 81756 59876 81820 59940
rect 67036 57896 67100 57900
rect 67036 57840 67086 57896
rect 67086 57840 67100 57896
rect 67036 57836 67100 57840
rect 500356 57156 500420 57220
rect 499252 55176 499316 55180
rect 499252 55120 499266 55176
rect 499266 55120 499316 55176
rect 499252 55116 499316 55120
rect 74212 53076 74276 53140
rect 502748 51716 502812 51780
rect 67036 50960 67100 50964
rect 67036 50904 67086 50960
rect 67086 50904 67100 50960
rect 67036 50900 67100 50904
rect 486188 50356 486252 50420
rect 502564 50220 502628 50284
rect 81204 47500 81268 47564
rect 506612 46140 506676 46204
rect 499252 45792 499316 45796
rect 499252 45736 499266 45792
rect 499266 45736 499316 45792
rect 499252 45732 499316 45736
rect 496492 45460 496556 45524
rect 499252 45520 499316 45524
rect 499252 45464 499266 45520
rect 499266 45464 499316 45520
rect 499252 45460 499316 45464
rect 501092 45460 501156 45524
rect 506796 44780 506860 44844
rect 496308 40760 496372 40764
rect 496308 40704 496358 40760
rect 496358 40704 496372 40760
rect 496308 40700 496372 40704
rect 499252 40760 499316 40764
rect 499252 40704 499266 40760
rect 499266 40704 499316 40760
rect 499252 40700 499316 40704
rect 505508 36484 505572 36548
rect 64092 35804 64156 35868
rect 74396 35124 74460 35188
rect 509372 30908 509436 30972
rect 516732 29004 516796 29068
rect 498332 28868 498396 28932
rect 504036 26828 504100 26892
rect 70900 24108 70964 24172
rect 498516 21116 498580 21180
rect 496308 12548 496372 12612
rect 496124 12276 496188 12340
rect 75500 11732 75564 11796
rect 495940 11596 496004 11660
rect 66668 9284 66732 9348
rect 491340 9284 491404 9348
rect 497412 9012 497476 9076
rect 498516 8876 498580 8940
rect 494836 7516 494900 7580
rect 495572 6700 495636 6764
rect 507900 6564 507964 6628
rect 492628 6428 492692 6492
rect 72188 6292 72252 6356
rect 496860 6292 496924 6356
rect 69980 6156 70044 6220
rect 222148 6020 222212 6084
rect 230428 6020 230492 6084
rect 239996 6020 240060 6084
rect 249748 6020 249812 6084
rect 288388 6020 288452 6084
rect 297956 6020 298020 6084
rect 384988 6020 385052 6084
rect 405780 6020 405844 6084
rect 153148 5884 153212 5948
rect 211108 5944 211172 5948
rect 211108 5888 211122 5944
rect 211122 5888 211172 5944
rect 211108 5884 211172 5888
rect 77156 5748 77220 5812
rect 239996 5748 240060 5812
rect 249748 5748 249812 5812
rect 260972 5748 261036 5812
rect 269068 5748 269132 5812
rect 288388 5748 288452 5812
rect 297956 5748 298020 5812
rect 307708 5748 307772 5812
rect 317276 5748 317340 5812
rect 153148 5612 153212 5676
rect 260788 5612 260852 5676
rect 360148 5748 360212 5812
rect 360332 5748 360396 5812
rect 365668 5748 365732 5812
rect 384988 5748 385052 5812
rect 405780 5612 405844 5676
rect 456748 5748 456812 5812
rect 456932 5748 456996 5812
rect 222148 5476 222212 5540
rect 230428 5476 230492 5540
rect 269068 5476 269132 5540
rect 307708 5476 307772 5540
rect 317276 5476 317340 5540
rect 365668 5476 365732 5540
rect 535500 5748 535564 5812
rect 211108 5340 211172 5404
rect 499252 4796 499316 4860
rect 169524 3980 169588 4044
rect 488580 3980 488644 4044
rect 535500 3980 535564 4044
rect 490236 3844 490300 3908
rect 75132 3708 75196 3772
rect 75684 3708 75748 3772
rect 486004 3708 486068 3772
rect 491892 3572 491956 3636
rect 67404 3436 67468 3500
rect 72556 3436 72620 3500
rect 501460 3436 501524 3500
rect 466132 2756 466196 2820
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 10182 452573 10242 485742
rect 11604 481254 12204 516698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 10179 452572 10245 452573
rect 10179 452508 10180 452572
rect 10244 452508 10245 452572
rect 10179 452507 10245 452508
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 21219 278900 21285 278901
rect 21219 278836 21220 278900
rect 21284 278836 21285 278900
rect 21219 278835 21285 278836
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 21222 206498 21282 278835
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 27478 485893 27538 487102
rect 27475 485892 27541 485893
rect 27475 485828 27476 485892
rect 27540 485828 27541 485892
rect 27475 485827 27541 485828
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 463254 30204 498698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 46795 487252 46861 487253
rect 46795 487188 46796 487252
rect 46860 487188 46861 487252
rect 46795 487187 46861 487188
rect 46798 484618 46858 487187
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 68875 700364 68941 700365
rect 68875 700300 68876 700364
rect 68940 700300 68941 700364
rect 68875 700299 68941 700300
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 61334 205733 61394 206262
rect 61331 205732 61397 205733
rect 61331 205668 61332 205732
rect 61396 205668 61397 205732
rect 61331 205667 61397 205668
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 64094 35869 64154 605422
rect 65604 571254 66204 606698
rect 67403 604892 67469 604893
rect 67403 604828 67404 604892
rect 67468 604828 67469 604892
rect 67403 604827 67469 604828
rect 67002 598710 67282 598770
rect 67222 591970 67282 598710
rect 66854 591910 67282 591970
rect 66854 582453 66914 591910
rect 66851 582452 66917 582453
rect 66851 582388 66852 582452
rect 66916 582388 66917 582452
rect 66851 582387 66917 582388
rect 67035 582180 67101 582181
rect 67035 582116 67036 582180
rect 67100 582116 67101 582180
rect 67035 582115 67101 582116
rect 67038 578237 67098 582115
rect 67035 578236 67101 578237
rect 67035 578172 67036 578236
rect 67100 578172 67101 578236
rect 67035 578171 67101 578172
rect 67035 572660 67101 572661
rect 67035 572596 67036 572660
rect 67100 572596 67101 572660
rect 67035 572595 67101 572596
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 67038 562730 67098 572595
rect 66854 562670 67098 562730
rect 66854 553485 66914 562670
rect 66851 553484 66917 553485
rect 66851 553420 66852 553484
rect 66916 553420 66917 553484
rect 66851 553419 66917 553420
rect 67035 553212 67101 553213
rect 67035 553148 67036 553212
rect 67100 553148 67101 553212
rect 67035 553147 67101 553148
rect 67038 543965 67098 553147
rect 67035 543964 67101 543965
rect 67035 543900 67036 543964
rect 67100 543900 67101 543964
rect 67035 543899 67101 543900
rect 67035 543556 67101 543557
rect 67035 543492 67036 543556
rect 67100 543492 67101 543556
rect 67035 543491 67101 543492
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 67038 534309 67098 543491
rect 67035 534308 67101 534309
rect 67035 534244 67036 534308
rect 67100 534244 67101 534308
rect 67035 534243 67101 534244
rect 67035 531452 67101 531453
rect 67035 531388 67036 531452
rect 67100 531388 67101 531452
rect 67035 531387 67101 531388
rect 67038 524789 67098 531387
rect 67035 524788 67101 524789
rect 67035 524724 67036 524788
rect 67100 524724 67101 524788
rect 67035 524723 67101 524724
rect 66667 524244 66733 524245
rect 66667 524180 66668 524244
rect 66732 524180 66733 524244
rect 66667 524179 66733 524180
rect 66670 521661 66730 524179
rect 66667 521660 66733 521661
rect 66667 521596 66668 521660
rect 66732 521596 66733 521660
rect 66667 521595 66733 521596
rect 66483 512140 66549 512141
rect 66483 512076 66484 512140
rect 66548 512076 66549 512140
rect 66483 512075 66549 512076
rect 66486 510509 66546 512075
rect 66483 510508 66549 510509
rect 66483 510444 66484 510508
rect 66548 510444 66549 510508
rect 66483 510443 66549 510444
rect 67035 500988 67101 500989
rect 67035 500924 67036 500988
rect 67100 500924 67101 500988
rect 67035 500923 67101 500924
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 67038 491197 67098 500923
rect 67035 491196 67101 491197
rect 67035 491132 67036 491196
rect 67100 491132 67101 491196
rect 67035 491131 67101 491132
rect 67035 483716 67101 483717
rect 67035 483652 67036 483716
rect 67100 483652 67101 483716
rect 67035 483651 67101 483652
rect 67038 478821 67098 483651
rect 67035 478820 67101 478821
rect 67035 478756 67036 478820
rect 67100 478756 67101 478820
rect 67035 478755 67101 478756
rect 67035 469436 67101 469437
rect 67035 469372 67036 469436
rect 67100 469372 67101 469436
rect 67035 469371 67101 469372
rect 67038 469165 67098 469371
rect 67035 469164 67101 469165
rect 67035 469100 67036 469164
rect 67100 469100 67101 469164
rect 67035 469099 67101 469100
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 66851 459644 66917 459645
rect 66851 459580 66852 459644
rect 66916 459580 66917 459644
rect 66851 459579 66917 459580
rect 66854 455970 66914 459579
rect 66854 455910 67098 455970
rect 67038 446453 67098 455910
rect 67035 446452 67101 446453
rect 67035 446388 67036 446452
rect 67100 446388 67101 446452
rect 67035 446387 67101 446388
rect 66667 434756 66733 434757
rect 66667 434692 66668 434756
rect 66732 434692 66733 434756
rect 66667 434691 66733 434692
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 66670 426730 66730 434691
rect 67406 434621 67466 604827
rect 67403 434620 67469 434621
rect 67403 434556 67404 434620
rect 67468 434556 67469 434620
rect 67403 434555 67469 434556
rect 67403 429860 67469 429861
rect 67403 429796 67404 429860
rect 67468 429796 67469 429860
rect 67403 429795 67469 429796
rect 66670 426670 67282 426730
rect 67222 398989 67282 426670
rect 67219 398988 67285 398989
rect 67219 398924 67220 398988
rect 67284 398924 67285 398988
rect 67219 398923 67285 398924
rect 66851 396132 66917 396133
rect 66851 396068 66852 396132
rect 66916 396068 66917 396132
rect 66851 396067 66917 396068
rect 66854 394637 66914 396067
rect 66851 394636 66917 394637
rect 66851 394572 66852 394636
rect 66916 394572 66917 394636
rect 66851 394571 66917 394572
rect 67035 394500 67101 394501
rect 67035 394436 67036 394500
rect 67100 394436 67101 394500
rect 67035 394435 67101 394436
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 67038 383621 67098 394435
rect 67035 383620 67101 383621
rect 67035 383556 67036 383620
rect 67100 383556 67101 383620
rect 67035 383555 67101 383556
rect 67219 374100 67285 374101
rect 67219 374036 67220 374100
rect 67284 374036 67285 374100
rect 67219 374035 67285 374036
rect 67222 373829 67282 374035
rect 66851 373828 66917 373829
rect 66851 373764 66852 373828
rect 66916 373764 66917 373828
rect 66851 373763 66917 373764
rect 67219 373828 67285 373829
rect 67219 373764 67220 373828
rect 67284 373764 67285 373828
rect 67219 373763 67285 373764
rect 66854 368930 66914 373763
rect 66854 368870 67282 368930
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 67222 350709 67282 368870
rect 67219 350708 67285 350709
rect 67219 350644 67220 350708
rect 67284 350644 67285 350708
rect 67219 350643 67285 350644
rect 66851 350572 66917 350573
rect 66851 350508 66852 350572
rect 66916 350508 66917 350572
rect 66851 350507 66917 350508
rect 66854 341053 66914 350507
rect 66851 341052 66917 341053
rect 66851 340988 66852 341052
rect 66916 340988 66917 341052
rect 66851 340987 66917 340988
rect 67035 340780 67101 340781
rect 67035 340716 67036 340780
rect 67100 340716 67101 340780
rect 67035 340715 67101 340716
rect 67038 336701 67098 340715
rect 67035 336700 67101 336701
rect 67035 336636 67036 336700
rect 67100 336636 67101 336700
rect 67035 336635 67101 336636
rect 67406 328405 67466 429795
rect 67403 328404 67469 328405
rect 67403 328340 67404 328404
rect 67468 328340 67469 328404
rect 67403 328339 67469 328340
rect 66667 327180 66733 327181
rect 66667 327116 66668 327180
rect 66732 327116 66733 327180
rect 66667 327115 66733 327116
rect 66670 321330 66730 327115
rect 67403 323644 67469 323645
rect 67403 323580 67404 323644
rect 67468 323580 67469 323644
rect 67403 323579 67469 323580
rect 66670 321270 67098 321330
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 67038 312085 67098 321270
rect 67035 312084 67101 312085
rect 67035 312020 67036 312084
rect 67100 312020 67101 312084
rect 67035 312019 67101 312020
rect 66851 311812 66917 311813
rect 66851 311748 66852 311812
rect 66916 311748 66917 311812
rect 66851 311747 66917 311748
rect 66854 309090 66914 311747
rect 66670 309030 66914 309090
rect 66670 302293 66730 309030
rect 66667 302292 66733 302293
rect 66667 302228 66668 302292
rect 66732 302228 66733 302292
rect 66667 302227 66733 302228
rect 66851 302156 66917 302157
rect 66851 302092 66852 302156
rect 66916 302092 66917 302156
rect 66851 302091 66917 302092
rect 66854 300250 66914 302091
rect 66854 300190 67052 300250
rect 66992 299570 67052 300190
rect 66992 299510 67098 299570
rect 67038 299437 67098 299510
rect 67035 299436 67101 299437
rect 67035 299372 67036 299436
rect 67100 299372 67101 299436
rect 67035 299371 67101 299372
rect 67035 289916 67101 289917
rect 67035 289852 67036 289916
rect 67100 289852 67101 289916
rect 67035 289851 67101 289852
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 67038 280125 67098 289851
rect 67035 280124 67101 280125
rect 67035 280060 67036 280124
rect 67100 280060 67101 280124
rect 67035 280059 67101 280060
rect 66851 270604 66917 270605
rect 66851 270540 66852 270604
rect 66916 270540 66917 270604
rect 66851 270539 66917 270540
rect 66854 264210 66914 270539
rect 66486 264150 66914 264210
rect 66486 263530 66546 264150
rect 66486 263470 66730 263530
rect 66670 260813 66730 263470
rect 66667 260812 66733 260813
rect 66667 260748 66668 260812
rect 66732 260748 66733 260812
rect 66667 260747 66733 260748
rect 67035 260812 67101 260813
rect 67035 260748 67036 260812
rect 67100 260748 67101 260812
rect 67035 260747 67101 260748
rect 67038 252650 67098 260747
rect 67038 252590 67282 252650
rect 67222 251157 67282 252590
rect 67219 251156 67285 251157
rect 67219 251092 67220 251156
rect 67284 251092 67285 251156
rect 67219 251091 67285 251092
rect 67035 251020 67101 251021
rect 67035 250956 67036 251020
rect 67100 250956 67101 251020
rect 67035 250955 67101 250956
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 67038 241770 67098 250955
rect 67406 242045 67466 323579
rect 67403 242044 67469 242045
rect 67403 241980 67404 242044
rect 67468 241980 67469 242044
rect 67403 241979 67469 241980
rect 67038 241710 67282 241770
rect 67222 240141 67282 241710
rect 67403 241636 67469 241637
rect 67403 241572 67404 241636
rect 67468 241572 67469 241636
rect 67403 241571 67469 241572
rect 67219 240140 67285 240141
rect 67219 240076 67220 240140
rect 67284 240076 67285 240140
rect 67219 240075 67285 240076
rect 67035 222324 67101 222325
rect 67035 222260 67036 222324
rect 67100 222260 67101 222324
rect 67035 222259 67101 222260
rect 67038 215525 67098 222259
rect 67035 215524 67101 215525
rect 67035 215460 67036 215524
rect 67100 215460 67101 215524
rect 67035 215459 67101 215460
rect 66851 215252 66917 215253
rect 66851 215188 66852 215252
rect 66916 215188 66917 215252
rect 66851 215187 66917 215188
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 66854 205730 66914 215187
rect 67406 206005 67466 241571
rect 67403 206004 67469 206005
rect 67403 205940 67404 206004
rect 67468 205940 67469 206004
rect 67403 205939 67469 205940
rect 66670 205670 66914 205730
rect 66670 201381 66730 205670
rect 67403 205460 67469 205461
rect 67403 205396 67404 205460
rect 67468 205396 67469 205460
rect 67403 205395 67469 205396
rect 66667 201380 66733 201381
rect 66667 201316 66668 201380
rect 66732 201316 66733 201380
rect 66667 201315 66733 201316
rect 66483 195532 66549 195533
rect 66483 195468 66484 195532
rect 66548 195468 66549 195532
rect 66483 195467 66549 195468
rect 66486 191725 66546 195467
rect 66483 191724 66549 191725
rect 66483 191660 66484 191724
rect 66548 191660 66549 191724
rect 66483 191659 66549 191660
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 67219 174044 67285 174045
rect 67219 173980 67220 174044
rect 67284 173980 67285 174044
rect 67219 173979 67285 173980
rect 67222 166970 67282 173979
rect 67038 166910 67282 166970
rect 67038 157450 67098 166910
rect 66854 157390 67098 157450
rect 66854 144941 66914 157390
rect 66667 144940 66733 144941
rect 66667 144876 66668 144940
rect 66732 144876 66733 144940
rect 66667 144875 66733 144876
rect 66851 144940 66917 144941
rect 66851 144876 66852 144940
rect 66916 144876 66917 144940
rect 66851 144875 66917 144876
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 66670 137869 66730 144875
rect 66667 137868 66733 137869
rect 66667 137804 66668 137868
rect 66732 137804 66733 137868
rect 66667 137803 66733 137804
rect 67219 137868 67285 137869
rect 67219 137804 67220 137868
rect 67284 137804 67285 137868
rect 67219 137803 67285 137804
rect 67222 128210 67282 137803
rect 67038 128150 67282 128210
rect 67038 114477 67098 128150
rect 67035 114476 67101 114477
rect 67035 114412 67036 114476
rect 67100 114412 67101 114476
rect 67035 114411 67101 114412
rect 67035 113252 67101 113253
rect 67035 113188 67036 113252
rect 67100 113188 67101 113252
rect 67035 113187 67101 113188
rect 67038 103461 67098 113187
rect 67035 103460 67101 103461
rect 67035 103396 67036 103460
rect 67100 103396 67101 103460
rect 67035 103395 67101 103396
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 67035 89724 67101 89725
rect 67035 89660 67036 89724
rect 67100 89660 67101 89724
rect 67035 89659 67101 89660
rect 67038 77890 67098 89659
rect 67038 77830 67282 77890
rect 67222 72453 67282 77830
rect 67219 72452 67285 72453
rect 67219 72388 67220 72452
rect 67284 72388 67285 72452
rect 67219 72387 67285 72388
rect 67219 67692 67285 67693
rect 67219 67628 67220 67692
rect 67284 67628 67285 67692
rect 67219 67627 67285 67628
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 64091 35868 64157 35869
rect 64091 35804 64092 35868
rect 64156 35804 64157 35868
rect 64091 35803 64157 35804
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 31254 66204 66698
rect 67222 60893 67282 67627
rect 67219 60892 67285 60893
rect 67219 60828 67220 60892
rect 67284 60828 67285 60892
rect 67219 60827 67285 60828
rect 67035 60620 67101 60621
rect 67035 60556 67036 60620
rect 67100 60556 67101 60620
rect 67035 60555 67101 60556
rect 67038 57901 67098 60555
rect 67035 57900 67101 57901
rect 67035 57836 67036 57900
rect 67100 57836 67101 57900
rect 67035 57835 67101 57836
rect 67035 50964 67101 50965
rect 67035 50900 67036 50964
rect 67100 50900 67101 50964
rect 67035 50899 67101 50900
rect 67038 41170 67098 50899
rect 66854 41110 67098 41170
rect 66854 32330 66914 41110
rect 66486 32270 66914 32330
rect 66486 31650 66546 32270
rect 66486 31590 66730 31650
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 66670 22130 66730 31590
rect 66670 22070 66914 22130
rect 66854 12610 66914 22070
rect 66670 12550 66914 12610
rect 66670 9349 66730 12550
rect 66667 9348 66733 9349
rect 66667 9284 66668 9348
rect 66732 9284 66733 9348
rect 66667 9283 66733 9284
rect 67406 3501 67466 205395
rect 68878 100741 68938 700299
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 70163 673572 70229 673573
rect 70163 673508 70164 673572
rect 70228 673508 70229 673572
rect 70163 673507 70229 673508
rect 69979 288556 70045 288557
rect 69979 288492 69980 288556
rect 70044 288492 70045 288556
rect 69979 288491 70045 288492
rect 68875 100740 68941 100741
rect 68875 100676 68876 100740
rect 68940 100676 68941 100740
rect 68875 100675 68941 100676
rect 69982 6221 70042 288491
rect 70166 205597 70226 673507
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 70899 603668 70965 603669
rect 70899 603604 70900 603668
rect 70964 603604 70965 603668
rect 70899 603603 70965 603604
rect 70163 205596 70229 205597
rect 70163 205532 70164 205596
rect 70228 205532 70229 205596
rect 70163 205531 70229 205532
rect 70902 24173 70962 603603
rect 72371 603396 72437 603397
rect 72371 603332 72372 603396
rect 72436 603332 72437 603396
rect 72371 603331 72437 603332
rect 71083 365804 71149 365805
rect 71083 365740 71084 365804
rect 71148 365740 71149 365804
rect 71083 365739 71149 365740
rect 71086 96525 71146 365739
rect 72187 155276 72253 155277
rect 72187 155212 72188 155276
rect 72252 155212 72253 155276
rect 72187 155211 72253 155212
rect 71083 96524 71149 96525
rect 71083 96460 71084 96524
rect 71148 96460 71149 96524
rect 71083 96459 71149 96460
rect 70899 24172 70965 24173
rect 70899 24108 70900 24172
rect 70964 24108 70965 24172
rect 70899 24107 70965 24108
rect 72190 6357 72250 155211
rect 72374 98701 72434 603331
rect 72555 602172 72621 602173
rect 72555 602108 72556 602172
rect 72620 602108 72621 602172
rect 72555 602107 72621 602108
rect 72371 98700 72437 98701
rect 72371 98636 72372 98700
rect 72436 98636 72437 98700
rect 72371 98635 72437 98636
rect 72187 6356 72253 6357
rect 72187 6292 72188 6356
rect 72252 6292 72253 6356
rect 72187 6291 72253 6292
rect 69979 6220 70045 6221
rect 69979 6156 69980 6220
rect 70044 6156 70045 6220
rect 69979 6155 70045 6156
rect 72558 3501 72618 602107
rect 72804 578454 73404 613898
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 75131 602036 75197 602037
rect 75131 601972 75132 602036
rect 75196 601972 75197 602036
rect 75131 601971 75197 601972
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 74211 543828 74277 543829
rect 74211 543764 74212 543828
rect 74276 543764 74277 543828
rect 74211 543763 74277 543764
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 74027 423740 74093 423741
rect 74027 423676 74028 423740
rect 74092 423676 74093 423740
rect 74027 423675 74093 423676
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 74030 77893 74090 423675
rect 74027 77892 74093 77893
rect 74027 77828 74028 77892
rect 74092 77828 74093 77892
rect 74027 77827 74093 77828
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 74214 53141 74274 543763
rect 74395 541108 74461 541109
rect 74395 541044 74396 541108
rect 74460 541044 74461 541108
rect 74395 541043 74461 541044
rect 74211 53140 74277 53141
rect 74211 53076 74212 53140
rect 74276 53076 74277 53140
rect 74211 53075 74277 53076
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 67403 3500 67469 3501
rect 67403 3436 67404 3500
rect 67468 3436 67469 3500
rect 67403 3435 67469 3436
rect 72555 3500 72621 3501
rect 72555 3436 72556 3500
rect 72620 3436 72621 3500
rect 72555 3435 72621 3436
rect 72804 2454 73404 37898
rect 74398 35189 74458 541043
rect 74395 35188 74461 35189
rect 74395 35124 74396 35188
rect 74460 35124 74461 35188
rect 74395 35123 74461 35124
rect 75134 3773 75194 601971
rect 75867 601356 75933 601357
rect 75867 601292 75868 601356
rect 75932 601292 75933 601356
rect 75867 601291 75933 601292
rect 75870 601085 75930 601291
rect 75867 601084 75933 601085
rect 75867 601020 75868 601084
rect 75932 601020 75933 601084
rect 75867 601019 75933 601020
rect 75683 600132 75749 600133
rect 75683 600068 75684 600132
rect 75748 600068 75749 600132
rect 75683 600067 75749 600068
rect 75499 187780 75565 187781
rect 75499 187716 75500 187780
rect 75564 187716 75565 187780
rect 75499 187715 75565 187716
rect 75502 11797 75562 187715
rect 75499 11796 75565 11797
rect 75499 11732 75500 11796
rect 75564 11732 75565 11796
rect 75499 11731 75565 11732
rect 75686 3773 75746 600067
rect 76404 582054 77004 617498
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 78443 588436 78509 588437
rect 78443 588372 78444 588436
rect 78508 588372 78509 588436
rect 78443 588371 78509 588372
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 77155 551988 77221 551989
rect 77155 551924 77156 551988
rect 77220 551924 77221 551988
rect 77155 551923 77221 551924
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76235 537300 76301 537301
rect 76235 537236 76236 537300
rect 76300 537236 76301 537300
rect 76235 537235 76301 537236
rect 75867 205732 75933 205733
rect 75867 205668 75868 205732
rect 75932 205668 75933 205732
rect 75867 205667 75933 205668
rect 75870 205053 75930 205667
rect 75867 205052 75933 205053
rect 75867 204988 75868 205052
rect 75932 204988 75933 205052
rect 75867 204987 75933 204988
rect 76238 69597 76298 537235
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 77158 206005 77218 551923
rect 78259 548452 78325 548453
rect 78259 548388 78260 548452
rect 78324 548388 78325 548452
rect 78259 548387 78325 548388
rect 78075 365668 78141 365669
rect 78075 365604 78076 365668
rect 78140 365604 78141 365668
rect 78075 365603 78141 365604
rect 77155 206004 77221 206005
rect 77155 205940 77156 206004
rect 77220 205940 77221 206004
rect 77155 205939 77221 205940
rect 77155 205460 77221 205461
rect 77155 205396 77156 205460
rect 77220 205396 77221 205460
rect 77155 205395 77221 205396
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76235 69596 76301 69597
rect 76235 69532 76236 69596
rect 76300 69532 76301 69596
rect 76235 69531 76301 69532
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 77158 5813 77218 205395
rect 78078 66877 78138 365603
rect 78262 94485 78322 548387
rect 78259 94484 78325 94485
rect 78259 94420 78260 94484
rect 78324 94420 78325 94484
rect 78259 94419 78325 94420
rect 78446 71365 78506 588371
rect 80004 585654 80604 621098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 82859 603260 82925 603261
rect 82859 603196 82860 603260
rect 82924 603196 82925 603260
rect 82859 603195 82925 603196
rect 82862 600269 82922 603195
rect 82859 600268 82925 600269
rect 82859 600204 82860 600268
rect 82924 600204 82925 600268
rect 82859 600203 82925 600204
rect 80835 600132 80901 600133
rect 80835 600068 80836 600132
rect 80900 600068 80901 600132
rect 80835 600067 80901 600068
rect 80838 598858 80898 600067
rect 83230 596050 83290 604062
rect 83604 602000 84204 624698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 86907 604076 86973 604077
rect 86907 604012 86908 604076
rect 86972 604012 86973 604076
rect 86907 604011 86973 604012
rect 86910 603805 86970 604011
rect 86907 603804 86973 603805
rect 86907 603740 86908 603804
rect 86972 603740 86973 603804
rect 86907 603739 86973 603740
rect 89667 603532 89733 603533
rect 89667 603468 89668 603532
rect 89732 603468 89733 603532
rect 89667 603467 89733 603468
rect 86907 601220 86973 601221
rect 86907 601156 86908 601220
rect 86972 601156 86973 601220
rect 86907 601155 86973 601156
rect 86910 600949 86970 601155
rect 86907 600948 86973 600949
rect 86907 600884 86908 600948
rect 86972 600884 86973 600948
rect 86907 600883 86973 600884
rect 89670 600133 89730 603467
rect 90804 602000 91404 631898
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 602000 95004 635498
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 602000 98604 603098
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 602000 102204 606698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 602000 109404 613898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 109723 605572 109789 605573
rect 109723 605508 109724 605572
rect 109788 605508 109789 605572
rect 109723 605507 109789 605508
rect 109726 604978 109786 605507
rect 112404 602000 113004 617498
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 602000 116604 621098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 118923 606116 118989 606117
rect 118923 606052 118924 606116
rect 118988 606052 118989 606116
rect 118923 606051 118989 606052
rect 118926 605658 118986 606051
rect 119604 602000 120204 624698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 602000 127404 631898
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 128675 606116 128741 606117
rect 128675 606052 128676 606116
rect 128740 606052 128741 606116
rect 128675 606051 128741 606052
rect 128678 605658 128738 606051
rect 130404 602000 131004 635498
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 602000 134604 603098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 602000 138204 606698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 138427 606116 138493 606117
rect 138427 606052 138428 606116
rect 138492 606052 138493 606116
rect 138427 606051 138493 606052
rect 138430 605658 138490 606051
rect 144804 602000 145404 613898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 602000 149004 617498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 602000 152604 621098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 153147 604076 153213 604077
rect 153147 604012 153148 604076
rect 153212 604012 153213 604076
rect 153147 604011 153213 604012
rect 153150 603805 153210 604011
rect 153147 603804 153213 603805
rect 153147 603740 153148 603804
rect 153212 603740 153213 603804
rect 153147 603739 153213 603740
rect 155604 602000 156204 624698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 157195 606116 157261 606117
rect 157195 606052 157196 606116
rect 157260 606052 157261 606116
rect 157195 606051 157261 606052
rect 157198 605658 157258 606051
rect 157934 604213 157994 604742
rect 157931 604212 157997 604213
rect 157931 604148 157932 604212
rect 157996 604148 157997 604212
rect 157931 604147 157997 604148
rect 162804 602000 163404 631898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 602000 167004 635498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 602000 170604 603098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 602000 174204 606698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 183507 674116 183573 674117
rect 183507 674052 183508 674116
rect 183572 674052 183573 674116
rect 183507 674051 183573 674052
rect 183510 673845 183570 674051
rect 183507 673844 183573 673845
rect 183507 673780 183508 673844
rect 183572 673780 183573 673844
rect 183507 673779 183573 673780
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 176883 606116 176949 606117
rect 176883 606052 176884 606116
rect 176948 606052 176949 606116
rect 176883 606051 176949 606052
rect 176886 605658 176946 606051
rect 180804 602000 181404 613898
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 602000 185004 617498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 602000 188604 621098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 602000 192204 624698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 195835 606116 195901 606117
rect 195835 606052 195836 606116
rect 195900 606052 195901 606116
rect 195835 606051 195901 606052
rect 196571 606116 196637 606117
rect 196571 606052 196572 606116
rect 196636 606052 196637 606116
rect 196571 606051 196637 606052
rect 195838 605658 195898 606051
rect 196574 605658 196634 606051
rect 198804 602000 199404 631898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 602000 203004 635498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 205186 604150 205686 604210
rect 206004 603654 206604 639098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 207059 606116 207125 606117
rect 207059 606052 207060 606116
rect 207124 606052 207125 606116
rect 207059 606051 207125 606052
rect 207062 604978 207122 606051
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 602000 206604 603098
rect 209604 602000 210204 606698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 602000 217404 613898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 602000 221004 617498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 602000 224604 621098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 602000 228204 624698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 602000 235404 631898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 235947 606252 236013 606253
rect 235947 606188 235948 606252
rect 236012 606188 236013 606252
rect 235947 606187 236013 606188
rect 235950 605658 236010 606187
rect 238404 602000 239004 635498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 244411 606252 244477 606253
rect 244411 606188 244412 606252
rect 244476 606188 244477 606252
rect 244411 606187 244477 606188
rect 244414 605658 244474 606187
rect 243826 604150 244326 604210
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 602000 242604 603098
rect 245604 602000 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 602000 253404 613898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 253979 606252 254045 606253
rect 253979 606188 253980 606252
rect 254044 606188 254045 606252
rect 253979 606187 254045 606188
rect 253982 605658 254042 606187
rect 256404 602000 257004 617498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 602000 260604 621098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 602000 264204 624698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 602000 271404 631898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 272931 606252 272997 606253
rect 272931 606188 272932 606252
rect 272996 606188 272997 606252
rect 272931 606187 272997 606188
rect 273299 606252 273365 606253
rect 273299 606188 273300 606252
rect 273364 606188 273365 606252
rect 273299 606187 273365 606188
rect 272934 605658 272994 606187
rect 273302 605658 273362 606187
rect 274404 602000 275004 635498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 602000 278604 603098
rect 281604 602000 282204 606698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 602000 289404 613898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 602000 293004 617498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 602000 296604 621098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 602000 300204 624698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 301786 604150 302286 604210
rect 306804 602000 307404 631898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 602000 311004 635498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 602000 314604 603098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 602000 318204 606698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 321106 604150 321606 604210
rect 324804 602000 325404 613898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 602000 329004 617498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 602000 332604 621098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 602000 336204 624698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 340426 604150 340926 604210
rect 342804 602000 343404 631898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 602000 347004 635498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 602000 350604 603098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 602000 354204 606698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 359746 604150 360246 604210
rect 360804 602000 361404 613898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 602000 365004 617498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 602000 368604 621098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 602000 372204 624698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 602000 379404 631898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 602000 383004 635498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 384987 603940 385053 603941
rect 384987 603876 384988 603940
rect 385052 603876 385053 603940
rect 384987 603875 385053 603876
rect 384990 603669 385050 603875
rect 384987 603668 385053 603669
rect 384987 603604 384988 603668
rect 385052 603604 385053 603668
rect 384987 603603 385053 603604
rect 386004 603654 386604 639098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 602000 386604 603098
rect 389604 602000 390204 606698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 602000 397404 613898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 602000 401004 617498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 602000 404604 621098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 602000 408204 624698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 602000 415404 631898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 602000 419004 635498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 602000 422604 603098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 602000 426204 606698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 428227 606660 428293 606661
rect 428227 606596 428228 606660
rect 428292 606596 428293 606660
rect 428227 606595 428293 606596
rect 428230 604978 428290 606595
rect 432804 602000 433404 613898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 602000 437004 617498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 437795 606660 437861 606661
rect 437795 606596 437796 606660
rect 437860 606596 437861 606660
rect 437795 606595 437861 606596
rect 437798 604978 437858 606595
rect 440004 602000 440604 621098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 602000 444204 624698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 602000 451404 631898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 453987 604212 454053 604213
rect 453987 604148 453988 604212
rect 454052 604148 454053 604212
rect 453987 604147 454053 604148
rect 453990 603805 454050 604147
rect 453987 603804 454053 603805
rect 453987 603740 453988 603804
rect 454052 603740 454053 603804
rect 453987 603739 454053 603740
rect 454404 602000 455004 635498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 458771 606660 458837 606661
rect 458771 606596 458772 606660
rect 458836 606596 458837 606660
rect 458771 606595 458837 606596
rect 458774 604978 458834 606595
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 602000 458604 603098
rect 461604 602000 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 602000 469404 613898
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 602000 473004 617498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 602000 476604 621098
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486371 700364 486437 700365
rect 486371 700300 486372 700364
rect 486436 700300 486437 700364
rect 486371 700299 486437 700300
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 602000 480204 624698
rect 486003 603396 486069 603397
rect 486003 603332 486004 603396
rect 486068 603332 486069 603396
rect 486003 603331 486069 603332
rect 482875 602444 482941 602445
rect 482875 602380 482876 602444
rect 482940 602380 482941 602444
rect 482875 602379 482941 602380
rect 162899 601356 162965 601357
rect 162899 601292 162900 601356
rect 162964 601292 162965 601356
rect 162899 601291 162965 601292
rect 200619 601356 200685 601357
rect 200619 601292 200620 601356
rect 200684 601292 200685 601356
rect 200619 601291 200685 601292
rect 200803 601356 200869 601357
rect 200803 601292 200804 601356
rect 200868 601292 200869 601356
rect 200803 601291 200869 601292
rect 258763 601356 258829 601357
rect 258763 601292 258764 601356
rect 258828 601292 258829 601356
rect 258763 601291 258829 601292
rect 260787 601356 260853 601357
rect 260787 601292 260788 601356
rect 260852 601292 260853 601356
rect 260787 601291 260853 601292
rect 270355 601356 270421 601357
rect 270355 601292 270356 601356
rect 270420 601292 270421 601356
rect 270355 601291 270421 601292
rect 270539 601356 270605 601357
rect 270539 601292 270540 601356
rect 270604 601292 270605 601356
rect 270539 601291 270605 601292
rect 301451 601356 301517 601357
rect 301451 601292 301452 601356
rect 301516 601292 301517 601356
rect 301451 601291 301517 601292
rect 405043 601356 405109 601357
rect 405043 601292 405044 601356
rect 405108 601292 405109 601356
rect 405043 601291 405109 601292
rect 409091 601356 409157 601357
rect 409091 601292 409092 601356
rect 409156 601292 409157 601356
rect 409091 601291 409157 601292
rect 476987 601356 477053 601357
rect 476987 601292 476988 601356
rect 477052 601292 477053 601356
rect 476987 601291 477053 601292
rect 135115 601220 135181 601221
rect 135115 601156 135116 601220
rect 135180 601156 135181 601220
rect 135115 601155 135181 601156
rect 153147 601220 153213 601221
rect 153147 601156 153148 601220
rect 153212 601156 153213 601220
rect 153147 601155 153213 601156
rect 124259 601084 124325 601085
rect 124259 601020 124260 601084
rect 124324 601020 124325 601084
rect 124259 601019 124325 601020
rect 124075 600948 124141 600949
rect 124075 600884 124076 600948
rect 124140 600884 124141 600948
rect 124075 600883 124141 600884
rect 124078 600810 124138 600883
rect 124262 600810 124322 601019
rect 135118 600949 135178 601155
rect 153150 600949 153210 601155
rect 135115 600948 135181 600949
rect 135115 600884 135116 600948
rect 135180 600884 135181 600948
rect 135115 600883 135181 600884
rect 153147 600948 153213 600949
rect 153147 600884 153148 600948
rect 153212 600884 153213 600948
rect 153147 600883 153213 600884
rect 124078 600750 124322 600810
rect 89667 600132 89733 600133
rect 89667 600068 89668 600132
rect 89732 600068 89733 600132
rect 89667 600067 89733 600068
rect 162902 599997 162962 601291
rect 167683 601220 167749 601221
rect 167683 601156 167684 601220
rect 167748 601156 167749 601220
rect 167683 601155 167749 601156
rect 172283 601220 172349 601221
rect 172283 601156 172284 601220
rect 172348 601156 172349 601220
rect 172283 601155 172349 601156
rect 167686 600813 167746 601155
rect 172286 600949 172346 601155
rect 172283 600948 172349 600949
rect 172283 600884 172284 600948
rect 172348 600884 172349 600948
rect 172283 600883 172349 600884
rect 195835 600948 195901 600949
rect 195835 600884 195836 600948
rect 195900 600884 195901 600948
rect 195835 600883 195901 600884
rect 167683 600812 167749 600813
rect 167683 600748 167684 600812
rect 167748 600748 167749 600812
rect 167683 600747 167749 600748
rect 167683 600676 167749 600677
rect 167683 600612 167684 600676
rect 167748 600612 167749 600676
rect 167683 600611 167749 600612
rect 172283 600676 172349 600677
rect 172283 600612 172284 600676
rect 172348 600612 172349 600676
rect 172283 600611 172349 600612
rect 167686 600269 167746 600611
rect 172286 600269 172346 600611
rect 195838 600269 195898 600883
rect 200622 600405 200682 601291
rect 200806 600677 200866 601291
rect 215339 601084 215405 601085
rect 215339 601020 215340 601084
rect 215404 601020 215405 601084
rect 215339 601019 215405 601020
rect 234659 601084 234725 601085
rect 234659 601020 234660 601084
rect 234724 601020 234725 601084
rect 234659 601019 234725 601020
rect 253979 601084 254045 601085
rect 253979 601020 253980 601084
rect 254044 601020 254045 601084
rect 253979 601019 254045 601020
rect 202827 600948 202893 600949
rect 202827 600884 202828 600948
rect 202892 600884 202893 600948
rect 202827 600883 202893 600884
rect 215155 600948 215221 600949
rect 215155 600884 215156 600948
rect 215220 600884 215221 600948
rect 215155 600883 215221 600884
rect 202830 600810 202890 600883
rect 202646 600750 202890 600810
rect 215158 600810 215218 600883
rect 215342 600810 215402 601019
rect 234475 600948 234541 600949
rect 234475 600884 234476 600948
rect 234540 600884 234541 600948
rect 234475 600883 234541 600884
rect 215158 600750 215402 600810
rect 234478 600810 234538 600883
rect 234662 600810 234722 601019
rect 253795 600948 253861 600949
rect 253795 600884 253796 600948
rect 253860 600884 253861 600948
rect 253795 600883 253861 600884
rect 234478 600750 234722 600810
rect 253798 600810 253858 600883
rect 253982 600810 254042 601019
rect 253798 600750 254042 600810
rect 200803 600676 200869 600677
rect 200803 600612 200804 600676
rect 200868 600612 200869 600676
rect 200803 600611 200869 600612
rect 200619 600404 200685 600405
rect 200619 600340 200620 600404
rect 200684 600340 200685 600404
rect 200619 600339 200685 600340
rect 202646 600269 202706 600750
rect 258766 600677 258826 601291
rect 260790 601085 260850 601291
rect 270358 601085 270418 601291
rect 260787 601084 260853 601085
rect 260787 601020 260788 601084
rect 260852 601020 260853 601084
rect 260787 601019 260853 601020
rect 270355 601084 270421 601085
rect 270355 601020 270356 601084
rect 270420 601020 270421 601084
rect 270355 601019 270421 601020
rect 270542 600949 270602 601291
rect 270539 600948 270605 600949
rect 270539 600884 270540 600948
rect 270604 600884 270605 600948
rect 270539 600883 270605 600884
rect 258763 600676 258829 600677
rect 258763 600612 258764 600676
rect 258828 600612 258829 600676
rect 258763 600611 258829 600612
rect 301454 600541 301514 601291
rect 301451 600540 301517 600541
rect 301451 600476 301452 600540
rect 301516 600476 301517 600540
rect 301451 600475 301517 600476
rect 167683 600268 167749 600269
rect 167683 600204 167684 600268
rect 167748 600204 167749 600268
rect 167683 600203 167749 600204
rect 172283 600268 172349 600269
rect 172283 600204 172284 600268
rect 172348 600204 172349 600268
rect 172283 600203 172349 600204
rect 195835 600268 195901 600269
rect 195835 600204 195836 600268
rect 195900 600204 195901 600268
rect 195835 600203 195901 600204
rect 202643 600268 202709 600269
rect 202643 600204 202644 600268
rect 202708 600204 202709 600268
rect 202643 600203 202709 600204
rect 405046 599997 405106 601291
rect 409094 600541 409154 601291
rect 476990 600898 477050 601291
rect 409091 600540 409157 600541
rect 409091 600476 409092 600540
rect 409156 600476 409157 600540
rect 409091 600475 409157 600476
rect 482878 599997 482938 602379
rect 162899 599996 162965 599997
rect 162899 599932 162900 599996
rect 162964 599932 162965 599996
rect 162899 599931 162965 599932
rect 405043 599996 405109 599997
rect 405043 599932 405044 599996
rect 405108 599932 405109 599996
rect 405043 599931 405109 599932
rect 482875 599996 482941 599997
rect 482875 599932 482876 599996
rect 482940 599932 482941 599996
rect 482875 599931 482941 599932
rect 82862 595990 83290 596050
rect 82491 595508 82557 595509
rect 82491 595444 82492 595508
rect 82556 595444 82557 595508
rect 82491 595443 82557 595444
rect 82494 595370 82554 595443
rect 82862 595370 82922 595990
rect 82494 595310 82922 595370
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 81387 581364 81453 581365
rect 81387 581300 81388 581364
rect 81452 581300 81453 581364
rect 81387 581299 81453 581300
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 79731 522884 79797 522885
rect 79731 522820 79732 522884
rect 79796 522820 79797 522884
rect 79731 522819 79797 522820
rect 79547 489972 79613 489973
rect 79547 489908 79548 489972
rect 79612 489908 79613 489972
rect 79547 489907 79613 489908
rect 79363 245172 79429 245173
rect 79363 245108 79364 245172
rect 79428 245108 79429 245172
rect 79363 245107 79429 245108
rect 79366 90541 79426 245107
rect 79363 90540 79429 90541
rect 79363 90476 79364 90540
rect 79428 90476 79429 90540
rect 79363 90475 79429 90476
rect 78443 71364 78509 71365
rect 78443 71300 78444 71364
rect 78508 71300 78509 71364
rect 78443 71299 78509 71300
rect 79550 71093 79610 489907
rect 79734 87549 79794 522819
rect 80004 513654 80604 549098
rect 81203 533764 81269 533765
rect 81203 533700 81204 533764
rect 81268 533700 81269 533764
rect 81203 533699 81269 533700
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 81019 256052 81085 256053
rect 81019 255988 81020 256052
rect 81084 255988 81085 256052
rect 81019 255987 81085 255988
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 79731 87548 79797 87549
rect 79731 87484 79732 87548
rect 79796 87484 79797 87548
rect 79731 87483 79797 87484
rect 80004 81654 80604 117098
rect 81022 93125 81082 255987
rect 81019 93124 81085 93125
rect 81019 93060 81020 93124
rect 81084 93060 81085 93124
rect 81019 93059 81085 93060
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 79547 71092 79613 71093
rect 79547 71028 79548 71092
rect 79612 71028 79613 71092
rect 79547 71027 79613 71028
rect 78075 66876 78141 66877
rect 78075 66812 78076 66876
rect 78140 66812 78141 66876
rect 78075 66811 78141 66812
rect 80004 45654 80604 81098
rect 81206 47565 81266 533699
rect 81390 86189 81450 581299
rect 81571 515540 81637 515541
rect 81571 515476 81572 515540
rect 81636 515476 81637 515540
rect 81571 515475 81637 515476
rect 81574 98837 81634 515475
rect 82491 475012 82557 475013
rect 82491 474948 82492 475012
rect 82556 475010 82557 475012
rect 82556 474950 82922 475010
rect 82556 474948 82557 474950
rect 82491 474947 82557 474948
rect 82862 473650 82922 474950
rect 82862 473590 83474 473650
rect 82491 467668 82557 467669
rect 82491 467604 82492 467668
rect 82556 467604 82557 467668
rect 82491 467603 82557 467604
rect 82494 467530 82554 467603
rect 82494 467470 83290 467530
rect 81755 373012 81821 373013
rect 81755 372948 81756 373012
rect 81820 372948 81821 373012
rect 81755 372947 81821 372948
rect 81571 98836 81637 98837
rect 81571 98772 81572 98836
rect 81636 98772 81637 98836
rect 81571 98771 81637 98772
rect 81387 86188 81453 86189
rect 81387 86124 81388 86188
rect 81452 86124 81453 86188
rect 81387 86123 81453 86124
rect 81758 59941 81818 372947
rect 82491 284884 82557 284885
rect 82491 284820 82492 284884
rect 82556 284820 82557 284884
rect 82491 284819 82557 284820
rect 82494 284610 82554 284819
rect 82494 284550 82922 284610
rect 82862 102509 82922 284550
rect 82859 102508 82925 102509
rect 82859 102444 82860 102508
rect 82924 102444 82925 102508
rect 82859 102443 82925 102444
rect 83230 98973 83290 467470
rect 83227 98972 83293 98973
rect 83227 98908 83228 98972
rect 83292 98908 83293 98972
rect 83227 98907 83293 98908
rect 83414 86325 83474 473590
rect 144867 102644 144933 102645
rect 144867 102580 144868 102644
rect 144932 102580 144933 102644
rect 144867 102579 144933 102580
rect 144870 102373 144930 102579
rect 144867 102372 144933 102373
rect 144867 102308 144868 102372
rect 144932 102308 144933 102372
rect 144867 102307 144933 102308
rect 83411 86324 83477 86325
rect 83411 86260 83412 86324
rect 83476 86260 83477 86324
rect 83411 86259 83477 86260
rect 83604 85254 84204 102000
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 81755 59940 81821 59941
rect 81755 59876 81756 59940
rect 81820 59876 81821 59940
rect 81755 59875 81821 59876
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 81203 47564 81269 47565
rect 81203 47500 81204 47564
rect 81268 47500 81269 47564
rect 81203 47499 81269 47500
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 77155 5812 77221 5813
rect 77155 5748 77156 5812
rect 77220 5748 77221 5812
rect 77155 5747 77221 5748
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 75131 3772 75197 3773
rect 75131 3708 75132 3772
rect 75196 3708 75197 3772
rect 75131 3707 75197 3708
rect 75683 3772 75749 3773
rect 75683 3708 75684 3772
rect 75748 3708 75749 3772
rect 75683 3707 75749 3708
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 92454 91404 102000
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 96054 95004 102000
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 99654 98604 102000
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 67254 102204 102000
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 74454 109404 102000
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 78054 113004 102000
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 81654 116604 102000
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 85254 120204 102000
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 92454 127404 102000
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 96054 131004 102000
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 99654 134604 102000
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 67254 138204 102000
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 74454 145404 102000
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 78054 149004 102000
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 81654 152604 102000
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 155604 85254 156204 102000
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 153147 5948 153213 5949
rect 153147 5884 153148 5948
rect 153212 5884 153213 5948
rect 153147 5883 153213 5884
rect 153150 5677 153210 5883
rect 153147 5676 153213 5677
rect 153147 5612 153148 5676
rect 153212 5612 153213 5676
rect 153147 5611 153213 5612
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 92454 163404 102000
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 96054 167004 102000
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 169526 4045 169586 101542
rect 170004 99654 170604 102000
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 169523 4044 169589 4045
rect 169523 3980 169524 4044
rect 169588 3980 169589 4044
rect 169523 3979 169589 3980
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 67254 174204 102000
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 74454 181404 102000
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 78054 185004 102000
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 81654 188604 102000
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 85254 192204 102000
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 92454 199404 102000
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 96054 203004 102000
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 99654 206604 102000
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 67254 210204 102000
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 74454 217404 102000
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 211107 5948 211173 5949
rect 211107 5884 211108 5948
rect 211172 5884 211173 5948
rect 211107 5883 211173 5884
rect 211110 5405 211170 5883
rect 211107 5404 211173 5405
rect 211107 5340 211108 5404
rect 211172 5340 211173 5404
rect 211107 5339 211173 5340
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 78054 221004 102000
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 224004 81654 224604 102000
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 222147 6084 222213 6085
rect 222147 6020 222148 6084
rect 222212 6020 222213 6084
rect 222147 6019 222213 6020
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 222150 5541 222210 6019
rect 220404 -2186 221004 5498
rect 222147 5540 222213 5541
rect 222147 5476 222148 5540
rect 222212 5476 222213 5540
rect 222147 5475 222213 5476
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 85254 228204 102000
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 92454 235404 102000
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 230427 6084 230493 6085
rect 230427 6020 230428 6084
rect 230492 6020 230493 6084
rect 230427 6019 230493 6020
rect 230430 5541 230490 6019
rect 230427 5540 230493 5541
rect 230427 5476 230428 5540
rect 230492 5476 230493 5540
rect 230427 5475 230493 5476
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 96054 239004 102000
rect 241286 100333 241346 100862
rect 241283 100332 241349 100333
rect 241283 100268 241284 100332
rect 241348 100268 241349 100332
rect 241283 100267 241349 100268
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 242004 99654 242604 102000
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 239995 6084 240061 6085
rect 239995 6020 239996 6084
rect 240060 6020 240061 6084
rect 239995 6019 240061 6020
rect 239998 5813 240058 6019
rect 239995 5812 240061 5813
rect 239995 5748 239996 5812
rect 240060 5748 240061 5812
rect 239995 5747 240061 5748
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 67254 246204 102000
rect 251035 101692 251101 101693
rect 251035 101628 251036 101692
rect 251100 101628 251101 101692
rect 251035 101627 251101 101628
rect 251038 100418 251098 101627
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 74454 253404 102000
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 249747 6084 249813 6085
rect 249747 6020 249748 6084
rect 249812 6020 249813 6084
rect 249747 6019 249813 6020
rect 249750 5813 249810 6019
rect 249747 5812 249813 5813
rect 249747 5748 249748 5812
rect 249812 5748 249813 5812
rect 249747 5747 249813 5748
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 78054 257004 102000
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 81654 260604 102000
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 263604 85254 264204 102000
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 260971 5812 261037 5813
rect 260971 5810 260972 5812
rect 260790 5750 260972 5810
rect 260790 5677 260850 5750
rect 260971 5748 260972 5750
rect 261036 5748 261037 5812
rect 260971 5747 261037 5748
rect 260787 5676 260853 5677
rect 260787 5612 260788 5676
rect 260852 5612 260853 5676
rect 260787 5611 260853 5612
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 92454 271404 102000
rect 273854 100333 273914 100862
rect 273851 100332 273917 100333
rect 273851 100268 273852 100332
rect 273916 100268 273917 100332
rect 273851 100267 273917 100268
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 269067 5812 269133 5813
rect 269067 5748 269068 5812
rect 269132 5748 269133 5812
rect 269067 5747 269133 5748
rect 269070 5541 269130 5747
rect 269067 5540 269133 5541
rect 269067 5476 269068 5540
rect 269132 5476 269133 5540
rect 269067 5475 269133 5476
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 96054 275004 102000
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 99654 278604 102000
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 67254 282204 102000
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 102000
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288387 6084 288453 6085
rect 288387 6020 288388 6084
rect 288452 6020 288453 6084
rect 288387 6019 288453 6020
rect 288390 5813 288450 6019
rect 288387 5812 288453 5813
rect 288387 5748 288388 5812
rect 288452 5748 288453 5812
rect 288387 5747 288453 5748
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 78054 293004 102000
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 81654 296604 102000
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 299604 85254 300204 102000
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 297955 6084 298021 6085
rect 297955 6020 297956 6084
rect 298020 6020 298021 6084
rect 297955 6019 298021 6020
rect 297958 5813 298018 6019
rect 297955 5812 298021 5813
rect 297955 5748 297956 5812
rect 298020 5748 298021 5812
rect 297955 5747 298021 5748
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 92454 307404 102000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 310404 96054 311004 102000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 307707 5812 307773 5813
rect 307707 5748 307708 5812
rect 307772 5748 307773 5812
rect 307707 5747 307773 5748
rect 307710 5541 307770 5747
rect 307707 5540 307773 5541
rect 307707 5476 307708 5540
rect 307772 5476 307773 5540
rect 307707 5475 307773 5476
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 99654 314604 102000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 317604 67254 318204 102000
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 317275 5812 317341 5813
rect 317275 5748 317276 5812
rect 317340 5748 317341 5812
rect 317275 5747 317341 5748
rect 317278 5541 317338 5747
rect 317275 5540 317341 5541
rect 317275 5476 317276 5540
rect 317340 5476 317341 5540
rect 317275 5475 317341 5476
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 74454 325404 102000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 78054 329004 102000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 81654 332604 102000
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 85254 336204 102000
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 92454 343404 102000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 96054 347004 102000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 99654 350604 102000
rect 351134 100333 351194 100862
rect 351131 100332 351197 100333
rect 351131 100268 351132 100332
rect 351196 100268 351197 100332
rect 351131 100267 351197 100268
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 67254 354204 102000
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 74454 361404 102000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360147 5812 360213 5813
rect 360147 5748 360148 5812
rect 360212 5810 360213 5812
rect 360331 5812 360397 5813
rect 360331 5810 360332 5812
rect 360212 5750 360332 5810
rect 360212 5748 360213 5750
rect 360147 5747 360213 5748
rect 360331 5748 360332 5750
rect 360396 5748 360397 5812
rect 360331 5747 360397 5748
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 78054 365004 102000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 368004 81654 368604 102000
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 365667 5812 365733 5813
rect 365667 5748 365668 5812
rect 365732 5748 365733 5812
rect 365667 5747 365733 5748
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 365670 5541 365730 5747
rect 364404 -2186 365004 5498
rect 365667 5540 365733 5541
rect 365667 5476 365668 5540
rect 365732 5476 365733 5540
rect 365667 5475 365733 5476
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 85254 372204 102000
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 92454 379404 102000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 96054 383004 102000
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 386004 99654 386604 102000
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 384987 6084 385053 6085
rect 384987 6020 384988 6084
rect 385052 6020 385053 6084
rect 384987 6019 385053 6020
rect 384990 5813 385050 6019
rect 384987 5812 385053 5813
rect 384987 5748 384988 5812
rect 385052 5748 385053 5812
rect 384987 5747 385053 5748
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 67254 390204 102000
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 74454 397404 102000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 78054 401004 102000
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 81654 404604 102000
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 407604 85254 408204 102000
rect 412406 101013 412466 101542
rect 412403 101012 412469 101013
rect 412403 100948 412404 101012
rect 412468 100948 412469 101012
rect 412403 100947 412469 100948
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 405779 6084 405845 6085
rect 405779 6020 405780 6084
rect 405844 6020 405845 6084
rect 405779 6019 405845 6020
rect 405782 5677 405842 6019
rect 405779 5676 405845 5677
rect 405779 5612 405780 5676
rect 405844 5612 405845 5676
rect 405779 5611 405845 5612
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 92454 415404 102000
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 96054 419004 102000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 99654 422604 102000
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 67254 426204 102000
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 74454 433404 102000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 78054 437004 102000
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 81654 440604 102000
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 85254 444204 102000
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 92454 451404 102000
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 96054 455004 102000
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 458004 99654 458604 102000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 456747 5812 456813 5813
rect 456747 5748 456748 5812
rect 456812 5810 456813 5812
rect 456931 5812 456997 5813
rect 456931 5810 456932 5812
rect 456812 5750 456932 5810
rect 456812 5748 456813 5750
rect 456747 5747 456813 5748
rect 456931 5748 456932 5750
rect 456996 5748 456997 5812
rect 456931 5747 456997 5748
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 67254 462204 102000
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 74454 469404 102000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 466134 2821 466194 3622
rect 466131 2820 466197 2821
rect 466131 2756 466132 2820
rect 466196 2756 466197 2820
rect 466131 2755 466197 2756
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 78054 473004 102000
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 81654 476604 102000
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 85254 480204 102000
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486006 3773 486066 603331
rect 486187 601356 486253 601357
rect 486187 601292 486188 601356
rect 486252 601292 486253 601356
rect 486187 601291 486253 601292
rect 486190 50421 486250 601291
rect 486374 100741 486434 700299
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 602000 487404 631898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 489867 607612 489933 607613
rect 489867 607548 489868 607612
rect 489932 607548 489933 607612
rect 489867 607547 489933 607548
rect 487843 607476 487909 607477
rect 487843 607412 487844 607476
rect 487908 607412 487909 607476
rect 487843 607411 487909 607412
rect 487846 600133 487906 607411
rect 488579 604012 488580 604062
rect 488644 604012 488645 604062
rect 488579 604011 488645 604012
rect 488579 602172 488645 602173
rect 488579 602108 488580 602172
rect 488644 602108 488645 602172
rect 488579 602107 488645 602108
rect 487843 600132 487909 600133
rect 487843 600068 487844 600132
rect 487908 600068 487909 600132
rect 487843 600067 487909 600068
rect 488211 600132 488277 600133
rect 488211 600068 488212 600132
rect 488276 600068 488277 600132
rect 488211 600067 488277 600068
rect 488214 596050 488274 600067
rect 487846 595990 488274 596050
rect 487846 547770 487906 595990
rect 487478 547710 487906 547770
rect 487478 538250 487538 547710
rect 487478 538190 487906 538250
rect 487846 451210 487906 538190
rect 487478 451150 487906 451210
rect 487478 441690 487538 451150
rect 487478 441630 487906 441690
rect 487846 404290 487906 441630
rect 487846 404230 488274 404290
rect 488214 401570 488274 404230
rect 488030 401510 488274 401570
rect 488030 395450 488090 401510
rect 487846 395390 488090 395450
rect 487294 365530 487354 374902
rect 487846 374370 487906 395390
rect 488582 375730 488642 602107
rect 489870 601490 489930 607547
rect 490404 602000 491004 635498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 491155 607340 491221 607341
rect 491155 607276 491156 607340
rect 491220 607276 491221 607340
rect 491155 607275 491221 607276
rect 489686 601430 489930 601490
rect 489686 591970 489746 601430
rect 491158 600130 491218 607275
rect 492811 605028 492877 605029
rect 492811 604964 492812 605028
rect 492876 604964 492877 605028
rect 492811 604963 492877 604964
rect 491891 604892 491957 604893
rect 491891 604828 491892 604892
rect 491956 604828 491957 604892
rect 491891 604827 491957 604828
rect 491158 600070 491586 600130
rect 489867 599996 489933 599997
rect 489867 599932 489868 599996
rect 489932 599932 489933 599996
rect 489867 599931 489933 599932
rect 491155 599996 491221 599997
rect 491155 599932 491156 599996
rect 491220 599932 491221 599996
rect 491155 599931 491221 599932
rect 489318 591910 489746 591970
rect 489318 581770 489378 591910
rect 489318 581710 489562 581770
rect 489502 402250 489562 581710
rect 489870 404290 489930 599931
rect 491158 598178 491218 599931
rect 491526 594690 491586 600070
rect 491526 594630 491770 594690
rect 491710 583810 491770 594630
rect 491526 583750 491770 583810
rect 491526 547770 491586 583750
rect 491526 547710 491770 547770
rect 491710 542330 491770 547710
rect 491342 542270 491770 542330
rect 491342 532810 491402 542270
rect 491342 532750 491770 532810
rect 491710 511730 491770 532750
rect 491342 511670 491770 511730
rect 491342 508330 491402 511670
rect 491894 510370 491954 604827
rect 492627 602308 492693 602309
rect 492627 602244 492628 602308
rect 492692 602244 492693 602308
rect 492627 602243 492693 602244
rect 491526 510310 491954 510370
rect 491526 509010 491586 510310
rect 491526 508950 491954 509010
rect 491342 508270 491770 508330
rect 491710 485890 491770 508270
rect 491526 485830 491770 485890
rect 491526 479770 491586 485830
rect 490974 479710 491586 479770
rect 490974 475690 491034 479710
rect 490974 475630 491770 475690
rect 491710 447130 491770 475630
rect 491526 447070 491770 447130
rect 491526 433530 491586 447070
rect 491894 436250 491954 508950
rect 491894 436190 492322 436250
rect 492262 434890 492322 436190
rect 491894 434830 492322 434890
rect 491526 433470 491770 433530
rect 491710 405650 491770 433470
rect 491342 405590 491770 405650
rect 491342 404378 491402 405590
rect 489870 404230 490114 404290
rect 489134 402190 489562 402250
rect 489134 390010 489194 402190
rect 490054 400210 490114 404230
rect 489870 400150 490114 400210
rect 489134 389950 489746 390010
rect 489686 384570 489746 389950
rect 487662 374310 487906 374370
rect 488398 375670 488642 375730
rect 488766 384510 489746 384570
rect 487662 366210 487722 374310
rect 488398 373690 488458 375670
rect 488766 375138 488826 384510
rect 488398 373630 489010 373690
rect 488950 368250 489010 373630
rect 488582 368190 489010 368250
rect 487662 366150 487906 366210
rect 487294 365470 487538 365530
rect 487478 360090 487538 365470
rect 487478 360030 487722 360090
rect 487662 356010 487722 360030
rect 487478 355950 487722 356010
rect 487478 348530 487538 355950
rect 487294 348470 487538 348530
rect 487294 341730 487354 348470
rect 487294 341670 487722 341730
rect 487662 336970 487722 341670
rect 487478 336910 487722 336970
rect 487478 331530 487538 336910
rect 487478 331470 487722 331530
rect 487662 324050 487722 331470
rect 487846 324730 487906 366150
rect 487846 324670 488274 324730
rect 487662 323990 488090 324050
rect 488030 318610 488090 323990
rect 487662 318550 488090 318610
rect 487662 305690 487722 318550
rect 488214 317930 488274 324670
rect 487846 317870 488274 317930
rect 487846 309090 487906 317870
rect 487846 309030 488274 309090
rect 487478 305630 487722 305690
rect 487478 298210 487538 305630
rect 488214 299570 488274 309030
rect 487294 298150 487538 298210
rect 487846 299510 488274 299570
rect 486742 206498 486802 208302
rect 487294 205730 487354 298150
rect 487846 260810 487906 299510
rect 487662 260750 487906 260810
rect 487662 251290 487722 260750
rect 487662 251230 487906 251290
rect 487294 205670 487722 205730
rect 487662 196210 487722 205670
rect 487110 196150 487722 196210
rect 487110 185330 487170 196150
rect 487110 185270 487354 185330
rect 487294 181930 487354 185270
rect 487294 181870 487722 181930
rect 487662 171050 487722 181870
rect 487478 170990 487722 171050
rect 487478 157450 487538 170990
rect 487294 157390 487538 157450
rect 487294 154050 487354 157390
rect 486926 153990 487354 154050
rect 486926 145298 486986 153990
rect 486926 135690 486986 144382
rect 486926 135630 487722 135690
rect 487662 124130 487722 135630
rect 487478 124070 487722 124130
rect 487478 114610 487538 124070
rect 487110 114550 487538 114610
rect 487110 102237 487170 114550
rect 487107 102236 487173 102237
rect 487107 102172 487108 102236
rect 487172 102172 487173 102236
rect 487107 102171 487173 102172
rect 486371 100740 486437 100741
rect 486371 100676 486372 100740
rect 486436 100676 486437 100740
rect 486371 100675 486437 100676
rect 486804 92454 487404 102000
rect 487846 96661 487906 251230
rect 488214 188138 488274 232102
rect 488582 195530 488642 368190
rect 488582 195470 489010 195530
rect 488950 194170 489010 195470
rect 488582 194110 489010 194170
rect 487843 96660 487909 96661
rect 487843 96596 487844 96660
rect 487908 96596 487909 96660
rect 487843 96595 487909 96596
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486187 50420 486253 50421
rect 486187 50356 486188 50420
rect 486252 50356 486253 50420
rect 486187 50355 486253 50356
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486003 3772 486069 3773
rect 486003 3708 486004 3772
rect 486068 3708 486069 3772
rect 486003 3707 486069 3708
rect 486804 -1266 487404 19898
rect 488582 4045 488642 194110
rect 489134 101829 489194 378302
rect 489131 101828 489197 101829
rect 489131 101764 489132 101828
rect 489196 101764 489197 101828
rect 489131 101763 489197 101764
rect 489870 96661 489930 400150
rect 491894 390010 491954 434830
rect 490974 389950 491954 390010
rect 490974 386698 491034 389950
rect 492262 387290 492322 404142
rect 491526 387230 492322 387290
rect 491526 382530 491586 387230
rect 491158 382470 491586 382530
rect 491158 381850 491218 382470
rect 490974 381790 491218 381850
rect 490974 370970 491034 381790
rect 490974 370910 491218 370970
rect 491158 370290 491218 370910
rect 491158 370230 491586 370290
rect 491526 364850 491586 370230
rect 491526 364790 491770 364850
rect 491710 314530 491770 364790
rect 491526 314470 491770 314530
rect 491526 295490 491586 314470
rect 491526 295430 491770 295490
rect 491710 264890 491770 295430
rect 491526 264830 491770 264890
rect 491526 254010 491586 264830
rect 491342 253950 491586 254010
rect 491342 251290 491402 253950
rect 491342 251230 491586 251290
rect 489867 96660 489933 96661
rect 489867 96596 489868 96660
rect 489932 96596 489933 96660
rect 489867 96595 489933 96596
rect 488579 4044 488645 4045
rect 488579 3980 488580 4044
rect 488644 3980 488645 4044
rect 488579 3979 488645 3980
rect 490238 3909 490298 240942
rect 491526 232338 491586 251230
rect 491894 188138 491954 386462
rect 492262 205818 492322 208302
rect 490404 96054 491004 102000
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490235 3908 490301 3909
rect 490235 3844 490236 3908
rect 490300 3844 490301 3908
rect 490235 3843 490301 3844
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 -3106 491004 23498
rect 491342 9349 491402 187222
rect 491339 9348 491405 9349
rect 491339 9284 491340 9348
rect 491404 9284 491405 9348
rect 491339 9283 491405 9284
rect 491894 3637 491954 183822
rect 492630 6493 492690 602243
rect 492814 102509 492874 604963
rect 494004 603654 494604 639098
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 496859 604756 496925 604757
rect 496859 604692 496860 604756
rect 496924 604692 496925 604756
rect 496859 604691 496925 604692
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 602000 494604 603098
rect 495939 603124 496005 603125
rect 495939 603060 495940 603124
rect 496004 603060 496005 603124
rect 495939 603059 496005 603060
rect 494835 601356 494901 601357
rect 494835 601292 494836 601356
rect 494900 601292 494901 601356
rect 494835 601291 494901 601292
rect 494283 600540 494349 600541
rect 494283 600476 494284 600540
rect 494348 600476 494349 600540
rect 494283 600475 494349 600476
rect 493179 599996 493245 599997
rect 493179 599932 493180 599996
rect 493244 599932 493245 599996
rect 493179 599931 493245 599932
rect 493182 598858 493242 599931
rect 494286 594690 494346 600475
rect 494286 594630 494530 594690
rect 494470 589250 494530 594630
rect 494286 589190 494530 589250
rect 494286 585170 494346 589190
rect 494286 585110 494530 585170
rect 494470 582450 494530 585110
rect 494102 582390 494530 582450
rect 494102 568170 494162 582390
rect 493918 568110 494162 568170
rect 493918 564090 493978 568110
rect 493918 564030 494162 564090
rect 494102 563410 494162 564030
rect 494102 563350 494530 563410
rect 494470 553210 494530 563350
rect 494286 553150 494530 553210
rect 494286 521250 494346 553150
rect 494102 521190 494346 521250
rect 494102 504930 494162 521190
rect 493918 504870 494162 504930
rect 493918 480450 493978 504870
rect 493918 480390 494162 480450
rect 493550 469570 493610 476222
rect 494102 475690 494162 480390
rect 494470 476458 494530 507502
rect 494102 475630 494530 475690
rect 494470 473650 494530 475630
rect 494286 473590 494530 473650
rect 494286 470930 494346 473590
rect 494286 470870 494714 470930
rect 493550 469510 494530 469570
rect 494470 455970 494530 469510
rect 494102 455910 494530 455970
rect 494102 451298 494162 455910
rect 494654 455290 494714 470870
rect 494470 455230 494714 455290
rect 494470 450530 494530 455230
rect 494102 450470 494530 450530
rect 494102 449850 494162 450470
rect 494102 449790 494714 449850
rect 493550 448430 494014 448490
rect 493550 440330 493610 448430
rect 494654 447810 494714 449790
rect 494102 447750 494714 447810
rect 494102 445090 494162 447750
rect 494838 445770 494898 601291
rect 495387 600676 495453 600677
rect 495387 600612 495388 600676
rect 495452 600612 495453 600676
rect 495387 600611 495453 600612
rect 495390 598770 495450 600611
rect 495206 598710 495450 598770
rect 495206 589386 495266 598710
rect 495942 592650 496002 603059
rect 496862 602989 496922 604691
rect 496859 602988 496925 602989
rect 496859 602924 496860 602988
rect 496924 602924 496925 602988
rect 496859 602923 496925 602924
rect 497227 602852 497293 602853
rect 497227 602788 497228 602852
rect 497292 602788 497293 602852
rect 497227 602787 497293 602788
rect 497230 594010 497290 602787
rect 497604 602000 498204 606698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 500907 606524 500973 606525
rect 500907 606460 500908 606524
rect 500972 606460 500973 606524
rect 500907 606459 500973 606460
rect 499435 606116 499501 606117
rect 499435 606052 499436 606116
rect 499500 606052 499501 606116
rect 499435 606051 499501 606052
rect 497595 600948 497661 600949
rect 497595 600884 497596 600948
rect 497660 600884 497661 600948
rect 497595 600883 497661 600884
rect 496862 593950 497290 594010
rect 495942 592590 496370 592650
rect 496310 589386 496370 592590
rect 495206 589326 495450 589386
rect 495390 587890 495450 589326
rect 495022 587830 495450 587890
rect 495942 589326 496370 589386
rect 495022 578370 495082 587830
rect 495022 578310 495634 578370
rect 495574 570210 495634 578310
rect 495390 570150 495634 570210
rect 495390 549130 495450 570150
rect 495390 549070 495634 549130
rect 495574 539610 495634 549070
rect 495390 539550 495634 539610
rect 495390 452570 495450 539550
rect 495390 452510 495818 452570
rect 493918 445030 494162 445090
rect 494654 445710 494898 445770
rect 493918 441010 493978 445030
rect 494654 443730 494714 445710
rect 494654 443670 494898 443730
rect 493918 440950 494714 441010
rect 493550 440270 494162 440330
rect 494102 429450 494162 440270
rect 494654 435570 494714 440950
rect 493734 429390 494162 429450
rect 494286 435510 494714 435570
rect 493734 417210 493794 429390
rect 494286 428770 494346 435510
rect 494102 428710 494346 428770
rect 494838 428770 494898 443670
rect 495758 443050 495818 452510
rect 495390 442990 495818 443050
rect 494838 428710 495266 428770
rect 494102 425370 494162 428710
rect 494102 425310 494714 425370
rect 493734 417150 494346 417210
rect 494286 407010 494346 417150
rect 494654 411090 494714 425310
rect 495206 419930 495266 428710
rect 495390 424010 495450 442990
rect 495390 423950 495818 424010
rect 493550 406950 494346 407010
rect 494470 411030 494714 411090
rect 494838 419870 495266 419930
rect 493182 394858 493242 404142
rect 493550 396898 493610 406950
rect 494470 402250 494530 411030
rect 494286 402190 494530 402250
rect 494286 397490 494346 402190
rect 493918 397430 494346 397490
rect 493918 392730 493978 397430
rect 493918 392670 494346 392730
rect 494286 385930 494346 392670
rect 494102 385870 494346 385930
rect 494102 373690 494162 385870
rect 494470 375730 494530 396662
rect 494286 375670 494530 375730
rect 494286 374370 494346 375670
rect 494286 374310 494530 374370
rect 494102 373630 494346 373690
rect 494286 365530 494346 373630
rect 493734 365470 494346 365530
rect 493734 360178 493794 365470
rect 494470 362130 494530 374310
rect 494102 362070 494530 362130
rect 494102 353290 494162 362070
rect 494102 353230 494346 353290
rect 493918 339690 493978 342262
rect 494286 340370 494346 353230
rect 494470 352610 494530 359942
rect 494838 358138 494898 419870
rect 495758 415442 495818 423950
rect 495390 415382 495818 415442
rect 495390 413810 495450 415382
rect 495206 413750 495450 413810
rect 495206 404378 495266 413750
rect 495390 362130 495450 394622
rect 495206 362070 495450 362130
rect 495206 354650 495266 362070
rect 495206 354590 495450 354650
rect 494470 352550 494714 352610
rect 494654 342498 494714 352550
rect 495390 347170 495450 354590
rect 495022 347110 495450 347170
rect 495022 343178 495082 347110
rect 495574 343090 495634 357902
rect 495390 343030 495634 343090
rect 494286 340310 494898 340370
rect 493918 339630 494714 339690
rect 494654 334930 494714 339630
rect 494838 335610 494898 340310
rect 494838 335550 495266 335610
rect 493918 334870 494714 334930
rect 493918 333570 493978 334870
rect 495206 333570 495266 335550
rect 493918 333510 494162 333570
rect 494102 326090 494162 333510
rect 493734 326030 494162 326090
rect 494286 333510 495266 333570
rect 493366 318610 493426 321862
rect 493734 319970 493794 326030
rect 494286 322098 494346 333510
rect 495390 328130 495450 343030
rect 495942 335018 496002 589326
rect 496862 585170 496922 593950
rect 497598 585170 497658 600883
rect 498331 600812 498397 600813
rect 498331 600748 498332 600812
rect 498396 600748 498397 600812
rect 498331 600747 498397 600748
rect 496862 585110 497106 585170
rect 497046 577098 497106 585110
rect 497230 585110 497658 585170
rect 497230 579594 497290 585110
rect 497230 579534 497658 579594
rect 497598 572930 497658 579534
rect 497598 572870 498210 572930
rect 498150 566130 498210 572870
rect 497966 566070 498210 566130
rect 497966 564770 498026 566070
rect 497230 564710 498026 564770
rect 496862 548450 496922 564622
rect 496678 548390 496922 548450
rect 496678 543690 496738 548390
rect 497230 543690 497290 564710
rect 496678 543630 497106 543690
rect 497230 543630 497658 543690
rect 497046 542330 497106 543630
rect 496678 542270 497106 542330
rect 497598 542330 497658 543630
rect 497598 542270 498026 542330
rect 496678 533490 496738 542270
rect 497966 533490 498026 542270
rect 496678 533430 497106 533490
rect 497046 530090 497106 533430
rect 496678 530030 497106 530090
rect 497598 533430 498026 533490
rect 496678 523290 496738 530030
rect 496678 523230 497106 523290
rect 497046 515130 497106 523230
rect 496862 515070 497106 515130
rect 496862 453338 496922 515070
rect 497598 513090 497658 533430
rect 497230 513030 497658 513090
rect 497230 494050 497290 513030
rect 497046 493990 497290 494050
rect 497046 483170 497106 493990
rect 497046 483110 497290 483170
rect 497230 478410 497290 483110
rect 497230 478350 497658 478410
rect 497598 475010 497658 478350
rect 497598 474950 498210 475010
rect 497598 464750 498026 464810
rect 497598 452570 497658 464750
rect 497966 464130 498026 464750
rect 498150 464130 498210 474950
rect 497966 464070 498210 464130
rect 498334 458282 498394 600747
rect 498702 564858 498762 576862
rect 498334 458222 499314 458282
rect 499254 453250 499314 458222
rect 498334 453190 499314 453250
rect 497414 452510 497658 452570
rect 497414 450530 497474 452510
rect 497966 450530 498026 453102
rect 497414 450470 497658 450530
rect 497598 448490 497658 450470
rect 497414 448430 497658 448490
rect 497782 450470 498026 450530
rect 497414 447810 497474 448430
rect 497230 447750 497474 447810
rect 497230 436930 497290 447750
rect 497782 443730 497842 450470
rect 497782 443670 498026 443730
rect 497230 436870 497474 436930
rect 497046 415170 497106 432702
rect 497414 430130 497474 436870
rect 497966 432938 498026 443670
rect 497230 430070 497474 430130
rect 497230 421970 497290 430070
rect 497230 421910 497474 421970
rect 497414 421290 497474 421910
rect 497414 421230 497842 421290
rect 496862 415110 497106 415170
rect 496862 404290 496922 415110
rect 496126 404230 496922 404290
rect 496126 402930 496186 404230
rect 497782 403698 497842 421230
rect 496126 402870 496370 402930
rect 496310 394090 496370 402870
rect 496310 394030 496738 394090
rect 496678 387970 496738 394030
rect 497414 392050 497474 402782
rect 497230 391990 497474 392050
rect 497230 390098 497290 391990
rect 496678 387910 497106 387970
rect 497046 383210 497106 387910
rect 496862 383150 497106 383210
rect 496862 377090 496922 383150
rect 497230 378538 497290 381022
rect 496862 377030 497106 377090
rect 497046 358050 497106 377030
rect 497046 357990 497658 358050
rect 497598 348530 497658 357990
rect 497046 348470 497658 348530
rect 496310 334250 496370 342942
rect 496126 334190 496370 334250
rect 496126 333570 496186 334190
rect 496678 333570 496738 334782
rect 495206 328070 495450 328130
rect 495574 333510 496186 333570
rect 496310 333510 496738 333570
rect 495206 327450 495266 328070
rect 495574 327450 495634 333510
rect 494838 327390 495266 327450
rect 495390 327390 495634 327450
rect 493734 319910 494714 319970
rect 493366 318550 494530 318610
rect 494470 309090 494530 318550
rect 494102 309030 494530 309090
rect 494102 299658 494162 309030
rect 494654 295490 494714 319910
rect 494838 304330 494898 327390
rect 494838 304270 495082 304330
rect 495022 302290 495082 304270
rect 494286 295430 494714 295490
rect 494838 302230 495082 302290
rect 494286 284610 494346 295430
rect 494838 286650 494898 302230
rect 495390 300250 495450 327390
rect 496310 324730 496370 333510
rect 497046 329490 497106 348470
rect 495942 324670 496370 324730
rect 496862 329430 497106 329490
rect 495390 300190 495818 300250
rect 493734 284550 494346 284610
rect 494654 286590 494898 286650
rect 493734 266338 493794 284550
rect 494654 281978 494714 286590
rect 495206 281890 495266 299422
rect 495758 290730 495818 300190
rect 495022 281830 495266 281890
rect 495390 290670 495818 290730
rect 495022 281210 495082 281830
rect 494286 281150 495082 281210
rect 494286 275090 494346 281150
rect 495022 277130 495082 280382
rect 494838 277070 495082 277130
rect 494286 275030 494530 275090
rect 494470 270330 494530 275030
rect 494286 270270 494530 270330
rect 494286 265570 494346 270270
rect 494838 267018 494898 277070
rect 493918 265510 494346 265570
rect 494838 265570 494898 266102
rect 494838 265510 495266 265570
rect 493918 263530 493978 265510
rect 493918 263470 494346 263530
rect 494286 259538 494346 263470
rect 494838 258770 494898 264062
rect 494286 258710 494898 258770
rect 493366 247890 493426 253182
rect 493918 248570 493978 252502
rect 494286 251970 494346 258710
rect 495206 253330 495266 265510
rect 494838 253270 495266 253330
rect 494838 252738 494898 253270
rect 494286 251910 494898 251970
rect 493918 248510 494714 248570
rect 493366 247830 494530 247890
rect 494470 242450 494530 247830
rect 493550 242390 494530 242450
rect 493550 237778 493610 242390
rect 494654 241090 494714 248510
rect 493918 241030 494714 241090
rect 493918 236330 493978 241030
rect 493918 236270 494162 236330
rect 494102 229530 494162 236270
rect 494102 229470 494346 229530
rect 494286 226130 494346 229470
rect 494102 226070 494346 226130
rect 493734 213210 493794 217142
rect 494102 214570 494162 226070
rect 494470 217378 494530 237542
rect 494102 214510 494714 214570
rect 493734 213150 494530 213210
rect 494470 208450 494530 213150
rect 494286 208390 494530 208450
rect 494286 196210 494346 208390
rect 494286 196150 494530 196210
rect 494470 180570 494530 196150
rect 494102 180510 494530 180570
rect 494102 179978 494162 180510
rect 494654 179210 494714 214510
rect 494838 209130 494898 251910
rect 494838 209070 495266 209130
rect 495206 196210 495266 209070
rect 494102 179150 494714 179210
rect 494838 196150 495266 196210
rect 494102 177850 494162 179150
rect 493918 177790 494162 177850
rect 493182 156178 493242 165462
rect 493918 160850 493978 177790
rect 494838 177170 494898 196150
rect 495390 184058 495450 290670
rect 494838 177110 495266 177170
rect 493734 160790 493978 160850
rect 493734 160170 493794 160790
rect 493550 160110 493794 160170
rect 493550 153370 493610 160110
rect 493182 153310 493610 153370
rect 493182 126170 493242 153310
rect 493182 126110 493610 126170
rect 493182 120138 493242 123302
rect 493550 117330 493610 126110
rect 493550 117270 493794 117330
rect 493734 102509 493794 117270
rect 492811 102508 492877 102509
rect 492811 102444 492812 102508
rect 492876 102444 492877 102508
rect 492811 102443 492877 102444
rect 493731 102508 493797 102509
rect 493731 102444 493732 102508
rect 493796 102444 493797 102508
rect 493731 102443 493797 102444
rect 492995 102372 493061 102373
rect 492995 102308 492996 102372
rect 493060 102308 493061 102372
rect 494470 102370 494530 177022
rect 495206 175810 495266 177110
rect 494838 175750 495266 175810
rect 494838 165698 494898 175750
rect 495206 164930 495266 172942
rect 494654 164870 495266 164930
rect 494654 130250 494714 164870
rect 495022 154730 495082 155942
rect 494838 154670 495082 154730
rect 494838 130930 494898 154670
rect 494838 130870 495450 130930
rect 494654 130190 494898 130250
rect 494838 126986 494898 130190
rect 494654 126926 494898 126986
rect 494654 126850 494714 126926
rect 494654 126790 494898 126850
rect 494838 123538 494898 126790
rect 495390 120730 495450 130870
rect 494838 120670 495450 120730
rect 494838 120050 494898 120670
rect 494654 119990 494898 120050
rect 494654 110530 494714 119990
rect 494654 110470 494898 110530
rect 492995 102307 493061 102308
rect 493734 102310 494530 102370
rect 492811 102236 492877 102237
rect 492811 102172 492812 102236
rect 492876 102172 492877 102236
rect 492811 102171 492877 102172
rect 492814 95981 492874 102171
rect 492998 102101 493058 102307
rect 492995 102100 493061 102101
rect 492995 102036 492996 102100
rect 493060 102036 493061 102100
rect 492995 102035 493061 102036
rect 493734 101421 493794 102310
rect 493731 101420 493797 101421
rect 493731 101356 493732 101420
rect 493796 101356 493797 101420
rect 493731 101355 493797 101356
rect 494004 99654 494604 102000
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492811 95980 492877 95981
rect 492811 95916 492812 95980
rect 492876 95916 492877 95980
rect 492811 95915 492877 95916
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 492627 6492 492693 6493
rect 492627 6428 492628 6492
rect 492692 6428 492693 6492
rect 492627 6427 492693 6428
rect 491891 3636 491957 3637
rect 491891 3572 491892 3636
rect 491956 3572 491957 3636
rect 491891 3571 491957 3572
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 -4946 494604 27098
rect 494838 7581 494898 110470
rect 495206 109170 495266 119902
rect 495206 109110 495312 109170
rect 495252 108490 495312 109110
rect 495206 108430 495312 108490
rect 495206 102237 495266 108430
rect 495203 102236 495269 102237
rect 495203 102172 495204 102236
rect 495268 102172 495269 102236
rect 495203 102171 495269 102172
rect 495206 101013 495266 101542
rect 495203 101012 495269 101013
rect 495203 100948 495204 101012
rect 495268 100948 495269 101012
rect 495203 100947 495269 100948
rect 494835 7580 494901 7581
rect 494835 7516 494836 7580
rect 494900 7516 494901 7580
rect 494835 7515 494901 7516
rect 495574 6765 495634 180422
rect 495942 11661 496002 324670
rect 496862 314530 496922 329430
rect 496862 314470 497106 314530
rect 497046 290730 497106 314470
rect 496862 290670 497106 290730
rect 496862 266930 496922 290670
rect 496678 266870 496922 266930
rect 496310 264298 496370 266782
rect 496678 260810 496738 266870
rect 496494 260750 496738 260810
rect 496494 251970 496554 260750
rect 497046 253418 497106 259302
rect 496126 251910 496554 251970
rect 496126 212530 496186 251910
rect 496126 212470 496370 212530
rect 496310 203010 496370 212470
rect 496126 202950 496370 203010
rect 496126 187778 496186 202950
rect 496126 187718 496738 187778
rect 496678 183290 496738 187718
rect 496310 183230 496738 183290
rect 496310 179890 496370 183230
rect 496126 179830 496370 179890
rect 496126 169690 496186 179830
rect 496126 169630 496370 169690
rect 496310 135690 496370 169630
rect 496126 135630 496370 135690
rect 496126 132290 496186 135630
rect 496126 132230 496370 132290
rect 496310 102098 496370 132230
rect 496310 102038 496554 102098
rect 496494 93941 496554 102038
rect 496491 93940 496557 93941
rect 496491 93876 496492 93940
rect 496556 93876 496557 93940
rect 496491 93875 496557 93876
rect 496491 93668 496557 93669
rect 496491 93604 496492 93668
rect 496556 93604 496557 93668
rect 496491 93603 496557 93604
rect 496494 85645 496554 93603
rect 496491 85644 496557 85645
rect 496491 85580 496492 85644
rect 496556 85580 496557 85644
rect 496491 85579 496557 85580
rect 496491 85372 496557 85373
rect 496491 85308 496492 85372
rect 496556 85308 496557 85372
rect 496491 85307 496557 85308
rect 496494 63610 496554 85307
rect 496310 63550 496554 63610
rect 496310 61570 496370 63550
rect 496310 61510 496554 61570
rect 496494 45525 496554 61510
rect 496491 45524 496557 45525
rect 496491 45460 496492 45524
rect 496556 45460 496557 45524
rect 496491 45459 496557 45460
rect 496307 40764 496373 40765
rect 496307 40700 496308 40764
rect 496372 40700 496373 40764
rect 496307 40699 496373 40700
rect 496310 12613 496370 40699
rect 496307 12612 496373 12613
rect 496307 12548 496308 12612
rect 496372 12548 496373 12612
rect 496307 12547 496373 12548
rect 496123 12340 496189 12341
rect 496123 12276 496124 12340
rect 496188 12276 496189 12340
rect 496123 12275 496189 12276
rect 495939 11660 496005 11661
rect 495939 11596 495940 11660
rect 496004 11596 496005 11660
rect 495939 11595 496005 11596
rect 495571 6764 495637 6765
rect 495571 6700 495572 6764
rect 495636 6700 495637 6764
rect 495571 6699 495637 6700
rect 496126 3858 496186 12275
rect 496862 6357 496922 187902
rect 497966 184738 498026 245702
rect 498334 242538 498394 453190
rect 498702 381938 498762 389862
rect 498702 317930 498762 342942
rect 498518 317870 498762 317930
rect 498518 302290 498578 317870
rect 498518 302230 498762 302290
rect 498702 241770 498762 302230
rect 498702 241710 498946 241770
rect 498886 240410 498946 241710
rect 498702 240350 498946 240410
rect 498702 220690 498762 240350
rect 499438 239050 499498 606051
rect 499803 600268 499869 600269
rect 499803 600204 499804 600268
rect 499868 600204 499869 600268
rect 499803 600203 499869 600204
rect 499806 507738 499866 600203
rect 500910 592650 500970 606459
rect 502379 606388 502445 606389
rect 502379 606324 502380 606388
rect 502444 606324 502445 606388
rect 502379 606323 502445 606324
rect 501643 601764 501709 601765
rect 501643 601700 501644 601764
rect 501708 601700 501709 601764
rect 501643 601699 501709 601700
rect 500910 592590 501154 592650
rect 501094 587890 501154 592590
rect 501646 589389 501706 601699
rect 501643 589388 501709 589389
rect 501643 589324 501644 589388
rect 501708 589324 501709 589388
rect 501643 589323 501709 589324
rect 501827 589116 501893 589117
rect 501827 589052 501828 589116
rect 501892 589052 501893 589116
rect 501827 589051 501893 589052
rect 501830 587890 501890 589051
rect 501094 587830 501338 587890
rect 501278 579050 501338 587830
rect 501646 587830 501890 587890
rect 501646 579733 501706 587830
rect 501643 579732 501709 579733
rect 501643 579668 501644 579732
rect 501708 579668 501709 579732
rect 501643 579667 501709 579668
rect 501643 579596 501709 579597
rect 501643 579532 501644 579596
rect 501708 579532 501709 579596
rect 501643 579531 501709 579532
rect 500726 578990 501338 579050
rect 500726 569530 500786 578990
rect 500726 569470 501338 569530
rect 501278 526421 501338 569470
rect 501646 554981 501706 579531
rect 501643 554980 501709 554981
rect 501643 554916 501644 554980
rect 501708 554916 501709 554980
rect 501643 554915 501709 554916
rect 501827 554844 501893 554845
rect 501827 554780 501828 554844
rect 501892 554780 501893 554844
rect 501827 554779 501893 554780
rect 501830 533490 501890 554779
rect 501830 533430 502074 533490
rect 501275 526420 501341 526421
rect 501275 526356 501276 526420
rect 501340 526356 501341 526420
rect 501275 526355 501341 526356
rect 502014 524789 502074 533430
rect 502011 524788 502077 524789
rect 502011 524724 502012 524788
rect 502076 524724 502077 524788
rect 502011 524723 502077 524724
rect 501275 522884 501341 522885
rect 501275 522820 501276 522884
rect 501340 522820 501341 522884
rect 501275 522819 501341 522820
rect 501278 519890 501338 522819
rect 501827 522340 501893 522341
rect 501827 522276 501828 522340
rect 501892 522276 501893 522340
rect 501827 522275 501893 522276
rect 500910 519830 501338 519890
rect 500910 514450 500970 519830
rect 501830 515130 501890 522275
rect 501830 515070 502074 515130
rect 500910 514390 501706 514450
rect 501459 505612 501525 505613
rect 501459 505610 501460 505612
rect 500726 505550 501460 505610
rect 500726 502210 500786 505550
rect 501459 505548 501460 505550
rect 501524 505548 501525 505612
rect 501459 505547 501525 505548
rect 501646 502210 501706 514390
rect 502014 507789 502074 515070
rect 502011 507788 502077 507789
rect 502011 507724 502012 507788
rect 502076 507724 502077 507788
rect 502011 507723 502077 507724
rect 500358 502150 500786 502210
rect 500910 502150 501706 502210
rect 500358 497450 500418 502150
rect 500910 501530 500970 502150
rect 500174 497390 500418 497450
rect 500542 501470 500970 501530
rect 500174 485210 500234 497390
rect 500542 485210 500602 501470
rect 502011 498268 502077 498269
rect 502011 498204 502012 498268
rect 502076 498204 502077 498268
rect 502011 498203 502077 498204
rect 502014 498130 502074 498203
rect 501646 498070 502074 498130
rect 501459 491060 501525 491061
rect 501459 490996 501460 491060
rect 501524 490996 501525 491060
rect 501459 490995 501525 490996
rect 501462 487338 501522 490995
rect 501646 487525 501706 498070
rect 501643 487524 501709 487525
rect 501643 487460 501644 487524
rect 501708 487460 501709 487524
rect 501643 487459 501709 487460
rect 502011 487524 502077 487525
rect 502011 487460 502012 487524
rect 502076 487460 502077 487524
rect 502011 487459 502077 487460
rect 499990 485150 500234 485210
rect 500358 485150 500602 485210
rect 499990 459370 500050 485150
rect 500358 461410 500418 485150
rect 502014 481541 502074 487459
rect 502011 481540 502077 481541
rect 502011 481476 502012 481540
rect 502076 481476 502077 481540
rect 502011 481475 502077 481476
rect 502011 472020 502077 472021
rect 502011 471956 502012 472020
rect 502076 471956 502077 472020
rect 502011 471955 502077 471956
rect 502014 471885 502074 471955
rect 502011 471884 502077 471885
rect 502011 471820 502012 471884
rect 502076 471820 502077 471884
rect 502011 471819 502077 471820
rect 502011 462636 502077 462637
rect 502011 462572 502012 462636
rect 502076 462572 502077 462636
rect 502011 462571 502077 462572
rect 502014 462090 502074 462571
rect 501646 462030 502074 462090
rect 500358 461350 500786 461410
rect 499990 459310 500418 459370
rect 500358 430130 500418 459310
rect 500726 456650 500786 461350
rect 501646 458965 501706 462030
rect 501643 458964 501709 458965
rect 501643 458900 501644 458964
rect 501708 458900 501709 458964
rect 501643 458899 501709 458900
rect 501643 458284 501709 458285
rect 501643 458220 501644 458284
rect 501708 458220 501709 458284
rect 501643 458219 501709 458220
rect 500174 430070 500418 430130
rect 500542 456590 500786 456650
rect 500542 430130 500602 456590
rect 501646 444410 501706 458219
rect 502011 452708 502077 452709
rect 502011 452644 502012 452708
rect 502076 452644 502077 452708
rect 502011 452643 502077 452644
rect 501278 444350 501706 444410
rect 500542 430070 500970 430130
rect 500174 388650 500234 430070
rect 500910 414490 500970 430070
rect 500542 414430 500970 414490
rect 500542 390010 500602 414430
rect 501278 411770 501338 444350
rect 502014 442917 502074 452643
rect 502011 442916 502077 442917
rect 502011 442852 502012 442916
rect 502076 442852 502077 442916
rect 502011 442851 502077 442852
rect 502011 433396 502077 433397
rect 502011 433332 502012 433396
rect 502076 433332 502077 433396
rect 502011 433331 502077 433332
rect 502014 428501 502074 433331
rect 502011 428500 502077 428501
rect 502011 428436 502012 428500
rect 502076 428436 502077 428500
rect 502011 428435 502077 428436
rect 502011 415444 502077 415445
rect 502011 415380 502012 415444
rect 502076 415380 502077 415444
rect 502011 415379 502077 415380
rect 502014 413949 502074 415379
rect 502011 413948 502077 413949
rect 502011 413884 502012 413948
rect 502076 413884 502077 413948
rect 502011 413883 502077 413884
rect 501278 411710 501706 411770
rect 501646 401570 501706 411710
rect 502011 404428 502077 404429
rect 502011 404364 502012 404428
rect 502076 404364 502077 404428
rect 502011 404363 502077 404364
rect 501462 401510 501706 401570
rect 501462 396810 501522 401510
rect 501278 396750 501522 396810
rect 500542 389950 500786 390010
rect 500174 388590 500418 388650
rect 500358 374370 500418 388590
rect 499990 374310 500418 374370
rect 499990 360090 500050 374310
rect 500726 373690 500786 389950
rect 501278 382530 501338 396750
rect 502014 394637 502074 404363
rect 502011 394636 502077 394637
rect 502011 394572 502012 394636
rect 502076 394572 502077 394636
rect 502011 394571 502077 394572
rect 502011 385116 502077 385117
rect 502011 385052 502012 385116
rect 502076 385052 502077 385116
rect 502011 385051 502077 385052
rect 500358 373630 500786 373690
rect 501094 382470 501338 382530
rect 500358 360770 500418 373630
rect 501094 363490 501154 382470
rect 502014 381850 502074 385051
rect 501830 381790 502074 381850
rect 501094 363430 501338 363490
rect 500358 360710 500602 360770
rect 499990 360030 500234 360090
rect 500174 336970 500234 360030
rect 499806 336910 500234 336970
rect 499806 326090 499866 336910
rect 500542 333570 500602 360710
rect 501278 342410 501338 363430
rect 501830 360909 501890 381790
rect 501827 360908 501893 360909
rect 501827 360844 501828 360908
rect 501892 360844 501893 360908
rect 501827 360843 501893 360844
rect 502195 356148 502261 356149
rect 502195 356084 502196 356148
rect 502260 356084 502261 356148
rect 502195 356083 502261 356084
rect 502198 354653 502258 356083
rect 502195 354652 502261 354653
rect 502195 354588 502196 354652
rect 502260 354588 502261 354652
rect 502195 354587 502261 354588
rect 501643 348532 501709 348533
rect 501643 348468 501644 348532
rect 501708 348468 501709 348532
rect 501643 348467 501709 348468
rect 501646 343178 501706 348467
rect 502195 345132 502261 345133
rect 502195 345068 502196 345132
rect 502260 345068 502261 345132
rect 502195 345067 502261 345068
rect 501278 342350 501522 342410
rect 500358 333510 500602 333570
rect 500358 332890 500418 333510
rect 500174 332830 500418 332890
rect 499806 326030 500050 326090
rect 499990 317250 500050 326030
rect 500174 317930 500234 332830
rect 501462 321741 501522 342350
rect 502198 339693 502258 345067
rect 502195 339692 502261 339693
rect 502195 339628 502196 339692
rect 502260 339628 502261 339692
rect 502195 339627 502261 339628
rect 502011 339420 502077 339421
rect 502011 339356 502012 339420
rect 502076 339356 502077 339420
rect 502011 339355 502077 339356
rect 502014 335341 502074 339355
rect 502011 335340 502077 335341
rect 502011 335276 502012 335340
rect 502076 335276 502077 335340
rect 502011 335275 502077 335276
rect 502195 325820 502261 325821
rect 502195 325756 502196 325820
rect 502260 325756 502261 325820
rect 502195 325755 502261 325756
rect 501459 321740 501525 321741
rect 501459 321676 501460 321740
rect 501524 321676 501525 321740
rect 501459 321675 501525 321676
rect 502198 319970 502258 325755
rect 502014 319910 502258 319970
rect 500174 317870 500786 317930
rect 499990 317190 500418 317250
rect 500358 298210 500418 317190
rect 500726 314530 500786 317870
rect 500542 314470 500786 314530
rect 500542 313170 500602 314470
rect 500542 313110 500786 313170
rect 500358 298150 500602 298210
rect 500542 297530 500602 298150
rect 500358 297470 500602 297530
rect 500358 278490 500418 297470
rect 500726 296850 500786 313110
rect 501459 311948 501525 311949
rect 501459 311884 501460 311948
rect 501524 311884 501525 311948
rect 501459 311883 501525 311884
rect 499806 278430 500418 278490
rect 500542 296790 500786 296850
rect 499806 253330 499866 278430
rect 500542 277810 500602 296790
rect 501462 288010 501522 311883
rect 502014 297938 502074 319910
rect 502014 297878 502258 297938
rect 502198 292090 502258 297878
rect 499622 253270 499866 253330
rect 500174 277750 500602 277810
rect 500910 287950 501522 288010
rect 501830 292030 502258 292090
rect 499622 241090 499682 253270
rect 500174 246530 500234 277750
rect 500910 256050 500970 287950
rect 501830 269245 501890 292030
rect 501827 269244 501893 269245
rect 501827 269180 501828 269244
rect 501892 269180 501893 269244
rect 501827 269179 501893 269180
rect 502011 269244 502077 269245
rect 502011 269180 502012 269244
rect 502076 269180 502077 269244
rect 502011 269179 502077 269180
rect 501275 256052 501341 256053
rect 501275 256050 501276 256052
rect 500910 255990 501276 256050
rect 501275 255988 501276 255990
rect 501340 255988 501341 256052
rect 501275 255987 501341 255988
rect 501459 256052 501525 256053
rect 501459 255988 501460 256052
rect 501524 255988 501525 256052
rect 501459 255987 501525 255988
rect 500174 246470 500786 246530
rect 500726 245938 500786 246470
rect 499622 241030 500234 241090
rect 499438 238990 499866 239050
rect 499806 237010 499866 238990
rect 499438 236950 499866 237010
rect 498702 220630 498946 220690
rect 498886 219602 498946 220630
rect 498702 219542 498946 219602
rect 498702 166290 498762 219542
rect 499070 210490 499130 234822
rect 499438 219330 499498 236950
rect 499438 219270 499866 219330
rect 499806 217970 499866 219270
rect 499438 217910 499866 217970
rect 499070 210430 499314 210490
rect 499254 209810 499314 210430
rect 498886 209750 499314 209810
rect 498886 171050 498946 209750
rect 498886 170990 499130 171050
rect 498518 166230 498762 166290
rect 497414 9077 497474 155942
rect 497782 143938 497842 147782
rect 498518 147250 498578 166230
rect 499070 162298 499130 170990
rect 498886 154866 498946 161382
rect 499438 156178 499498 217910
rect 500174 197570 500234 241030
rect 501462 229261 501522 255987
rect 502014 255370 502074 269179
rect 501646 255310 502074 255370
rect 501459 229260 501525 229261
rect 501459 229196 501460 229260
rect 501524 229196 501525 229260
rect 501459 229195 501525 229196
rect 501459 228988 501525 228989
rect 501459 228924 501460 228988
rect 501524 228924 501525 228988
rect 501459 228923 501525 228924
rect 501462 228850 501522 228923
rect 501646 228853 501706 255310
rect 502011 238916 502077 238917
rect 502011 238852 502012 238916
rect 502076 238852 502077 238916
rect 502011 238851 502077 238852
rect 502014 235058 502074 238851
rect 501278 228790 501522 228850
rect 501643 228852 501709 228853
rect 501278 219605 501338 228790
rect 501643 228788 501644 228852
rect 501708 228788 501709 228852
rect 501643 228787 501709 228788
rect 501827 220930 501893 220931
rect 501827 220866 501828 220930
rect 501892 220866 501893 220930
rect 501827 220865 501893 220866
rect 501275 219604 501341 219605
rect 501275 219540 501276 219604
rect 501340 219540 501341 219604
rect 501275 219539 501341 219540
rect 501459 219468 501525 219469
rect 501459 219404 501460 219468
rect 501524 219404 501525 219468
rect 501459 219403 501525 219404
rect 501462 209810 501522 219403
rect 501462 209750 501706 209810
rect 501459 205732 501525 205733
rect 501459 205730 501460 205732
rect 501242 205670 501460 205730
rect 501459 205668 501460 205670
rect 501524 205668 501525 205732
rect 501459 205667 501525 205668
rect 501459 198932 501525 198933
rect 501459 198930 501460 198932
rect 499806 197510 500234 197570
rect 500726 198870 501460 198930
rect 499806 194170 499866 197510
rect 499806 194110 500234 194170
rect 500174 184650 500234 194110
rect 500726 189410 500786 198870
rect 501459 198868 501460 198870
rect 501524 198868 501525 198932
rect 501459 198867 501525 198868
rect 499990 184590 500234 184650
rect 500358 189350 500786 189410
rect 499990 171050 500050 184590
rect 499806 170990 500050 171050
rect 499806 161530 499866 170990
rect 500358 162978 500418 189350
rect 501278 183970 501338 184502
rect 501459 183972 501525 183973
rect 501459 183970 501460 183972
rect 501278 183910 501460 183970
rect 501459 183908 501460 183910
rect 501524 183908 501525 183972
rect 501459 183907 501525 183908
rect 501646 179890 501706 209750
rect 501830 206957 501890 220865
rect 501827 206956 501893 206957
rect 501827 206892 501828 206956
rect 501892 206892 501893 206956
rect 501827 206891 501893 206892
rect 502011 206820 502077 206821
rect 502011 206756 502012 206820
rect 502076 206756 502077 206820
rect 502011 206755 502077 206756
rect 502014 187781 502074 206755
rect 502011 187780 502077 187781
rect 502011 187716 502012 187780
rect 502076 187716 502077 187780
rect 502011 187715 502077 187716
rect 502195 187508 502261 187509
rect 502195 187444 502196 187508
rect 502260 187444 502261 187508
rect 502195 187443 502261 187444
rect 502198 182885 502258 187443
rect 501827 182884 501893 182885
rect 501827 182820 501828 182884
rect 501892 182820 501893 182884
rect 501827 182819 501893 182820
rect 502195 182884 502261 182885
rect 502195 182820 502196 182884
rect 502260 182820 502261 182884
rect 502195 182819 502261 182820
rect 501094 179830 501706 179890
rect 501094 179210 501154 179830
rect 500910 179150 501154 179210
rect 499806 161470 500050 161530
rect 498886 154806 499130 154866
rect 499070 154050 499130 154806
rect 498702 153990 499130 154050
rect 498702 151330 498762 153990
rect 498702 151270 498946 151330
rect 498886 148018 498946 151270
rect 499438 147338 499498 151862
rect 498518 147190 498762 147250
rect 498150 143258 498210 147102
rect 497782 102645 497842 136902
rect 497779 102644 497845 102645
rect 497779 102580 497780 102644
rect 497844 102580 497845 102644
rect 497779 102579 497845 102580
rect 497604 67254 498204 102000
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 498702 67010 498762 147190
rect 499990 145298 500050 161470
rect 500358 146570 500418 161382
rect 500358 146510 500786 146570
rect 499070 144470 499682 144530
rect 499070 143938 499130 144470
rect 499622 143850 499682 144470
rect 499622 143790 500418 143850
rect 499070 142490 499130 143022
rect 499070 142430 499498 142490
rect 499438 129570 499498 142430
rect 499990 137050 500050 142342
rect 499806 136990 500050 137050
rect 499806 134330 499866 136990
rect 500358 134330 500418 143790
rect 499806 134270 500050 134330
rect 499254 129510 499498 129570
rect 499254 128210 499314 129510
rect 499254 128150 499682 128210
rect 499254 115970 499314 126702
rect 499622 124810 499682 128150
rect 498886 115910 499314 115970
rect 499438 124750 499682 124810
rect 498886 100741 498946 115910
rect 498883 100740 498949 100741
rect 498883 100676 498884 100740
rect 498948 100676 498949 100740
rect 498883 100675 498949 100676
rect 499438 86730 499498 124750
rect 499990 120730 500050 134270
rect 500174 134270 500418 134330
rect 500174 130930 500234 134270
rect 500174 130870 500418 130930
rect 500358 126938 500418 130870
rect 500726 124810 500786 146510
rect 500910 127530 500970 179150
rect 501459 154868 501525 154869
rect 501459 154804 501460 154868
rect 501524 154804 501525 154868
rect 501459 154803 501525 154804
rect 501462 152098 501522 154803
rect 501459 151196 501525 151197
rect 501459 151132 501460 151196
rect 501524 151132 501525 151196
rect 501459 151131 501525 151132
rect 500910 127470 501338 127530
rect 501278 126850 501338 127470
rect 501462 126989 501522 151131
rect 501830 145890 501890 182819
rect 501830 145830 502074 145890
rect 501643 137868 501709 137869
rect 501643 137804 501644 137868
rect 501708 137804 501709 137868
rect 501643 137803 501709 137804
rect 501459 126988 501525 126989
rect 501459 126924 501460 126988
rect 501524 126924 501525 126988
rect 501459 126923 501525 126924
rect 501278 126790 501522 126850
rect 500358 124750 500786 124810
rect 500358 122770 500418 124750
rect 500358 122710 500602 122770
rect 499990 120670 500418 120730
rect 500358 115970 500418 120670
rect 500174 115910 500418 115970
rect 499806 97205 499866 115822
rect 500174 112570 500234 115910
rect 500174 112510 500418 112570
rect 500358 111210 500418 112510
rect 499990 111150 500418 111210
rect 499990 102373 500050 111150
rect 499987 102372 500053 102373
rect 499987 102308 499988 102372
rect 500052 102308 500053 102372
rect 499987 102307 500053 102308
rect 500171 102236 500237 102237
rect 500171 102172 500172 102236
rect 500236 102172 500237 102236
rect 500171 102171 500237 102172
rect 499803 97204 499869 97205
rect 499803 97140 499804 97204
rect 499868 97140 499869 97204
rect 499803 97139 499869 97140
rect 500174 87413 500234 102171
rect 500542 87685 500602 122710
rect 501462 121549 501522 126790
rect 501459 121548 501525 121549
rect 501459 121484 501460 121548
rect 501524 121484 501525 121548
rect 501459 121483 501525 121484
rect 501646 121410 501706 137803
rect 502014 137138 502074 145830
rect 502011 122772 502077 122773
rect 502011 122708 502012 122772
rect 502076 122708 502077 122772
rect 502011 122707 502077 122708
rect 501094 121350 501706 121410
rect 501094 120730 501154 121350
rect 501643 121276 501709 121277
rect 501643 121212 501644 121276
rect 501708 121212 501709 121276
rect 501643 121211 501709 121212
rect 500910 120670 501154 120730
rect 500910 102645 500970 120670
rect 501459 119372 501525 119373
rect 501459 119308 501460 119372
rect 501524 119308 501525 119372
rect 501459 119307 501525 119308
rect 500907 102644 500973 102645
rect 500907 102580 500908 102644
rect 500972 102580 500973 102644
rect 500907 102579 500973 102580
rect 501275 102644 501341 102645
rect 501275 102580 501276 102644
rect 501340 102580 501341 102644
rect 501275 102579 501341 102580
rect 501278 92445 501338 102579
rect 501275 92444 501341 92445
rect 501275 92380 501276 92444
rect 501340 92380 501341 92444
rect 501275 92379 501341 92380
rect 501091 92308 501157 92309
rect 501091 92244 501092 92308
rect 501156 92244 501157 92308
rect 501091 92243 501157 92244
rect 500539 87684 500605 87685
rect 500539 87620 500540 87684
rect 500604 87620 500605 87684
rect 500539 87619 500605 87620
rect 500171 87412 500237 87413
rect 500171 87348 500172 87412
rect 500236 87348 500237 87412
rect 500171 87347 500237 87348
rect 500723 87412 500789 87413
rect 500723 87348 500724 87412
rect 500788 87348 500789 87412
rect 500723 87347 500789 87348
rect 499438 86670 499682 86730
rect 499622 77485 499682 86670
rect 499619 77484 499685 77485
rect 499619 77420 499620 77484
rect 499684 77420 499685 77484
rect 499619 77419 499685 77420
rect 499435 77348 499501 77349
rect 499435 77284 499436 77348
rect 499500 77284 499501 77348
rect 499435 77283 499501 77284
rect 499438 75173 499498 77283
rect 499435 75172 499501 75173
rect 499435 75108 499436 75172
rect 499500 75108 499501 75172
rect 499435 75107 499501 75108
rect 499067 67692 499133 67693
rect 499067 67628 499068 67692
rect 499132 67628 499133 67692
rect 500726 67690 500786 87347
rect 499067 67627 499133 67628
rect 500542 67630 500786 67690
rect 499070 67013 499130 67627
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 498518 66950 498762 67010
rect 499067 67012 499133 67013
rect 498518 61570 498578 66950
rect 499067 66948 499068 67012
rect 499132 66948 499133 67012
rect 500542 67010 500602 67630
rect 501094 67010 501154 92243
rect 499067 66947 499133 66948
rect 500358 66950 500602 67010
rect 500910 66950 501154 67010
rect 498518 61510 498762 61570
rect 498702 31650 498762 61510
rect 499251 60076 499317 60077
rect 499251 60012 499252 60076
rect 499316 60012 499317 60076
rect 499251 60011 499317 60012
rect 499254 55181 499314 60011
rect 500358 57221 500418 66950
rect 500910 60893 500970 66950
rect 500907 60892 500973 60893
rect 500907 60828 500908 60892
rect 500972 60828 500973 60892
rect 500907 60827 500973 60828
rect 501091 60620 501157 60621
rect 501091 60556 501092 60620
rect 501156 60556 501157 60620
rect 501091 60555 501157 60556
rect 500355 57220 500421 57221
rect 500355 57156 500356 57220
rect 500420 57156 500421 57220
rect 500355 57155 500421 57156
rect 499251 55180 499317 55181
rect 499251 55116 499252 55180
rect 499316 55116 499317 55180
rect 499251 55115 499317 55116
rect 499251 45796 499317 45797
rect 499251 45732 499252 45796
rect 499316 45732 499317 45796
rect 499251 45731 499317 45732
rect 499254 45525 499314 45731
rect 501094 45525 501154 60555
rect 499251 45524 499317 45525
rect 499251 45460 499252 45524
rect 499316 45460 499317 45524
rect 499251 45459 499317 45460
rect 501091 45524 501157 45525
rect 501091 45460 501092 45524
rect 501156 45460 501157 45524
rect 501091 45459 501157 45460
rect 499251 40764 499317 40765
rect 499251 40700 499252 40764
rect 499316 40700 499317 40764
rect 499251 40699 499317 40700
rect 499254 31650 499314 40699
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 497411 9076 497477 9077
rect 497411 9012 497412 9076
rect 497476 9012 497477 9076
rect 497411 9011 497477 9012
rect 496859 6356 496925 6357
rect 496859 6292 496860 6356
rect 496924 6292 496925 6356
rect 496859 6291 496925 6292
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 498334 31590 498762 31650
rect 499070 31590 499314 31650
rect 498334 28933 498394 31590
rect 498331 28932 498397 28933
rect 498331 28868 498332 28932
rect 498396 28868 498397 28932
rect 498331 28867 498397 28868
rect 499070 22130 499130 31590
rect 498886 22070 499130 22130
rect 498886 21450 498946 22070
rect 498886 21390 499314 21450
rect 498515 21180 498581 21181
rect 498515 21116 498516 21180
rect 498580 21116 498581 21180
rect 498515 21115 498581 21116
rect 498518 19410 498578 21115
rect 498518 19350 498762 19410
rect 498702 14650 498762 19350
rect 498334 14590 498762 14650
rect 498334 11930 498394 14590
rect 498334 11870 498578 11930
rect 498518 8941 498578 11870
rect 498515 8940 498581 8941
rect 498515 8876 498516 8940
rect 498580 8876 498581 8940
rect 498515 8875 498581 8876
rect 499254 4861 499314 21390
rect 499251 4860 499317 4861
rect 499251 4796 499252 4860
rect 499316 4796 499317 4860
rect 499251 4795 499317 4796
rect 501462 3501 501522 119307
rect 501646 71229 501706 121211
rect 502014 116058 502074 122707
rect 502382 102781 502442 606323
rect 504804 578454 505404 613898
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 507899 606252 507965 606253
rect 507899 606188 507900 606252
rect 507964 606188 507965 606252
rect 507899 606187 507965 606188
rect 505507 579188 505573 579189
rect 505507 579124 505508 579188
rect 505572 579124 505573 579188
rect 505507 579123 505573 579124
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504219 531588 504285 531589
rect 504219 531524 504220 531588
rect 504284 531524 504285 531588
rect 504219 531523 504285 531524
rect 502563 517172 502629 517173
rect 502563 517108 502564 517172
rect 502628 517108 502629 517172
rect 502563 517107 502629 517108
rect 502379 102780 502445 102781
rect 502379 102716 502380 102780
rect 502444 102716 502445 102780
rect 502379 102715 502445 102716
rect 501643 71228 501709 71229
rect 501643 71164 501644 71228
rect 501708 71164 501709 71228
rect 501643 71163 501709 71164
rect 502566 50285 502626 517107
rect 502747 509828 502813 509829
rect 502747 509764 502748 509828
rect 502812 509764 502813 509828
rect 502747 509763 502813 509764
rect 502750 51781 502810 509763
rect 504035 297940 504101 297941
rect 504035 297876 504036 297940
rect 504100 297876 504101 297940
rect 504035 297875 504101 297876
rect 504038 283389 504098 297875
rect 504035 283388 504101 283389
rect 504035 283324 504036 283388
rect 504100 283324 504101 283388
rect 504035 283323 504101 283324
rect 504035 280260 504101 280261
rect 504035 280196 504036 280260
rect 504100 280196 504101 280260
rect 504035 280195 504101 280196
rect 504038 254421 504098 280195
rect 504035 254420 504101 254421
rect 504035 254356 504036 254420
rect 504100 254356 504101 254420
rect 504035 254355 504101 254356
rect 503667 253876 503733 253877
rect 503667 253812 503668 253876
rect 503732 253812 503733 253876
rect 503667 253811 503733 253812
rect 503670 232253 503730 253811
rect 503667 232252 503733 232253
rect 503667 232188 503668 232252
rect 503732 232188 503733 232252
rect 503667 232187 503733 232188
rect 503851 231878 503917 231879
rect 503851 231814 503852 231878
rect 503916 231814 503917 231878
rect 503851 231813 503917 231814
rect 503854 194581 503914 231813
rect 503851 194580 503917 194581
rect 503851 194516 503852 194580
rect 503916 194516 503917 194580
rect 503851 194515 503917 194516
rect 504035 192132 504101 192133
rect 504035 192068 504036 192132
rect 504100 192068 504101 192132
rect 504035 192067 504101 192068
rect 503851 185060 503917 185061
rect 503851 184996 503852 185060
rect 503916 184996 503917 185060
rect 503851 184995 503917 184996
rect 503854 175269 503914 184995
rect 503851 175268 503917 175269
rect 503851 175204 503852 175268
rect 503916 175204 503917 175268
rect 503851 175203 503917 175204
rect 503667 174044 503733 174045
rect 503667 173980 503668 174044
rect 503732 173980 503733 174044
rect 503667 173979 503733 173980
rect 503670 173770 503730 173979
rect 503486 173710 503730 173770
rect 503486 173178 503546 173710
rect 503851 165646 503917 165647
rect 503851 165582 503852 165646
rect 503916 165582 503917 165646
rect 503851 165581 503917 165582
rect 503854 164930 503914 165581
rect 503670 164870 503914 164930
rect 503670 145890 503730 164870
rect 503670 145830 503914 145890
rect 503854 126170 503914 145830
rect 503670 126110 503914 126170
rect 503670 87410 503730 126110
rect 503670 87350 503914 87410
rect 503854 79389 503914 87350
rect 503851 79388 503917 79389
rect 503851 79324 503852 79388
rect 503916 79324 503917 79388
rect 503851 79323 503917 79324
rect 502747 51780 502813 51781
rect 502747 51716 502748 51780
rect 502812 51716 502813 51780
rect 502747 51715 502813 51716
rect 502563 50284 502629 50285
rect 502563 50220 502564 50284
rect 502628 50220 502629 50284
rect 502563 50219 502629 50220
rect 504038 26893 504098 192067
rect 504222 186285 504282 531523
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504219 186284 504285 186285
rect 504219 186220 504220 186284
rect 504284 186220 504285 186284
rect 504219 186219 504285 186220
rect 504219 185332 504285 185333
rect 504219 185268 504220 185332
rect 504284 185268 504285 185332
rect 504219 185267 504285 185268
rect 504222 176629 504282 185267
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504219 176628 504285 176629
rect 504219 176564 504220 176628
rect 504284 176564 504285 176628
rect 504219 176563 504285 176564
rect 504219 175404 504285 175405
rect 504219 175340 504220 175404
rect 504284 175340 504285 175404
rect 504219 175339 504285 175340
rect 504222 99109 504282 175339
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504590 101013 504650 101542
rect 504587 101012 504653 101013
rect 504587 100948 504588 101012
rect 504652 100948 504653 101012
rect 504587 100947 504653 100948
rect 504219 99108 504285 99109
rect 504219 99044 504220 99108
rect 504284 99044 504285 99108
rect 504219 99043 504285 99044
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504035 26892 504101 26893
rect 504035 26828 504036 26892
rect 504100 26828 504101 26892
rect 504035 26827 504101 26828
rect 501459 3500 501525 3501
rect 501459 3436 501460 3500
rect 501524 3436 501525 3500
rect 501459 3435 501525 3436
rect 504804 2454 505404 37898
rect 505510 36549 505570 579123
rect 506427 557156 506493 557157
rect 506427 557092 506428 557156
rect 506492 557092 506493 557156
rect 506427 557091 506493 557092
rect 505691 513364 505757 513365
rect 505691 513300 505692 513364
rect 505756 513300 505757 513364
rect 505691 513299 505757 513300
rect 505694 86325 505754 513299
rect 505875 480452 505941 480453
rect 505875 480388 505876 480452
rect 505940 480388 505941 480452
rect 505875 480387 505941 480388
rect 505691 86324 505757 86325
rect 505691 86260 505692 86324
rect 505756 86260 505757 86324
rect 505691 86259 505757 86260
rect 505878 72453 505938 480387
rect 506430 87821 506490 557091
rect 506611 466036 506677 466037
rect 506611 465972 506612 466036
rect 506676 465972 506677 466036
rect 506611 465971 506677 465972
rect 506427 87820 506493 87821
rect 506427 87756 506428 87820
rect 506492 87756 506493 87820
rect 506427 87755 506493 87756
rect 505875 72452 505941 72453
rect 505875 72388 505876 72452
rect 505940 72388 505941 72452
rect 505875 72387 505941 72388
rect 506614 46205 506674 465971
rect 506795 454884 506861 454885
rect 506795 454820 506796 454884
rect 506860 454820 506861 454884
rect 506795 454819 506861 454820
rect 506611 46204 506677 46205
rect 506611 46140 506612 46204
rect 506676 46140 506677 46204
rect 506611 46139 506677 46140
rect 506798 44845 506858 454819
rect 507163 228172 507229 228173
rect 507163 228108 507164 228172
rect 507228 228108 507229 228172
rect 507163 228107 507229 228108
rect 507166 226898 507226 228107
rect 506795 44844 506861 44845
rect 506795 44780 506796 44844
rect 506860 44780 506861 44844
rect 506795 44779 506861 44780
rect 505507 36548 505573 36549
rect 505507 36484 505508 36548
rect 505572 36484 505573 36548
rect 505507 36483 505573 36484
rect 507902 6629 507962 606187
rect 508404 582054 509004 617498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 519491 697236 519557 697237
rect 519491 697172 519492 697236
rect 519556 697172 519557 697236
rect 519491 697171 519557 697172
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 512683 681868 512749 681869
rect 512683 681804 512684 681868
rect 512748 681804 512749 681868
rect 512683 681803 512749 681804
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 509190 90405 509250 600662
rect 511211 600404 511277 600405
rect 511211 600340 511212 600404
rect 511276 600340 511277 600404
rect 511211 600339 511277 600340
rect 510659 502484 510725 502485
rect 510659 502420 510660 502484
rect 510724 502420 510725 502484
rect 510659 502419 510725 502420
rect 509371 418436 509437 418437
rect 509371 418372 509372 418436
rect 509436 418372 509437 418436
rect 509371 418371 509437 418372
rect 509187 90404 509253 90405
rect 509187 90340 509188 90404
rect 509252 90340 509253 90404
rect 509187 90339 509253 90340
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 507899 6628 507965 6629
rect 507899 6564 507900 6628
rect 507964 6564 507965 6628
rect 507899 6563 507965 6564
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 6054 509004 41498
rect 509374 30973 509434 418371
rect 510662 80069 510722 502419
rect 511214 87005 511274 600339
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 511579 227492 511645 227493
rect 511579 227428 511580 227492
rect 511644 227428 511645 227492
rect 511579 227427 511645 227428
rect 511582 226898 511642 227427
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 511211 87004 511277 87005
rect 511211 86940 511212 87004
rect 511276 86940 511277 87004
rect 511211 86939 511277 86940
rect 512004 81654 512604 117098
rect 512686 114613 512746 681803
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 513419 596324 513485 596325
rect 513419 596260 513420 596324
rect 513484 596260 513485 596324
rect 513419 596259 513485 596260
rect 512683 114612 512749 114613
rect 512683 114548 512684 114612
rect 512748 114548 512749 114612
rect 512683 114547 512749 114548
rect 513422 101098 513482 596259
rect 515604 589254 516204 624698
rect 516731 605980 516797 605981
rect 516731 605916 516732 605980
rect 516796 605916 516797 605980
rect 516731 605915 516797 605916
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 510659 80068 510725 80069
rect 510659 80004 510660 80068
rect 510724 80004 510725 80068
rect 510659 80003 510725 80004
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 509371 30972 509437 30973
rect 509371 30908 509372 30972
rect 509436 30908 509437 30972
rect 509371 30907 509437 30908
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 516734 29069 516794 605915
rect 519494 97885 519554 697171
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522070 592109 522130 597942
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522067 592108 522133 592109
rect 522067 592044 522068 592108
rect 522132 592044 522133 592108
rect 522067 592043 522133 592044
rect 521883 591836 521949 591837
rect 521883 591772 521884 591836
rect 521948 591772 521949 591836
rect 521883 591771 521949 591772
rect 521886 582453 521946 591771
rect 521883 582452 521949 582453
rect 521883 582388 521884 582452
rect 521948 582388 521949 582452
rect 521883 582387 521949 582388
rect 522067 582180 522133 582181
rect 522067 582116 522068 582180
rect 522132 582116 522133 582180
rect 522067 582115 522133 582116
rect 522070 579597 522130 582115
rect 522067 579596 522133 579597
rect 522067 579532 522068 579596
rect 522132 579532 522133 579596
rect 522067 579531 522133 579532
rect 521883 570076 521949 570077
rect 521883 570012 521884 570076
rect 521948 570012 521949 570076
rect 521883 570011 521949 570012
rect 521886 563141 521946 570011
rect 521883 563140 521949 563141
rect 521883 563076 521884 563140
rect 521948 563076 521949 563140
rect 521883 563075 521949 563076
rect 522067 562868 522133 562869
rect 522067 562804 522068 562868
rect 522132 562804 522133 562868
rect 522067 562803 522133 562804
rect 522070 560285 522130 562803
rect 522804 560454 523404 595898
rect 522067 560284 522133 560285
rect 522067 560220 522068 560284
rect 522132 560220 522133 560284
rect 522067 560219 522133 560220
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522251 550764 522317 550765
rect 522251 550700 522252 550764
rect 522316 550700 522317 550764
rect 522251 550699 522317 550700
rect 522254 543965 522314 550699
rect 522251 543964 522317 543965
rect 522251 543900 522252 543964
rect 522316 543900 522317 543964
rect 522251 543899 522317 543900
rect 522067 543692 522133 543693
rect 522067 543628 522068 543692
rect 522132 543628 522133 543692
rect 522067 543627 522133 543628
rect 522070 540973 522130 543627
rect 522067 540972 522133 540973
rect 522067 540908 522068 540972
rect 522132 540908 522133 540972
rect 522067 540907 522133 540908
rect 521883 531452 521949 531453
rect 521883 531388 521884 531452
rect 521948 531388 521949 531452
rect 521883 531387 521949 531388
rect 521886 524517 521946 531387
rect 521883 524516 521949 524517
rect 521883 524452 521884 524516
rect 521948 524452 521949 524516
rect 521883 524451 521949 524452
rect 522804 524454 523404 559898
rect 522067 524244 522133 524245
rect 522067 524180 522068 524244
rect 522132 524180 522133 524244
rect 522067 524179 522133 524180
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522070 521661 522130 524179
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522067 521660 522133 521661
rect 522067 521596 522068 521660
rect 522132 521596 522133 521660
rect 522067 521595 522133 521596
rect 521883 512140 521949 512141
rect 521883 512076 521884 512140
rect 521948 512076 521949 512140
rect 521883 512075 521949 512076
rect 521886 505205 521946 512075
rect 521883 505204 521949 505205
rect 521883 505140 521884 505204
rect 521948 505140 521949 505204
rect 521883 505139 521949 505140
rect 521699 504932 521765 504933
rect 521699 504868 521700 504932
rect 521764 504868 521765 504932
rect 521699 504867 521765 504868
rect 521702 502349 521762 504867
rect 521699 502348 521765 502349
rect 521699 502284 521700 502348
rect 521764 502284 521765 502348
rect 521699 502283 521765 502284
rect 521883 492692 521949 492693
rect 521883 492628 521884 492692
rect 521948 492628 521949 492692
rect 521883 492627 521949 492628
rect 521886 485893 521946 492627
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 521883 485892 521949 485893
rect 521883 485828 521884 485892
rect 521948 485828 521949 485892
rect 521883 485827 521949 485828
rect 521699 485620 521765 485621
rect 521699 485556 521700 485620
rect 521764 485556 521765 485620
rect 521699 485555 521765 485556
rect 521702 476101 521762 485555
rect 521699 476100 521765 476101
rect 521699 476036 521700 476100
rect 521764 476036 521765 476100
rect 521699 476035 521765 476036
rect 522435 476100 522501 476101
rect 522435 476036 522436 476100
rect 522500 476036 522501 476100
rect 522435 476035 522501 476036
rect 522438 466581 522498 476035
rect 522435 466580 522501 466581
rect 522435 466516 522436 466580
rect 522500 466516 522501 466580
rect 522435 466515 522501 466516
rect 522251 466308 522317 466309
rect 522251 466244 522252 466308
rect 522316 466244 522317 466308
rect 522251 466243 522317 466244
rect 522254 463589 522314 466243
rect 522251 463588 522317 463589
rect 522251 463524 522252 463588
rect 522316 463524 522317 463588
rect 522251 463523 522317 463524
rect 521883 454068 521949 454069
rect 521883 454004 521884 454068
rect 521948 454004 521949 454068
rect 521883 454003 521949 454004
rect 521886 447269 521946 454003
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 521883 447268 521949 447269
rect 521883 447204 521884 447268
rect 521948 447204 521949 447268
rect 521883 447203 521949 447204
rect 522067 446996 522133 446997
rect 522067 446932 522068 446996
rect 522132 446932 522133 446996
rect 522067 446931 522133 446932
rect 522070 437610 522130 446931
rect 521702 437550 522130 437610
rect 521702 437477 521762 437550
rect 521699 437476 521765 437477
rect 521699 437412 521700 437476
rect 521764 437412 521765 437476
rect 521699 437411 521765 437412
rect 522251 437476 522317 437477
rect 522251 437412 522252 437476
rect 522316 437412 522317 437476
rect 522251 437411 522317 437412
rect 522254 427957 522314 437411
rect 522251 427956 522317 427957
rect 522251 427892 522252 427956
rect 522316 427892 522317 427956
rect 522251 427891 522317 427892
rect 522067 427684 522133 427685
rect 522067 427620 522068 427684
rect 522132 427620 522133 427684
rect 522067 427619 522133 427620
rect 522070 424965 522130 427619
rect 522067 424964 522133 424965
rect 522067 424900 522068 424964
rect 522132 424900 522133 424964
rect 522067 424899 522133 424900
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 521883 415444 521949 415445
rect 521883 415380 521884 415444
rect 521948 415380 521949 415444
rect 521883 415379 521949 415380
rect 521886 408645 521946 415379
rect 521883 408644 521949 408645
rect 521883 408580 521884 408644
rect 521948 408580 521949 408644
rect 521883 408579 521949 408580
rect 521699 408372 521765 408373
rect 521699 408308 521700 408372
rect 521764 408308 521765 408372
rect 521699 408307 521765 408308
rect 521702 405653 521762 408307
rect 521699 405652 521765 405653
rect 521699 405588 521700 405652
rect 521764 405588 521765 405652
rect 521699 405587 521765 405588
rect 521883 396132 521949 396133
rect 521883 396068 521884 396132
rect 521948 396068 521949 396132
rect 521883 396067 521949 396068
rect 521886 389333 521946 396067
rect 521883 389332 521949 389333
rect 521883 389268 521884 389332
rect 521948 389268 521949 389332
rect 521883 389267 521949 389268
rect 522067 389060 522133 389061
rect 522067 388996 522068 389060
rect 522132 388996 522133 389060
rect 522067 388995 522133 388996
rect 522070 386341 522130 388995
rect 522067 386340 522133 386341
rect 522067 386276 522068 386340
rect 522132 386276 522133 386340
rect 522067 386275 522133 386276
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522251 376820 522317 376821
rect 522251 376756 522252 376820
rect 522316 376756 522317 376820
rect 522251 376755 522317 376756
rect 522254 370021 522314 376755
rect 522251 370020 522317 370021
rect 522251 369956 522252 370020
rect 522316 369956 522317 370020
rect 522251 369955 522317 369956
rect 522067 369748 522133 369749
rect 522067 369684 522068 369748
rect 522132 369684 522133 369748
rect 522067 369683 522133 369684
rect 522070 360090 522130 369683
rect 521886 360030 522130 360090
rect 521886 357373 521946 360030
rect 521883 357372 521949 357373
rect 521883 357308 521884 357372
rect 521948 357308 521949 357372
rect 521883 357307 521949 357308
rect 521699 350572 521765 350573
rect 521699 350508 521700 350572
rect 521764 350508 521765 350572
rect 521699 350507 521765 350508
rect 521702 347717 521762 350507
rect 521699 347716 521765 347717
rect 521699 347652 521700 347716
rect 521764 347652 521765 347716
rect 521699 347651 521765 347652
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 521883 338196 521949 338197
rect 521883 338132 521884 338196
rect 521948 338132 521949 338196
rect 521883 338131 521949 338132
rect 521886 331397 521946 338131
rect 521883 331396 521949 331397
rect 521883 331332 521884 331396
rect 521948 331332 521949 331396
rect 521883 331331 521949 331332
rect 522067 331124 522133 331125
rect 522067 331060 522068 331124
rect 522132 331060 522133 331124
rect 522067 331059 522133 331060
rect 522070 328405 522130 331059
rect 522067 328404 522133 328405
rect 522067 328340 522068 328404
rect 522132 328340 522133 328404
rect 522067 328339 522133 328340
rect 521883 318884 521949 318885
rect 521883 318820 521884 318884
rect 521948 318820 521949 318884
rect 521883 318819 521949 318820
rect 521886 312085 521946 318819
rect 521883 312084 521949 312085
rect 521883 312020 521884 312084
rect 521948 312020 521949 312084
rect 521883 312019 521949 312020
rect 522067 311812 522133 311813
rect 522067 311748 522068 311812
rect 522132 311748 522133 311812
rect 522067 311747 522133 311748
rect 522070 309093 522130 311747
rect 522067 309092 522133 309093
rect 522067 309028 522068 309092
rect 522132 309028 522133 309092
rect 522067 309027 522133 309028
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 521883 302156 521949 302157
rect 521883 302092 521884 302156
rect 521948 302092 521949 302156
rect 521883 302091 521949 302092
rect 521886 292770 521946 302091
rect 521886 292710 522130 292770
rect 522070 289781 522130 292710
rect 522067 289780 522133 289781
rect 522067 289716 522068 289780
rect 522132 289716 522133 289780
rect 522067 289715 522133 289716
rect 521883 280260 521949 280261
rect 521883 280196 521884 280260
rect 521948 280196 521949 280260
rect 521883 280195 521949 280196
rect 521886 273461 521946 280195
rect 521883 273460 521949 273461
rect 521883 273396 521884 273460
rect 521948 273396 521949 273460
rect 521883 273395 521949 273396
rect 522067 273052 522133 273053
rect 522067 272988 522068 273052
rect 522132 272988 522133 273052
rect 522067 272987 522133 272988
rect 522070 270469 522130 272987
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522067 270468 522133 270469
rect 522067 270404 522068 270468
rect 522132 270404 522133 270468
rect 522067 270403 522133 270404
rect 521883 260948 521949 260949
rect 521883 260884 521884 260948
rect 521948 260884 521949 260948
rect 521883 260883 521949 260884
rect 521886 254013 521946 260883
rect 521883 254012 521949 254013
rect 521883 253948 521884 254012
rect 521948 253948 521949 254012
rect 521883 253947 521949 253948
rect 522067 253740 522133 253741
rect 522067 253676 522068 253740
rect 522132 253676 522133 253740
rect 522067 253675 522133 253676
rect 522070 251157 522130 253675
rect 522067 251156 522133 251157
rect 522067 251092 522068 251156
rect 522132 251092 522133 251156
rect 522067 251091 522133 251092
rect 521883 241636 521949 241637
rect 521883 241572 521884 241636
rect 521948 241572 521949 241636
rect 521883 241571 521949 241572
rect 521886 234701 521946 241571
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 521883 234700 521949 234701
rect 521883 234636 521884 234700
rect 521948 234636 521949 234700
rect 521883 234635 521949 234636
rect 522067 234428 522133 234429
rect 522067 234364 522068 234428
rect 522132 234364 522133 234428
rect 522067 234363 522133 234364
rect 522070 227490 522130 234363
rect 521518 227430 522130 227490
rect 522251 227492 522317 227493
rect 521518 224770 521578 227430
rect 522251 227428 522252 227492
rect 522316 227428 522317 227492
rect 522251 227427 522317 227428
rect 521518 224710 521946 224770
rect 521886 222189 521946 224710
rect 521883 222188 521949 222189
rect 521883 222124 521884 222188
rect 521948 222124 521949 222188
rect 521883 222123 521949 222124
rect 522067 212668 522133 212669
rect 522067 212604 522068 212668
rect 522132 212604 522133 212668
rect 522067 212603 522133 212604
rect 522070 212533 522130 212603
rect 522067 212532 522133 212533
rect 522067 212468 522068 212532
rect 522132 212468 522133 212532
rect 522067 212467 522133 212468
rect 521883 206276 521949 206277
rect 521883 206212 521884 206276
rect 521948 206212 521949 206276
rect 521883 206211 521949 206212
rect 521886 200021 521946 206211
rect 521883 200020 521949 200021
rect 521883 199956 521884 200020
rect 521948 199956 521949 200020
rect 521883 199955 521949 199956
rect 521699 190500 521765 190501
rect 521699 190436 521700 190500
rect 521764 190436 521765 190500
rect 521699 190435 521765 190436
rect 521702 186010 521762 190435
rect 521702 185950 521946 186010
rect 521886 176765 521946 185950
rect 522254 181117 522314 227427
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522251 181116 522317 181117
rect 522251 181052 522252 181116
rect 522316 181052 522317 181116
rect 522251 181051 522317 181052
rect 521883 176764 521949 176765
rect 521883 176700 521884 176764
rect 521948 176700 521949 176764
rect 521883 176699 521949 176700
rect 521699 176492 521765 176493
rect 521699 176428 521700 176492
rect 521764 176428 521765 176492
rect 521699 176427 521765 176428
rect 521702 173909 521762 176427
rect 521699 173908 521765 173909
rect 521699 173844 521700 173908
rect 521764 173844 521765 173908
rect 521699 173843 521765 173844
rect 522804 164454 523404 199898
rect 521883 164252 521949 164253
rect 521883 164188 521884 164252
rect 521948 164188 521949 164252
rect 521883 164187 521949 164188
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 521886 157453 521946 164187
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 521883 157452 521949 157453
rect 521883 157388 521884 157452
rect 521948 157388 521949 157452
rect 521883 157387 521949 157388
rect 521699 157180 521765 157181
rect 521699 157116 521700 157180
rect 521764 157116 521765 157180
rect 521699 157115 521765 157116
rect 521702 147661 521762 157115
rect 521699 147660 521765 147661
rect 521699 147596 521700 147660
rect 521764 147596 521765 147660
rect 521699 147595 521765 147596
rect 522435 147660 522501 147661
rect 522435 147596 522436 147660
rect 522500 147596 522501 147660
rect 522435 147595 522501 147596
rect 522438 138141 522498 147595
rect 522435 138140 522501 138141
rect 522435 138076 522436 138140
rect 522500 138076 522501 138140
rect 522435 138075 522501 138076
rect 522251 137868 522317 137869
rect 522251 137804 522252 137868
rect 522316 137804 522317 137868
rect 522251 137803 522317 137804
rect 522254 135149 522314 137803
rect 522251 135148 522317 135149
rect 522251 135084 522252 135148
rect 522316 135084 522317 135148
rect 522251 135083 522317 135084
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 521883 125628 521949 125629
rect 521883 125564 521884 125628
rect 521948 125564 521949 125628
rect 521883 125563 521949 125564
rect 521886 118829 521946 125563
rect 521883 118828 521949 118829
rect 521883 118764 521884 118828
rect 521948 118764 521949 118828
rect 521883 118763 521949 118764
rect 522067 118556 522133 118557
rect 522067 118492 522068 118556
rect 522132 118492 522133 118556
rect 522067 118491 522133 118492
rect 522070 115837 522130 118491
rect 522067 115836 522133 115837
rect 522067 115772 522068 115836
rect 522132 115772 522133 115836
rect 522067 115771 522133 115772
rect 521883 106316 521949 106317
rect 521883 106252 521884 106316
rect 521948 106252 521949 106316
rect 521883 106251 521949 106252
rect 521886 98837 521946 106251
rect 521883 98836 521949 98837
rect 521883 98772 521884 98836
rect 521948 98772 521949 98836
rect 521883 98771 521949 98772
rect 519491 97884 519557 97885
rect 519491 97820 519492 97884
rect 519556 97820 519557 97884
rect 519491 97819 519557 97820
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 516731 29068 516797 29069
rect 516731 29004 516732 29068
rect 516796 29004 516797 29068
rect 516731 29003 516797 29004
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 529062 263669 529122 377622
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 529059 263668 529125 263669
rect 529059 263604 529060 263668
rect 529124 263604 529125 263668
rect 529059 263603 529125 263604
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 531267 181388 531333 181389
rect 531267 181324 531268 181388
rect 531332 181324 531333 181388
rect 531267 181323 531333 181324
rect 531270 180981 531330 181323
rect 531267 180980 531333 180981
rect 531267 180916 531268 180980
rect 531332 180916 531333 180980
rect 531267 180915 531333 180916
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 535499 5812 535565 5813
rect 535499 5748 535500 5812
rect 535564 5748 535565 5812
rect 535499 5747 535565 5748
rect 535502 4045 535562 5747
rect 535499 4044 535565 4045
rect 535499 3980 535500 4044
rect 535564 3980 535565 4044
rect 535499 3979 535565 3980
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 10094 485742 10330 485978
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 17822 485892 18058 485978
rect 17822 485828 17908 485892
rect 17908 485828 17972 485892
rect 17972 485828 18058 485892
rect 17822 485742 18058 485828
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 21134 206262 21370 206498
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 27390 487102 27626 487338
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 33646 487252 33882 487338
rect 33646 487188 33732 487252
rect 33732 487188 33796 487252
rect 33796 487188 33882 487252
rect 33646 487102 33882 487188
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 46710 484382 46946 484618
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 64006 605422 64242 605658
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 61246 206262 61482 206498
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 66766 598622 67002 598858
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83142 604062 83378 604298
rect 80750 598622 80986 598858
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 89030 605572 89266 605658
rect 89030 605508 89116 605572
rect 89116 605508 89180 605572
rect 89180 605508 89266 605572
rect 89030 605422 89266 605508
rect 90134 605572 90370 605658
rect 90134 605508 90220 605572
rect 90220 605508 90284 605572
rect 90284 605508 90370 605572
rect 90134 605422 90370 605508
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108350 604212 108586 604298
rect 108350 604148 108436 604212
rect 108436 604148 108500 604212
rect 108500 604148 108586 604212
rect 108350 604062 108586 604148
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 109638 604742 109874 604978
rect 109638 604212 109874 604298
rect 109638 604148 109724 604212
rect 109724 604148 109788 604212
rect 109788 604148 109874 604212
rect 109638 604062 109874 604148
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 118470 605572 118706 605658
rect 118470 605508 118556 605572
rect 118556 605508 118620 605572
rect 118620 605508 118706 605572
rect 118470 605422 118706 605508
rect 118838 605422 119074 605658
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 128590 605422 128826 605658
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 138342 605422 138578 605658
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 147358 604212 147594 604298
rect 147358 604148 147444 604212
rect 147444 604148 147508 604212
rect 147508 604148 147594 604212
rect 147358 604062 147594 604148
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 157110 605422 157346 605658
rect 157662 605572 157898 605658
rect 157662 605508 157748 605572
rect 157748 605508 157812 605572
rect 157812 605508 157898 605572
rect 157662 605422 157898 605508
rect 157846 604742 158082 604978
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 176430 605572 176666 605658
rect 176430 605508 176516 605572
rect 176516 605508 176580 605572
rect 176580 605508 176666 605572
rect 176430 605422 176666 605508
rect 176798 605422 177034 605658
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 195750 605422 195986 605658
rect 196486 605422 196722 605658
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 204950 604062 205186 604298
rect 205686 604062 205922 604298
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 206974 604742 207210 604978
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 223534 604212 223770 604298
rect 223534 604148 223620 604212
rect 223620 604148 223684 604212
rect 223684 604148 223770 604212
rect 223534 604062 223770 604148
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 224822 604212 225058 604298
rect 224822 604148 224908 604212
rect 224908 604148 224972 604212
rect 224972 604148 225058 604212
rect 224822 604062 225058 604148
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 235862 605422 236098 605658
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 244326 605422 244562 605658
rect 243590 604062 243826 604298
rect 244326 604062 244562 604298
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 253894 605422 254130 605658
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263278 604212 263514 604298
rect 263278 604148 263364 604212
rect 263364 604148 263428 604212
rect 263428 604148 263514 604212
rect 263278 604062 263514 604148
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 264382 604212 264618 604298
rect 264382 604148 264468 604212
rect 264468 604148 264532 604212
rect 264532 604148 264618 604212
rect 264382 604062 264618 604148
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 272846 605422 273082 605658
rect 273214 605422 273450 605658
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281126 604212 281362 604298
rect 281126 604148 281212 604212
rect 281212 604148 281276 604212
rect 281276 604148 281362 604212
rect 281126 604062 281362 604148
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 282966 604212 283202 604298
rect 282966 604148 283052 604212
rect 283052 604148 283116 604212
rect 283116 604148 283202 604212
rect 282966 604062 283202 604148
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 301550 604062 301786 604298
rect 302286 604062 302522 604298
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 320870 604062 321106 604298
rect 321606 604062 321842 604298
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 340190 604062 340426 604298
rect 340926 604062 341162 604298
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 359510 604062 359746 604298
rect 360246 604062 360482 604298
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378462 604212 378698 604298
rect 378462 604148 378548 604212
rect 378548 604148 378612 604212
rect 378612 604148 378698 604212
rect 378462 604062 378698 604148
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 388950 604212 389186 604298
rect 388950 604148 389036 604212
rect 389036 604148 389100 604212
rect 389100 604148 389186 604212
rect 388950 604062 389186 604148
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414342 604212 414578 604298
rect 414342 604148 414428 604212
rect 414428 604148 414492 604212
rect 414492 604148 414578 604212
rect 414342 604062 414578 604148
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 421518 604212 421754 604298
rect 421518 604148 421604 604212
rect 421604 604148 421668 604212
rect 421668 604148 421754 604212
rect 421518 604062 421754 604148
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 428142 604742 428378 604978
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 437710 604742 437946 604978
rect 437158 604212 437394 604298
rect 437158 604148 437244 604212
rect 437244 604148 437308 604212
rect 437308 604148 437394 604212
rect 437158 604062 437394 604148
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 458686 604742 458922 604978
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 476902 600662 477138 600898
rect 404958 599452 405194 599538
rect 404958 599388 405044 599452
rect 405044 599388 405108 599452
rect 405108 599388 405194 599452
rect 404958 599302 405194 599388
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 78910 205052 79146 205138
rect 78910 204988 78996 205052
rect 78996 204988 79060 205052
rect 79060 204988 79146 205052
rect 78910 204902 79146 204988
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 82406 377092 82642 377178
rect 82406 377028 82492 377092
rect 82492 377028 82556 377092
rect 82556 377028 82642 377092
rect 82406 376942 82642 377028
rect 82406 227492 82642 227578
rect 82406 227428 82492 227492
rect 82492 227428 82556 227492
rect 82556 227428 82642 227492
rect 82406 227342 82642 227428
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 76586 5498 76822 5734
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 169438 101542 169674 101778
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 231814 100332 232050 100418
rect 231814 100268 231900 100332
rect 231900 100268 231964 100332
rect 231964 100268 232050 100332
rect 231814 100182 232050 100268
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 241382 101692 241618 101778
rect 241382 101628 241468 101692
rect 241468 101628 241532 101692
rect 241532 101628 241618 101692
rect 241382 101542 241618 101628
rect 241198 100862 241434 101098
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 250950 100182 251186 100418
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 270454 100332 270690 100418
rect 270454 100268 270540 100332
rect 270540 100268 270604 100332
rect 270604 100268 270690 100332
rect 270454 100182 270690 100268
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 273766 100862 274002 101098
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 347734 100332 347970 100418
rect 347734 100268 347820 100332
rect 347820 100268 347884 100332
rect 347884 100268 347970 100332
rect 347734 100182 347970 100268
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 351046 100862 351282 101098
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 395758 101012 395994 101098
rect 395758 100948 395844 101012
rect 395844 100948 395908 101012
rect 395908 100948 395994 101012
rect 395758 100862 395994 100948
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 402750 101012 402986 101098
rect 402750 100948 402836 101012
rect 402836 100948 402900 101012
rect 402900 100948 402986 101012
rect 402750 100862 402986 100948
rect 403670 101012 403906 101098
rect 403670 100948 403756 101012
rect 403756 100948 403820 101012
rect 403820 100948 403906 101012
rect 403670 100862 403906 100948
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 412318 101542 412554 101778
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 466046 3622 466282 3858
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 481502 101012 481738 101098
rect 481502 100948 481588 101012
rect 481588 100948 481652 101012
rect 481652 100948 481738 101012
rect 481502 100862 481738 100948
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 488494 604076 488730 604298
rect 488494 604062 488580 604076
rect 488580 604062 488644 604076
rect 488644 604062 488730 604076
rect 487206 374902 487442 375138
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 491070 597942 491306 598178
rect 491254 404142 491490 404378
rect 489046 378302 489282 378538
rect 488678 374902 488914 375138
rect 486654 208302 486890 208538
rect 486654 206262 486890 206498
rect 486838 145062 487074 145298
rect 486838 144382 487074 144618
rect 488126 232102 488362 232338
rect 488126 187902 488362 188138
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 492174 404142 492410 404378
rect 490886 386462 491122 386698
rect 491806 386462 492042 386698
rect 490150 240942 490386 241178
rect 491438 232102 491674 232338
rect 492174 208302 492410 208538
rect 492174 205582 492410 205818
rect 491806 187902 492042 188138
rect 491254 187222 491490 187458
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 491806 183822 492042 184058
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 493094 598622 493330 598858
rect 494382 507502 494618 507738
rect 493462 476222 493698 476458
rect 494382 476222 494618 476458
rect 494014 451062 494250 451298
rect 494014 448342 494250 448578
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 493094 404142 493330 404378
rect 493462 396662 493698 396898
rect 493094 394622 493330 394858
rect 494382 396662 494618 396898
rect 493646 359942 493882 360178
rect 494382 359942 494618 360178
rect 493830 342262 494066 342498
rect 495118 404142 495354 404378
rect 495302 394622 495538 394858
rect 494750 357902 494986 358138
rect 495486 357902 495722 358138
rect 494934 342942 495170 343178
rect 494566 342262 494802 342498
rect 493278 321862 493514 322098
rect 496958 576862 497194 577098
rect 496774 564622 497010 564858
rect 496774 453102 497010 453338
rect 498614 576862 498850 577098
rect 498614 564622 498850 564858
rect 497878 453102 498114 453338
rect 496958 432702 497194 432938
rect 497878 432702 498114 432938
rect 497694 403462 497930 403698
rect 497326 402782 497562 403018
rect 497142 389862 497378 390098
rect 497142 381022 497378 381258
rect 497142 378302 497378 378538
rect 496222 342942 496458 343178
rect 495854 334782 496090 335018
rect 496590 334782 496826 335018
rect 494198 321862 494434 322098
rect 494014 299422 494250 299658
rect 495118 299422 495354 299658
rect 494566 281742 494802 281978
rect 494934 280382 495170 280618
rect 493646 266102 493882 266338
rect 494750 266782 494986 267018
rect 494750 266102 494986 266338
rect 494750 264062 494986 264298
rect 494198 259302 494434 259538
rect 493278 253182 493514 253418
rect 493830 252502 494066 252738
rect 494750 252502 494986 252738
rect 493462 237542 493698 237778
rect 494382 237542 494618 237778
rect 493646 217142 493882 217378
rect 494382 217142 494618 217378
rect 494014 179742 494250 179978
rect 493094 165462 493330 165698
rect 494382 177022 494618 177258
rect 495302 183822 495538 184058
rect 495486 180422 495722 180658
rect 493094 155942 493330 156178
rect 493094 123302 493330 123538
rect 493094 119902 493330 120138
rect 495118 172942 495354 173178
rect 494750 165462 494986 165698
rect 494934 155942 495170 156178
rect 494750 123302 494986 123538
rect 495118 119902 495354 120138
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 495118 101542 495354 101778
rect 496222 266782 496458 267018
rect 496222 264062 496458 264298
rect 496958 259302 497194 259538
rect 496958 253182 497194 253418
rect 497878 245702 498114 245938
rect 496774 187902 497010 188138
rect 498614 389862 498850 390098
rect 498614 381702 498850 381938
rect 498614 342942 498850 343178
rect 498246 242302 498482 242538
rect 499718 507502 499954 507738
rect 501374 487102 501610 487338
rect 501558 342942 501794 343178
rect 500638 245702 500874 245938
rect 498982 234822 499218 235058
rect 497878 184502 498114 184738
rect 497326 155942 497562 156178
rect 497694 147782 497930 148018
rect 498062 147102 498298 147338
rect 498982 162062 499218 162298
rect 498798 161382 499034 161618
rect 501926 234822 502162 235058
rect 501742 228172 501978 228258
rect 501742 228108 501828 228172
rect 501828 228108 501892 228172
rect 501892 228108 501978 228172
rect 501742 228022 501978 228108
rect 501006 205582 501242 205818
rect 501190 184502 501426 184738
rect 500270 162742 500506 162978
rect 499350 155942 499586 156178
rect 499350 151862 499586 152098
rect 498798 147782 499034 148018
rect 497694 143702 497930 143938
rect 498062 143022 498298 143258
rect 497694 136902 497930 137138
rect 497786 67018 498022 67254
rect 499350 147102 499586 147338
rect 500270 161382 500506 161618
rect 499902 145062 500138 145298
rect 498982 143702 499218 143938
rect 498982 143022 499218 143258
rect 499902 142342 500138 142578
rect 499166 126702 499402 126938
rect 500270 126702 500506 126938
rect 501374 151862 501610 152098
rect 499718 115822 499954 116058
rect 501926 136902 502162 137138
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 496038 3622 496274 3858
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 501926 115822 502162 116058
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 503214 181252 503450 181338
rect 503214 181188 503300 181252
rect 503300 181188 503364 181252
rect 503364 181188 503450 181252
rect 503214 181102 503450 181188
rect 503398 172942 503634 173178
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504502 101542 504738 101778
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 507078 226662 507314 226898
rect 507078 101012 507314 101098
rect 507078 100948 507164 101012
rect 507164 100948 507228 101012
rect 507228 100948 507314 101012
rect 507078 100862 507314 100948
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 515786 696698 516022 696934
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 509102 600662 509338 600898
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 511494 598092 511730 598178
rect 511494 598028 511580 598092
rect 511580 598028 511644 598092
rect 511644 598028 511730 598092
rect 511494 597942 511730 598028
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 511494 226662 511730 226898
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515174 598092 515410 598178
rect 515174 598028 515260 598092
rect 515260 598028 515324 598092
rect 515324 598028 515410 598092
rect 515174 597942 515410 598028
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 513334 100862 513570 101098
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 521982 597942 522218 598178
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 528974 377622 529210 377858
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect 63964 605658 89308 605700
rect 63964 605422 64006 605658
rect 64242 605422 89030 605658
rect 89266 605422 89308 605658
rect 63964 605380 89308 605422
rect 90092 605658 99612 605700
rect 90092 605422 90134 605658
rect 90370 605422 99612 605658
rect 90092 605380 99612 605422
rect 118428 605658 119116 605700
rect 118428 605422 118470 605658
rect 118706 605422 118838 605658
rect 119074 605422 119116 605658
rect 118428 605380 119116 605422
rect 128548 605658 138620 605700
rect 128548 605422 128590 605658
rect 128826 605422 138342 605658
rect 138578 605422 138620 605658
rect 128548 605380 138620 605422
rect 157068 605658 157940 605700
rect 157068 605422 157110 605658
rect 157346 605422 157662 605658
rect 157898 605422 157940 605658
rect 157068 605380 157940 605422
rect 176388 605658 177076 605700
rect 176388 605422 176430 605658
rect 176666 605422 176798 605658
rect 177034 605422 177076 605658
rect 176388 605380 177076 605422
rect 195708 605658 196764 605700
rect 195708 605422 195750 605658
rect 195986 605422 196486 605658
rect 196722 605422 196764 605658
rect 195708 605380 196764 605422
rect 224964 605658 236140 605700
rect 224964 605422 235862 605658
rect 236098 605422 236140 605658
rect 224964 605380 236140 605422
rect 244284 605658 254172 605700
rect 244284 605422 244326 605658
rect 244562 605422 253894 605658
rect 254130 605422 254172 605658
rect 244284 605380 254172 605422
rect 272804 605658 273492 605700
rect 272804 605422 272846 605658
rect 273082 605422 273214 605658
rect 273450 605422 273492 605658
rect 272804 605380 273492 605422
rect 99292 605020 99612 605380
rect 224964 605020 225284 605380
rect 99292 604978 109916 605020
rect 99292 604742 109638 604978
rect 109874 604742 109916 604978
rect 99292 604700 109916 604742
rect 157804 604978 176892 605020
rect 157804 604742 157846 604978
rect 158082 604742 176892 604978
rect 157804 604700 176892 604742
rect 206932 604978 225284 605020
rect 206932 604742 206974 604978
rect 207210 604742 225284 604978
rect 206932 604700 225284 604742
rect 176572 604340 176892 604700
rect 398476 604340 398980 605020
rect 428100 604978 437988 605020
rect 428100 604742 428142 604978
rect 428378 604742 437710 604978
rect 437946 604742 437988 604978
rect 428100 604700 437988 604742
rect 458644 604978 476444 605020
rect 458644 604742 458686 604978
rect 458922 604742 476444 604978
rect 458644 604700 476444 604742
rect 476124 604340 476444 604700
rect 83100 604298 108628 604340
rect 83100 604062 83142 604298
rect 83378 604062 108350 604298
rect 108586 604062 108628 604298
rect 83100 604020 108628 604062
rect 109596 604298 147636 604340
rect 109596 604062 109638 604298
rect 109874 604062 147358 604298
rect 147594 604062 147636 604298
rect 109596 604020 147636 604062
rect 176572 604298 205228 604340
rect 176572 604062 204950 604298
rect 205186 604062 205228 604298
rect 176572 604020 205228 604062
rect 205644 604298 223812 604340
rect 205644 604062 205686 604298
rect 205922 604062 223534 604298
rect 223770 604062 223812 604298
rect 205644 604020 223812 604062
rect 224780 604298 243868 604340
rect 224780 604062 224822 604298
rect 225058 604062 243590 604298
rect 243826 604062 243868 604298
rect 224780 604020 243868 604062
rect 244284 604298 263556 604340
rect 244284 604062 244326 604298
rect 244562 604062 263278 604298
rect 263514 604062 263556 604298
rect 244284 604020 263556 604062
rect 264340 604298 281404 604340
rect 264340 604062 264382 604298
rect 264618 604062 281126 604298
rect 281362 604062 281404 604298
rect 264340 604020 281404 604062
rect 282924 604298 301828 604340
rect 282924 604062 282966 604298
rect 283202 604062 301550 604298
rect 301786 604062 301828 604298
rect 282924 604020 301828 604062
rect 302244 604298 321148 604340
rect 302244 604062 302286 604298
rect 302522 604062 320870 604298
rect 321106 604062 321148 604298
rect 302244 604020 321148 604062
rect 321564 604298 340468 604340
rect 321564 604062 321606 604298
rect 321842 604062 340190 604298
rect 340426 604062 340468 604298
rect 321564 604020 340468 604062
rect 340884 604298 359788 604340
rect 340884 604062 340926 604298
rect 341162 604062 359510 604298
rect 359746 604062 359788 604298
rect 340884 604020 359788 604062
rect 360204 604298 378740 604340
rect 360204 604062 360246 604298
rect 360482 604062 378462 604298
rect 378698 604062 378740 604298
rect 360204 604020 378740 604062
rect 388908 604298 414620 604340
rect 388908 604062 388950 604298
rect 389186 604062 414342 604298
rect 414578 604062 414620 604298
rect 388908 604020 414620 604062
rect 421476 604298 437436 604340
rect 421476 604062 421518 604298
rect 421754 604062 437158 604298
rect 437394 604062 437436 604298
rect 421476 604020 437436 604062
rect 476124 604298 488772 604340
rect 476124 604062 488494 604298
rect 488730 604062 488772 604298
rect 476124 604020 488772 604062
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect 476860 600898 509380 600940
rect 476860 600662 476902 600898
rect 477138 600662 509102 600898
rect 509338 600662 509380 600898
rect 476860 600620 509380 600662
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599538 526586 599734
rect 58822 599498 404958 599538
rect -4756 599476 404958 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 404916 599302 404958 599476
rect 405194 599498 526586 599538
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect 405194 599476 588680 599498
rect 405194 599302 405236 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect 404916 599080 405236 599302
rect 404732 598900 405236 599080
rect 66724 598858 81028 598900
rect 66724 598622 66766 598858
rect 67002 598622 80750 598858
rect 80986 598622 81028 598858
rect 66724 598580 81028 598622
rect 404732 598580 420692 598900
rect 420372 598220 420692 598580
rect 424420 598580 426212 598900
rect 493052 598858 497236 598900
rect 493052 598622 493094 598858
rect 493330 598622 497236 598858
rect 493052 598580 497236 598622
rect 420372 597900 422348 598220
rect 422028 597540 422348 597900
rect 424420 597540 424740 598580
rect 425892 598220 426212 598580
rect 496916 598220 497236 598580
rect 425892 598178 491348 598220
rect 425892 597942 491070 598178
rect 491306 597942 491348 598178
rect 425892 597900 491348 597942
rect 496916 598178 511772 598220
rect 496916 597942 511494 598178
rect 511730 597942 511772 598178
rect 496916 597900 511772 597942
rect 515132 598178 522260 598220
rect 515132 597942 515174 598178
rect 515410 597942 521982 598178
rect 522218 597942 522260 598178
rect 515132 597900 522260 597942
rect 422028 597220 424740 597540
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect 496916 577098 498892 577140
rect 496916 576862 496958 577098
rect 497194 576862 498614 577098
rect 498850 576862 498892 577098
rect 496916 576820 498892 576862
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect 496732 564858 498892 564900
rect 496732 564622 496774 564858
rect 497010 564622 498614 564858
rect 498850 564622 498892 564858
rect 496732 564580 498892 564622
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect 494340 507738 499996 507780
rect 494340 507502 494382 507738
rect 494618 507502 499718 507738
rect 499954 507502 499996 507738
rect 494340 507460 499996 507502
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect 27348 487338 33924 487380
rect 27348 487102 27390 487338
rect 27626 487102 33646 487338
rect 33882 487102 33924 487338
rect 27348 487060 33924 487102
rect 489556 487060 495580 487380
rect 57708 486380 60420 486700
rect 57708 486020 58028 486380
rect 10052 485978 18100 486020
rect 10052 485742 10094 485978
rect 10330 485742 17822 485978
rect 18058 485742 18100 485978
rect 10052 485700 18100 485742
rect 52924 485700 58028 486020
rect 60100 486020 60420 486380
rect 60836 486380 62996 486700
rect 60836 486020 61156 486380
rect 60100 485700 61156 486020
rect 62676 486020 62996 486380
rect 95244 486380 98324 486700
rect 62676 485700 84892 486020
rect 52924 484660 53244 485700
rect 46668 484618 53244 484660
rect 46668 484382 46710 484618
rect 46946 484382 53244 484618
rect 46668 484340 53244 484382
rect 84572 484660 84892 485700
rect 95244 484660 95564 486380
rect 84572 484340 95564 484660
rect 98004 484660 98324 486380
rect 489556 484660 489876 487060
rect 495260 486700 495580 487060
rect 499492 487338 501652 487380
rect 499492 487102 501374 487338
rect 501610 487102 501652 487338
rect 499492 487060 501652 487102
rect 499492 486700 499812 487060
rect 495260 486380 499812 486700
rect 98004 484340 104948 484660
rect 104628 483980 104948 484340
rect 488268 484340 489876 484660
rect 488268 483980 488588 484340
rect 104628 483660 108444 483980
rect 108124 482620 108444 483660
rect 109044 483660 114700 483980
rect 109044 482620 109364 483660
rect 108124 482300 109364 482620
rect 114380 482620 114700 483660
rect 115116 483660 127764 483980
rect 115116 482620 115436 483660
rect 114380 482300 115436 482620
rect 127444 482620 127764 483660
rect 128364 483660 134020 483980
rect 128364 482620 128684 483660
rect 127444 482300 128684 482620
rect 133700 482620 134020 483660
rect 134436 483660 147084 483980
rect 134436 482620 134756 483660
rect 133700 482300 134756 482620
rect 146764 482620 147084 483660
rect 147684 483660 153340 483980
rect 147684 482620 148004 483660
rect 146764 482300 148004 482620
rect 153020 482620 153340 483660
rect 153756 483660 166404 483980
rect 153756 482620 154076 483660
rect 153020 482300 154076 482620
rect 166084 482620 166404 483660
rect 167004 483660 172660 483980
rect 167004 482620 167324 483660
rect 166084 482300 167324 482620
rect 172340 482620 172660 483660
rect 173076 483660 185724 483980
rect 173076 482620 173396 483660
rect 172340 482300 173396 482620
rect 185404 482620 185724 483660
rect 186324 483660 191980 483980
rect 186324 482620 186644 483660
rect 185404 482300 186644 482620
rect 191660 482620 191980 483660
rect 192396 483660 205044 483980
rect 192396 482620 192716 483660
rect 191660 482300 192716 482620
rect 204724 482620 205044 483660
rect 205644 483660 211300 483980
rect 205644 482620 205964 483660
rect 204724 482300 205964 482620
rect 210980 482620 211300 483660
rect 211716 483660 224364 483980
rect 211716 482620 212036 483660
rect 210980 482300 212036 482620
rect 224044 482620 224364 483660
rect 224964 483660 230620 483980
rect 224964 482620 225284 483660
rect 224044 482300 225284 482620
rect 230300 482620 230620 483660
rect 231036 483660 243684 483980
rect 231036 482620 231356 483660
rect 230300 482300 231356 482620
rect 243364 482620 243684 483660
rect 244284 483660 249940 483980
rect 244284 482620 244604 483660
rect 243364 482300 244604 482620
rect 249620 482620 249940 483660
rect 250356 483660 263004 483980
rect 250356 482620 250676 483660
rect 249620 482300 250676 482620
rect 262684 482620 263004 483660
rect 263604 483660 269260 483980
rect 263604 482620 263924 483660
rect 262684 482300 263924 482620
rect 268940 482620 269260 483660
rect 269676 483660 282324 483980
rect 269676 482620 269996 483660
rect 268940 482300 269996 482620
rect 282004 482620 282324 483660
rect 282924 483660 288580 483980
rect 282924 482620 283244 483660
rect 282004 482300 283244 482620
rect 288260 482620 288580 483660
rect 288996 483660 301644 483980
rect 288996 482620 289316 483660
rect 288260 482300 289316 482620
rect 301324 482620 301644 483660
rect 302244 483660 307900 483980
rect 302244 482620 302564 483660
rect 301324 482300 302564 482620
rect 307580 482620 307900 483660
rect 308316 483660 320964 483980
rect 308316 482620 308636 483660
rect 307580 482300 308636 482620
rect 320644 482620 320964 483660
rect 321564 483660 327220 483980
rect 321564 482620 321884 483660
rect 320644 482300 321884 482620
rect 326900 482620 327220 483660
rect 327636 483660 340284 483980
rect 327636 482620 327956 483660
rect 326900 482300 327956 482620
rect 339964 482620 340284 483660
rect 340884 483660 346540 483980
rect 340884 482620 341204 483660
rect 339964 482300 341204 482620
rect 346220 482620 346540 483660
rect 346956 483660 359604 483980
rect 346956 482620 347276 483660
rect 346220 482300 347276 482620
rect 359284 482620 359604 483660
rect 360204 483660 365860 483980
rect 360204 482620 360524 483660
rect 359284 482300 360524 482620
rect 365540 482620 365860 483660
rect 366276 483660 378924 483980
rect 366276 482620 366596 483660
rect 365540 482300 366596 482620
rect 378604 482620 378924 483660
rect 379524 483660 385180 483980
rect 379524 482620 379844 483660
rect 378604 482300 379844 482620
rect 384860 482620 385180 483660
rect 385596 483660 398244 483980
rect 385596 482620 385916 483660
rect 384860 482300 385916 482620
rect 397924 482620 398244 483660
rect 398844 483660 404500 483980
rect 398844 482620 399164 483660
rect 397924 482300 399164 482620
rect 404180 482620 404500 483660
rect 404916 483660 417564 483980
rect 404916 482620 405236 483660
rect 404180 482300 405236 482620
rect 417244 482620 417564 483660
rect 418164 483660 423820 483980
rect 418164 482620 418484 483660
rect 417244 482300 418484 482620
rect 423500 482620 423820 483660
rect 424236 483660 436884 483980
rect 424236 482620 424556 483660
rect 423500 482300 424556 482620
rect 436564 482620 436884 483660
rect 437484 483660 443140 483980
rect 437484 482620 437804 483660
rect 436564 482300 437804 482620
rect 442820 482620 443140 483660
rect 443556 483660 456204 483980
rect 443556 482620 443876 483660
rect 442820 482300 443876 482620
rect 455884 482620 456204 483660
rect 456804 483660 462460 483980
rect 456804 482620 457124 483660
rect 455884 482300 457124 482620
rect 462140 482620 462460 483660
rect 462876 483660 475524 483980
rect 462876 482620 463196 483660
rect 475204 483300 475524 483660
rect 478700 483660 488588 483980
rect 478700 483300 479020 483660
rect 475204 482980 479020 483300
rect 462140 482300 463196 482620
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect 493420 476458 494660 476500
rect 493420 476222 493462 476458
rect 493698 476222 494382 476458
rect 494618 476222 494660 476458
rect 493420 476180 494660 476222
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect 496732 453338 498156 453380
rect 496732 453102 496774 453338
rect 497010 453102 497878 453338
rect 498114 453102 498156 453338
rect 496732 453060 498156 453102
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect 493972 451298 494660 451340
rect 493972 451062 494014 451298
rect 494250 451062 494660 451298
rect 493972 451020 494660 451062
rect 494340 448620 494660 451020
rect 493972 448578 494660 448620
rect 493972 448342 494014 448578
rect 494250 448342 494660 448578
rect 493972 448300 494660 448342
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 496916 432938 498156 432980
rect 496916 432702 496958 432938
rect 497194 432702 497878 432938
rect 498114 432702 498156 432938
rect 496916 432660 498156 432702
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect 491212 404378 492452 404420
rect 491212 404142 491254 404378
rect 491490 404142 492174 404378
rect 492410 404142 492452 404378
rect 491212 404100 492452 404142
rect 493052 404378 495396 404420
rect 493052 404142 493094 404378
rect 493330 404142 495118 404378
rect 495354 404142 495396 404378
rect 493052 404100 495396 404142
rect 497100 403698 497972 403740
rect 497100 403462 497694 403698
rect 497930 403462 497972 403698
rect 497100 403420 497972 403462
rect 497100 403060 497420 403420
rect 497100 403018 497604 403060
rect 497100 402782 497326 403018
rect 497562 402782 497604 403018
rect 497100 402740 497604 402782
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 493420 396898 494660 396940
rect 493420 396662 493462 396898
rect 493698 396662 494382 396898
rect 494618 396662 494660 396898
rect 493420 396620 494660 396662
rect 493052 394858 495580 394900
rect 493052 394622 493094 394858
rect 493330 394622 495302 394858
rect 495538 394622 495580 394858
rect 493052 394580 495580 394622
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect 497100 390098 498892 390140
rect 497100 389862 497142 390098
rect 497378 389862 498614 390098
rect 498850 389862 498892 390098
rect 497100 389820 498892 389862
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect 490844 386698 492084 386740
rect 490844 386462 490886 386698
rect 491122 386462 491806 386698
rect 492042 386462 492084 386698
rect 490844 386420 492084 386462
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect 497100 381938 498892 381980
rect 497100 381702 498614 381938
rect 498850 381702 498892 381938
rect 497100 381660 498892 381702
rect 497100 381258 497420 381660
rect 497100 381022 497142 381258
rect 497378 381022 497420 381258
rect 497100 380980 497420 381022
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect 489004 378538 497420 378580
rect 489004 378302 489046 378538
rect 489282 378302 497142 378538
rect 497378 378302 497420 378538
rect 489004 378260 497420 378302
rect 510532 378260 520236 378580
rect 176572 377580 186276 377900
rect 82364 377178 89676 377220
rect 82364 376942 82406 377178
rect 82642 376942 89676 377178
rect 82364 376900 89676 376942
rect 89356 376540 89676 376900
rect 89356 376220 96852 376540
rect 96532 375180 96852 376220
rect 105916 376220 116172 376540
rect 105916 375180 106236 376220
rect 96532 374860 106236 375180
rect 115852 375180 116172 376220
rect 125236 376220 135492 376540
rect 125236 375180 125556 376220
rect 115852 374860 125556 375180
rect 135172 375180 135492 376220
rect 144556 376220 154812 376540
rect 144556 375180 144876 376220
rect 135172 374860 144876 375180
rect 154492 375180 154812 376220
rect 163876 376220 174132 376540
rect 163876 375180 164196 376220
rect 154492 374860 164196 375180
rect 173812 374500 174132 376220
rect 176572 374500 176892 377580
rect 185956 376540 186276 377580
rect 195892 377580 205596 377900
rect 185956 376220 193452 376540
rect 173812 374180 176892 374500
rect 193132 374500 193452 376220
rect 195892 374500 196212 377580
rect 205276 376540 205596 377580
rect 215212 377580 224916 377900
rect 205276 376220 212772 376540
rect 193132 374180 196212 374500
rect 212452 374500 212772 376220
rect 215212 374500 215532 377580
rect 224596 376540 224916 377580
rect 234532 377580 244236 377900
rect 224596 376220 232092 376540
rect 212452 374180 215532 374500
rect 231772 374500 232092 376220
rect 234532 374500 234852 377580
rect 243916 376540 244236 377580
rect 253852 377580 263556 377900
rect 243916 376220 251412 376540
rect 231772 374180 234852 374500
rect 251092 374500 251412 376220
rect 253852 374500 254172 377580
rect 263236 376540 263556 377580
rect 273172 377580 282876 377900
rect 263236 376220 270732 376540
rect 251092 374180 254172 374500
rect 270412 374500 270732 376220
rect 273172 374500 273492 377580
rect 282556 376540 282876 377580
rect 292492 377580 302196 377900
rect 282556 376220 290052 376540
rect 270412 374180 273492 374500
rect 289732 374500 290052 376220
rect 292492 374500 292812 377580
rect 301876 376540 302196 377580
rect 311812 377580 321516 377900
rect 301876 376220 309372 376540
rect 289732 374180 292812 374500
rect 309052 374500 309372 376220
rect 311812 374500 312132 377580
rect 321196 376540 321516 377580
rect 331132 377580 340836 377900
rect 321196 376220 328692 376540
rect 309052 374180 312132 374500
rect 328372 374500 328692 376220
rect 331132 374500 331452 377580
rect 340516 376540 340836 377580
rect 350452 377580 360156 377900
rect 340516 376220 348012 376540
rect 328372 374180 331452 374500
rect 347692 374500 348012 376220
rect 350452 374500 350772 377580
rect 359836 376540 360156 377580
rect 369772 377580 379476 377900
rect 359836 376220 367332 376540
rect 347692 374180 350772 374500
rect 367012 374500 367332 376220
rect 369772 374500 370092 377580
rect 379156 376540 379476 377580
rect 389092 377580 398796 377900
rect 379156 376220 386652 376540
rect 367012 374180 370092 374500
rect 386332 374500 386652 376220
rect 389092 374500 389412 377580
rect 398476 376540 398796 377580
rect 408412 377580 418116 377900
rect 398476 376220 405972 376540
rect 386332 374180 389412 374500
rect 405652 374500 405972 376220
rect 408412 374500 408732 377580
rect 417796 376540 418116 377580
rect 427732 377580 437436 377900
rect 417796 376220 425292 376540
rect 405652 374180 408732 374500
rect 424972 374500 425292 376220
rect 427732 374500 428052 377580
rect 437116 376540 437436 377580
rect 447052 377580 456756 377900
rect 437116 376220 444612 376540
rect 424972 374180 428052 374500
rect 444292 374500 444612 376220
rect 447052 374500 447372 377580
rect 456436 376540 456756 377580
rect 466372 377580 474972 377900
rect 456436 376220 463932 376540
rect 444292 374180 447372 374500
rect 463612 374500 463932 376220
rect 466372 374500 466692 377580
rect 474652 377220 474972 377580
rect 510532 377220 510852 378260
rect 474652 376900 476260 377220
rect 475940 376540 476260 376900
rect 481460 376900 486012 377220
rect 481460 376540 481780 376900
rect 475940 376220 481780 376540
rect 485692 376540 486012 376900
rect 491028 376900 510852 377220
rect 491028 376540 491348 376900
rect 485692 376220 491348 376540
rect 519916 376540 520236 378260
rect 524332 377858 529252 377900
rect 524332 377622 528974 377858
rect 529210 377622 529252 377858
rect 524332 377580 529252 377622
rect 524332 376540 524652 377580
rect 519916 376220 524652 376540
rect 487164 375138 488956 375180
rect 487164 374902 487206 375138
rect 487442 374902 488678 375138
rect 488914 374902 488956 375138
rect 487164 374860 488956 374902
rect 463612 374180 466692 374500
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect 493604 360178 494660 360220
rect 493604 359942 493646 360178
rect 493882 359942 494382 360178
rect 494618 359942 494660 360178
rect 493604 359900 494660 359942
rect 494708 358138 495764 358180
rect 494708 357902 494750 358138
rect 494986 357902 495486 358138
rect 495722 357902 495764 358138
rect 494708 357860 495764 357902
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect 494892 343178 496500 343220
rect 494892 342942 494934 343178
rect 495170 342942 496222 343178
rect 496458 342942 496500 343178
rect 494892 342900 496500 342942
rect 498572 343178 501836 343220
rect 498572 342942 498614 343178
rect 498850 342942 501558 343178
rect 501794 342942 501836 343178
rect 498572 342900 501836 342942
rect 493788 342498 494844 342540
rect 493788 342262 493830 342498
rect 494066 342262 494566 342498
rect 494802 342262 494844 342498
rect 493788 342220 494844 342262
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect 495812 335018 496868 335060
rect 495812 334782 495854 335018
rect 496090 334782 496590 335018
rect 496826 334782 496868 335018
rect 495812 334740 496868 334782
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect 493236 322098 494476 322140
rect 493236 321862 493278 322098
rect 493514 321862 494198 322098
rect 494434 321862 494476 322098
rect 493236 321820 494476 321862
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect 493972 299658 495396 299700
rect 493972 299422 494014 299658
rect 494250 299422 495118 299658
rect 495354 299422 495396 299658
rect 493972 299380 495396 299422
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect 494524 281978 494844 282020
rect 494524 281742 494566 281978
rect 494802 281742 494844 281978
rect 494524 280660 494844 281742
rect 494524 280618 495212 280660
rect 494524 280382 494934 280618
rect 495170 280382 495212 280618
rect 494524 280340 495212 280382
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect 494708 267018 496500 267060
rect 494708 266782 494750 267018
rect 494986 266782 496222 267018
rect 496458 266782 496500 267018
rect 494708 266740 496500 266782
rect 493604 266338 495028 266380
rect 493604 266102 493646 266338
rect 493882 266102 494750 266338
rect 494986 266102 495028 266338
rect 493604 266060 495028 266102
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect 494708 264298 496500 264340
rect 494708 264062 494750 264298
rect 494986 264062 496222 264298
rect 496458 264062 496500 264298
rect 494708 264020 496500 264062
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect 494156 259538 497236 259580
rect 494156 259302 494198 259538
rect 494434 259302 496958 259538
rect 497194 259302 497236 259538
rect 494156 259260 497236 259302
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect 493236 253418 497236 253460
rect 493236 253182 493278 253418
rect 493514 253182 496958 253418
rect 497194 253182 497236 253418
rect 493236 253140 497236 253182
rect 493788 252738 495028 252780
rect 493788 252502 493830 252738
rect 494066 252502 494750 252738
rect 494986 252502 495028 252738
rect 493788 252460 495028 252502
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect 497836 245938 500916 245980
rect 497836 245702 497878 245938
rect 498114 245702 500638 245938
rect 500874 245702 500916 245938
rect 497836 245660 500916 245702
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect 498204 242538 498708 242580
rect 498204 242302 498246 242538
rect 498482 242302 498708 242538
rect 498204 242260 498708 242302
rect 498388 241220 498708 242260
rect 490108 241178 498708 241220
rect 490108 240942 490150 241178
rect 490386 240942 498708 241178
rect 490108 240900 498708 240942
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect 493420 237778 494660 237820
rect 493420 237542 493462 237778
rect 493698 237542 494382 237778
rect 494618 237542 494660 237778
rect 493420 237500 494660 237542
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect 498940 235058 502204 235100
rect 498940 234822 498982 235058
rect 499218 234822 501926 235058
rect 502162 234822 502204 235058
rect 498940 234780 502204 234822
rect 488084 232338 491716 232380
rect 488084 232102 488126 232338
rect 488362 232102 491438 232338
rect 491674 232102 491716 232338
rect 488084 232060 491716 232102
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect 99108 227980 125556 228300
rect 82364 227578 96668 227620
rect 82364 227342 82406 227578
rect 82642 227342 96668 227578
rect 82364 227300 96668 227342
rect 96348 226940 96668 227300
rect 99108 226940 99428 227980
rect 96348 226620 99428 226940
rect 125236 226940 125556 227980
rect 127996 227980 144876 228300
rect 127996 226940 128316 227980
rect 125236 226620 128316 226940
rect 144556 226940 144876 227980
rect 147316 227980 164196 228300
rect 147316 226940 147636 227980
rect 144556 226620 147636 226940
rect 163876 226940 164196 227980
rect 166636 227980 183516 228300
rect 166636 226940 166956 227980
rect 163876 226620 166956 226940
rect 183196 226940 183516 227980
rect 185956 227980 196028 228300
rect 185956 226940 186276 227980
rect 183196 226620 186276 226940
rect 195708 226940 196028 227980
rect 199940 227980 209828 228300
rect 199940 226940 200260 227980
rect 195708 226620 200260 226940
rect 209508 226940 209828 227980
rect 219260 227980 229148 228300
rect 219260 226940 219580 227980
rect 209508 226620 219580 226940
rect 228828 226940 229148 227980
rect 238580 227980 248468 228300
rect 238580 226940 238900 227980
rect 228828 226620 238900 226940
rect 248148 226940 248468 227980
rect 257900 227980 267788 228300
rect 257900 226940 258220 227980
rect 248148 226620 258220 226940
rect 267468 226940 267788 227980
rect 277220 227980 287108 228300
rect 277220 226940 277540 227980
rect 267468 226620 277540 226940
rect 286788 226940 287108 227980
rect 296540 227980 306428 228300
rect 296540 226940 296860 227980
rect 286788 226620 296860 226940
rect 306108 226940 306428 227980
rect 315860 227980 325748 228300
rect 315860 226940 316180 227980
rect 306108 226620 316180 226940
rect 325428 226940 325748 227980
rect 335180 227980 345068 228300
rect 335180 226940 335500 227980
rect 325428 226620 335500 226940
rect 344748 226940 345068 227980
rect 354500 227980 364388 228300
rect 354500 226940 354820 227980
rect 344748 226620 354820 226940
rect 364068 226940 364388 227980
rect 373820 227980 383708 228300
rect 373820 226940 374140 227980
rect 364068 226620 374140 226940
rect 383388 226940 383708 227980
rect 393140 227980 403028 228300
rect 393140 226940 393460 227980
rect 383388 226620 393460 226940
rect 402708 226940 403028 227980
rect 412460 227980 422348 228300
rect 412460 226940 412780 227980
rect 402708 226620 412780 226940
rect 422028 226940 422348 227980
rect 431780 227980 441668 228300
rect 431780 226940 432100 227980
rect 422028 226620 432100 226940
rect 441348 226940 441668 227980
rect 451100 227980 460988 228300
rect 451100 226940 451420 227980
rect 441348 226620 451420 226940
rect 460668 226940 460988 227980
rect 470420 227980 472212 228300
rect 470420 226940 470740 227980
rect 471892 227620 472212 227980
rect 481460 228258 502020 228300
rect 481460 228022 501742 228258
rect 501978 228022 502020 228258
rect 481460 227980 502020 228022
rect 481460 227620 481780 227980
rect 471892 227300 481780 227620
rect 460668 226620 470740 226940
rect 481276 226620 481780 227300
rect 507036 226898 511772 226940
rect 507036 226662 507078 226898
rect 507314 226662 511494 226898
rect 511730 226662 511772 226898
rect 507036 226620 511772 226662
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect 493604 217378 494660 217420
rect 493604 217142 493646 217378
rect 493882 217142 494382 217378
rect 494618 217142 494660 217378
rect 493604 217100 494660 217142
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect 486612 208538 492452 208580
rect 486612 208302 486654 208538
rect 486890 208302 492174 208538
rect 492410 208302 492452 208538
rect 486612 208260 492452 208302
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -35879 206498 26380 206540
rect -35879 206262 21134 206498
rect 21370 206262 26380 206498
rect -35879 206220 26380 206262
rect 26060 205180 26380 206220
rect 50716 206498 61524 206540
rect 50716 206262 61246 206498
rect 61482 206262 61524 206498
rect 50716 206220 61524 206262
rect 91564 206220 94092 206540
rect 50716 205180 51036 206220
rect 91564 205180 91884 206220
rect 26060 204860 51036 205180
rect 78868 205138 91884 205180
rect 78868 204902 78910 205138
rect 79146 204902 91884 205138
rect 78868 204860 91884 204902
rect 93772 205180 94092 206220
rect 94692 206220 103660 206540
rect 94692 205180 95012 206220
rect 93772 204860 95012 205180
rect 103340 205180 103660 206220
rect 112908 206220 122980 206540
rect 112908 205180 113228 206220
rect 103340 204860 113228 205180
rect 122660 205180 122980 206220
rect 132228 206220 142300 206540
rect 132228 205180 132548 206220
rect 122660 204860 132548 205180
rect 141980 205180 142300 206220
rect 151548 206220 161620 206540
rect 151548 205180 151868 206220
rect 141980 204860 151868 205180
rect 161300 205180 161620 206220
rect 170868 206220 180940 206540
rect 170868 205180 171188 206220
rect 161300 204860 171188 205180
rect 180620 205180 180940 206220
rect 190188 206220 200260 206540
rect 190188 205180 190508 206220
rect 180620 204860 190508 205180
rect 199940 205180 200260 206220
rect 209508 206220 219580 206540
rect 209508 205180 209828 206220
rect 199940 204860 209828 205180
rect 219260 205180 219580 206220
rect 228828 206220 238900 206540
rect 228828 205180 229148 206220
rect 219260 204860 229148 205180
rect 238580 205180 238900 206220
rect 248148 206220 258220 206540
rect 248148 205180 248468 206220
rect 238580 204860 248468 205180
rect 257900 205180 258220 206220
rect 267468 206220 277540 206540
rect 267468 205180 267788 206220
rect 257900 204860 267788 205180
rect 277220 205180 277540 206220
rect 286788 206220 296860 206540
rect 286788 205180 287108 206220
rect 277220 204860 287108 205180
rect 296540 205180 296860 206220
rect 306108 206220 316180 206540
rect 306108 205180 306428 206220
rect 296540 204860 306428 205180
rect 315860 205180 316180 206220
rect 325428 206220 335500 206540
rect 325428 205180 325748 206220
rect 315860 204860 325748 205180
rect 335180 205180 335500 206220
rect 344748 206220 354820 206540
rect 344748 205180 345068 206220
rect 335180 204860 345068 205180
rect 354500 205180 354820 206220
rect 364068 206220 374140 206540
rect 364068 205180 364388 206220
rect 354500 204860 364388 205180
rect 373820 205180 374140 206220
rect 383388 206220 393460 206540
rect 383388 205180 383708 206220
rect 373820 204860 383708 205180
rect 393140 205180 393460 206220
rect 402708 206220 412780 206540
rect 402708 205180 403028 206220
rect 393140 204860 403028 205180
rect 412460 205180 412780 206220
rect 422028 206220 432100 206540
rect 422028 205180 422348 206220
rect 412460 204860 422348 205180
rect 431780 205180 432100 206220
rect 441348 206220 451420 206540
rect 441348 205180 441668 206220
rect 431780 204860 441668 205180
rect 451100 205180 451420 206220
rect 460668 206220 470740 206540
rect 460668 205180 460988 206220
rect 451100 204860 460988 205180
rect 470420 205180 470740 206220
rect 483116 206498 486932 206540
rect 483116 206262 486654 206498
rect 486890 206262 486932 206498
rect 483116 206220 486932 206262
rect 483116 205180 483436 206220
rect 492132 205818 501284 205860
rect 492132 205582 492174 205818
rect 492410 205582 501006 205818
rect 501242 205582 501284 205818
rect 492132 205540 501284 205582
rect 470420 204860 483436 205180
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect 488084 188138 488404 188180
rect 488084 187902 488126 188138
rect 488362 187902 488404 188138
rect 488084 187500 488404 187902
rect 491764 188138 497052 188180
rect 491764 187902 491806 188138
rect 492042 187902 496774 188138
rect 497010 187902 497052 188138
rect 491764 187860 497052 187902
rect 488084 187458 491532 187500
rect 488084 187222 491254 187458
rect 491490 187222 491532 187458
rect 488084 187180 491532 187222
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect 497836 184738 501468 184780
rect 497836 184502 497878 184738
rect 498114 184502 501190 184738
rect 501426 184502 501468 184738
rect 497836 184460 501468 184502
rect 491764 184058 495580 184100
rect 491764 183822 491806 184058
rect 492042 183822 495302 184058
rect 495538 183822 495580 184058
rect 491764 183780 495580 183822
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect 495444 181338 503492 181380
rect 495444 181102 503214 181338
rect 503450 181102 503492 181338
rect 495444 181060 503492 181102
rect 495444 180658 495764 181060
rect 495444 180422 495486 180658
rect 495722 180422 495764 180658
rect 495444 180380 495764 180422
rect 493972 179978 494660 180020
rect 493972 179742 494014 179978
rect 494250 179742 494660 179978
rect 493972 179700 494660 179742
rect 494340 177258 494660 179700
rect 494340 177022 494382 177258
rect 494618 177022 494660 177258
rect 494340 176980 494660 177022
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect 495076 173178 503676 173220
rect 495076 172942 495118 173178
rect 495354 172942 503398 173178
rect 503634 172942 503676 173178
rect 495076 172900 503676 172942
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect 493052 165698 495028 165740
rect 493052 165462 493094 165698
rect 493330 165462 494750 165698
rect 494986 165462 495028 165698
rect 493052 165420 495028 165462
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect 500228 162978 500548 163020
rect 500228 162742 500270 162978
rect 500506 162742 500548 162978
rect 498756 162298 499260 162340
rect 498756 162062 498982 162298
rect 499218 162062 499260 162298
rect 498756 162020 499260 162062
rect 498756 161618 499076 162020
rect 498756 161382 498798 161618
rect 499034 161382 499076 161618
rect 498756 161340 499076 161382
rect 500228 161618 500548 162742
rect 500228 161382 500270 161618
rect 500506 161382 500548 161618
rect 500228 161340 500548 161382
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect 493052 156178 495212 156220
rect 493052 155942 493094 156178
rect 493330 155942 494934 156178
rect 495170 155942 495212 156178
rect 493052 155900 495212 155942
rect 497284 156178 499628 156220
rect 497284 155942 497326 156178
rect 497562 155942 499350 156178
rect 499586 155942 499628 156178
rect 497284 155900 499628 155942
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect 499308 152098 501652 152140
rect 499308 151862 499350 152098
rect 499586 151862 501374 152098
rect 501610 151862 501652 152098
rect 499308 151820 501652 151862
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect 497652 148018 499076 148060
rect 497652 147782 497694 148018
rect 497930 147782 498798 148018
rect 499034 147782 499076 148018
rect 497652 147740 499076 147782
rect 498020 147338 499628 147380
rect 498020 147102 498062 147338
rect 498298 147102 499350 147338
rect 499586 147102 499628 147338
rect 498020 147060 499628 147102
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect 486796 145298 487668 145340
rect 486796 145062 486838 145298
rect 487074 145062 487668 145298
rect 486796 145020 487668 145062
rect 487348 144660 487668 145020
rect 499860 145298 500180 145340
rect 499860 145062 499902 145298
rect 500138 145062 500180 145298
rect 499860 144660 500180 145062
rect 486796 144618 487668 144660
rect 486796 144382 486838 144618
rect 487074 144382 487668 144618
rect 486796 144340 487668 144382
rect 499676 144340 500180 144660
rect 497652 143938 499260 143980
rect 497652 143702 497694 143938
rect 497930 143702 498982 143938
rect 499218 143702 499260 143938
rect 497652 143660 499260 143702
rect 498020 143258 499260 143300
rect 498020 143022 498062 143258
rect 498298 143022 498982 143258
rect 499218 143022 499260 143258
rect 498020 142980 499260 143022
rect 499676 142620 499996 144340
rect 499676 142578 500180 142620
rect 499676 142342 499902 142578
rect 500138 142342 500180 142578
rect 499676 142300 500180 142342
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect 497652 137138 502204 137180
rect 497652 136902 497694 137138
rect 497930 136902 501926 137138
rect 502162 136902 502204 137138
rect 497652 136860 502204 136902
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect 499124 126938 500548 126980
rect 499124 126702 499166 126938
rect 499402 126702 500270 126938
rect 500506 126702 500548 126938
rect 499124 126660 500548 126702
rect 493052 123538 495028 123580
rect 493052 123302 493094 123538
rect 493330 123302 494750 123538
rect 494986 123302 495028 123538
rect 493052 123260 495028 123302
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect 493052 120138 495396 120180
rect 493052 119902 493094 120138
rect 493330 119902 495118 120138
rect 495354 119902 495396 120138
rect 493052 119860 495396 119902
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect 499676 116058 502204 116100
rect 499676 115822 499718 116058
rect 499954 115822 501926 116058
rect 502162 115822 502204 116058
rect 499676 115780 502204 115822
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect 495076 101820 496132 101956
rect 169396 101778 181676 101820
rect 169396 101542 169438 101778
rect 169674 101542 181676 101778
rect 169396 101500 181676 101542
rect 181356 101140 181676 101500
rect 186324 101500 205228 101820
rect 186324 101140 186644 101500
rect 181356 100820 186644 101140
rect 204908 100460 205228 101500
rect 215028 101140 215532 101820
rect 241340 101778 241660 101820
rect 241340 101542 241382 101778
rect 241618 101542 241660 101778
rect 241340 101140 241660 101542
rect 215028 100820 224916 101140
rect 241156 101098 241660 101140
rect 241156 100862 241198 101098
rect 241434 100862 241660 101098
rect 241156 100820 241660 100862
rect 253668 101140 254172 101820
rect 286972 101500 296860 101820
rect 286972 101140 287292 101500
rect 253668 100820 263556 101140
rect 273724 101098 287292 101140
rect 273724 100862 273766 101098
rect 274002 100862 287292 101098
rect 273724 100820 287292 100862
rect 215028 100460 215348 100820
rect 204908 100140 215348 100460
rect 224596 100460 224916 100820
rect 253668 100460 253988 100820
rect 224596 100418 232092 100460
rect 224596 100182 231814 100418
rect 232050 100182 232092 100418
rect 224596 100140 232092 100182
rect 250908 100418 253988 100460
rect 250908 100182 250950 100418
rect 251186 100182 253988 100418
rect 250908 100140 253988 100182
rect 263236 100460 263556 100820
rect 296540 100460 296860 101500
rect 311628 101500 316364 101820
rect 311628 100460 311948 101500
rect 316044 101140 316364 101500
rect 325612 101500 335500 101820
rect 325612 101140 325932 101500
rect 316044 100820 325932 101140
rect 263236 100418 270732 100460
rect 263236 100182 270454 100418
rect 270690 100182 270732 100418
rect 263236 100140 270732 100182
rect 296540 100140 311948 100460
rect 335180 100460 335500 101500
rect 364252 101500 374324 101820
rect 412276 101778 415724 101820
rect 412276 101542 412318 101778
rect 412554 101542 415724 101778
rect 412276 101500 415724 101542
rect 364252 101140 364572 101500
rect 351004 101098 364572 101140
rect 351004 100862 351046 101098
rect 351282 100862 364572 101098
rect 351004 100820 364572 100862
rect 374004 101140 374324 101500
rect 374004 101098 396036 101140
rect 374004 100862 395758 101098
rect 395994 100862 396036 101098
rect 374004 100820 396036 100862
rect 402708 101098 403948 101140
rect 402708 100862 402750 101098
rect 402986 100862 403670 101098
rect 403906 100862 403948 101098
rect 402708 100820 403948 100862
rect 415404 100460 415724 101500
rect 427732 101500 437620 101820
rect 427732 101140 428052 101500
rect 424788 100820 428052 101140
rect 437300 101140 437620 101500
rect 447052 101500 457124 101820
rect 447052 101140 447372 101500
rect 437300 100820 447372 101140
rect 456804 101140 457124 101500
rect 466372 101500 473500 101820
rect 495076 101778 504780 101820
rect 495076 101542 495118 101778
rect 495354 101636 504502 101778
rect 495354 101542 495396 101636
rect 495076 101500 495396 101542
rect 495812 101542 504502 101636
rect 504738 101542 504780 101778
rect 495812 101500 504780 101542
rect 466372 101140 466692 101500
rect 456804 100820 466692 101140
rect 473180 101140 473500 101500
rect 473180 101098 481780 101140
rect 473180 100862 481502 101098
rect 481738 100862 481780 101098
rect 473180 100820 481780 100862
rect 507036 101098 513612 101140
rect 507036 100862 507078 101098
rect 507314 100862 513334 101098
rect 513570 100862 513612 101098
rect 507036 100820 513612 100862
rect 424788 100460 425108 100820
rect 335180 100418 348012 100460
rect 335180 100182 347734 100418
rect 347970 100182 348012 100418
rect 335180 100140 348012 100182
rect 415404 100140 425108 100460
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect 466004 3858 496316 3900
rect 466004 3622 466046 3858
rect 466282 3622 496038 3858
rect 496274 3622 496316 3858
rect 466004 3580 496316 3622
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use Ibtida_top_dffram_cv  mprj
timestamp 1607406405
transform 1 0 82000 0 1 102000
box 0 0 420000 500000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
