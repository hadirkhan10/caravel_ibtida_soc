VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2818.490 89.660 2818.810 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2818.490 89.520 2899.310 89.660 ;
        RECT 2818.490 89.460 2818.810 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2818.520 89.460 2818.780 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 518.510 3022.075 518.790 3022.445 ;
        RECT 2818.510 3022.075 2818.790 3022.445 ;
        RECT 518.580 3010.000 518.720 3022.075 ;
        RECT 518.580 3009.340 518.930 3010.000 ;
        RECT 518.650 3006.000 518.930 3009.340 ;
        RECT 2818.580 89.750 2818.720 3022.075 ;
        RECT 2818.520 89.430 2818.780 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 518.510 3022.120 518.790 3022.400 ;
        RECT 2818.510 3022.120 2818.790 3022.400 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 518.485 3022.410 518.815 3022.425 ;
        RECT 2818.485 3022.410 2818.815 3022.425 ;
        RECT 518.485 3022.110 2818.815 3022.410 ;
        RECT 518.485 3022.095 518.815 3022.110 ;
        RECT 2818.485 3022.095 2818.815 3022.110 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2839.190 2429.200 2839.510 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2839.190 2429.060 2901.150 2429.200 ;
        RECT 2839.190 2429.000 2839.510 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2520.410 1531.600 2520.730 1531.660 ;
        RECT 2839.190 1531.600 2839.510 1531.660 ;
        RECT 2520.410 1531.460 2839.510 1531.600 ;
        RECT 2520.410 1531.400 2520.730 1531.460 ;
        RECT 2839.190 1531.400 2839.510 1531.460 ;
      LAYER via ;
        RECT 2839.220 2429.000 2839.480 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2520.440 1531.400 2520.700 1531.660 ;
        RECT 2839.220 1531.400 2839.480 1531.660 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2839.220 2428.970 2839.480 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2839.280 1531.690 2839.420 2428.970 ;
        RECT 2520.440 1531.370 2520.700 1531.690 ;
        RECT 2839.220 1531.370 2839.480 1531.690 ;
        RECT 2520.500 1526.445 2520.640 1531.370 ;
        RECT 2520.430 1526.075 2520.710 1526.445 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2520.430 1526.120 2520.710 1526.400 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2506.000 1526.410 2510.000 1526.560 ;
        RECT 2520.405 1526.410 2520.735 1526.425 ;
        RECT 2506.000 1526.110 2520.735 1526.410 ;
        RECT 2506.000 1525.960 2510.000 1526.110 ;
        RECT 2520.405 1526.095 2520.735 1526.110 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2037.410 3015.700 2037.730 3015.760 ;
        RECT 2536.050 3015.700 2536.370 3015.760 ;
        RECT 2037.410 3015.560 2536.370 3015.700 ;
        RECT 2037.410 3015.500 2037.730 3015.560 ;
        RECT 2536.050 3015.500 2536.370 3015.560 ;
        RECT 2536.050 2670.260 2536.370 2670.320 ;
        RECT 2900.830 2670.260 2901.150 2670.320 ;
        RECT 2536.050 2670.120 2901.150 2670.260 ;
        RECT 2536.050 2670.060 2536.370 2670.120 ;
        RECT 2900.830 2670.060 2901.150 2670.120 ;
      LAYER via ;
        RECT 2037.440 3015.500 2037.700 3015.760 ;
        RECT 2536.080 3015.500 2536.340 3015.760 ;
        RECT 2536.080 2670.060 2536.340 2670.320 ;
        RECT 2900.860 2670.060 2901.120 2670.320 ;
      LAYER met2 ;
        RECT 2037.440 3015.470 2037.700 3015.790 ;
        RECT 2536.080 3015.470 2536.340 3015.790 ;
        RECT 2037.500 3010.000 2037.640 3015.470 ;
        RECT 2037.500 3009.340 2037.850 3010.000 ;
        RECT 2037.570 3006.000 2037.850 3009.340 ;
        RECT 2536.140 2670.350 2536.280 3015.470 ;
        RECT 2536.080 2670.030 2536.340 2670.350 ;
        RECT 2900.860 2670.030 2901.120 2670.350 ;
        RECT 2900.920 2669.525 2901.060 2670.030 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2804.690 2898.400 2805.010 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2804.690 2898.260 2901.150 2898.400 ;
        RECT 2804.690 2898.200 2805.010 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2054.890 502.760 2055.210 502.820 ;
        RECT 2804.690 502.760 2805.010 502.820 ;
        RECT 2054.890 502.620 2805.010 502.760 ;
        RECT 2054.890 502.560 2055.210 502.620 ;
        RECT 2804.690 502.560 2805.010 502.620 ;
      LAYER via ;
        RECT 2804.720 2898.200 2804.980 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2054.920 502.560 2055.180 502.820 ;
        RECT 2804.720 502.560 2804.980 502.820 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2804.720 2898.170 2804.980 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2055.050 510.340 2055.330 514.000 ;
        RECT 2054.980 510.000 2055.330 510.340 ;
        RECT 2054.980 502.850 2055.120 510.000 ;
        RECT 2804.780 502.850 2804.920 2898.170 ;
        RECT 2054.920 502.530 2055.180 502.850 ;
        RECT 2804.720 502.530 2804.980 502.850 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 408.550 3133.000 408.870 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 408.550 3132.860 2901.150 3133.000 ;
        RECT 408.550 3132.800 408.870 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 408.580 3132.800 408.840 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 408.580 3132.770 408.840 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 408.640 1901.805 408.780 3132.770 ;
        RECT 408.570 1901.435 408.850 1901.805 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 408.570 1901.480 408.850 1901.760 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 408.545 1901.770 408.875 1901.785 ;
        RECT 410.000 1901.770 414.000 1901.920 ;
        RECT 408.545 1901.470 414.000 1901.770 ;
        RECT 408.545 1901.455 408.875 1901.470 ;
        RECT 410.000 1901.320 414.000 1901.470 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.470 3369.980 869.790 3370.040 ;
        RECT 891.550 3369.980 891.870 3370.040 ;
        RECT 869.470 3369.840 891.870 3369.980 ;
        RECT 869.470 3369.780 869.790 3369.840 ;
        RECT 891.550 3369.780 891.870 3369.840 ;
        RECT 772.870 3368.960 773.190 3369.020 ;
        RECT 811.050 3368.960 811.370 3369.020 ;
        RECT 772.870 3368.820 811.370 3368.960 ;
        RECT 772.870 3368.760 773.190 3368.820 ;
        RECT 811.050 3368.760 811.370 3368.820 ;
      LAYER via ;
        RECT 869.500 3369.780 869.760 3370.040 ;
        RECT 891.580 3369.780 891.840 3370.040 ;
        RECT 772.900 3368.760 773.160 3369.020 ;
        RECT 811.080 3368.760 811.340 3369.020 ;
      LAYER met2 ;
        RECT 941.710 3370.235 941.990 3370.605 ;
        RECT 869.500 3369.925 869.760 3370.070 ;
        RECT 869.490 3369.555 869.770 3369.925 ;
        RECT 891.580 3369.750 891.840 3370.070 ;
        RECT 891.640 3369.245 891.780 3369.750 ;
        RECT 941.780 3369.245 941.920 3370.235 ;
        RECT 772.890 3368.875 773.170 3369.245 ;
        RECT 772.900 3368.730 773.160 3368.875 ;
        RECT 811.080 3368.730 811.340 3369.050 ;
        RECT 834.530 3368.875 834.810 3369.245 ;
        RECT 891.570 3368.875 891.850 3369.245 ;
        RECT 941.710 3368.875 941.990 3369.245 ;
        RECT 811.140 3367.885 811.280 3368.730 ;
        RECT 834.600 3367.885 834.740 3368.875 ;
        RECT 811.070 3367.515 811.350 3367.885 ;
        RECT 834.530 3367.515 834.810 3367.885 ;
      LAYER via2 ;
        RECT 941.710 3370.280 941.990 3370.560 ;
        RECT 869.490 3369.600 869.770 3369.880 ;
        RECT 772.890 3368.920 773.170 3369.200 ;
        RECT 834.530 3368.920 834.810 3369.200 ;
        RECT 891.570 3368.920 891.850 3369.200 ;
        RECT 941.710 3368.920 941.990 3369.200 ;
        RECT 811.070 3367.560 811.350 3367.840 ;
        RECT 834.530 3367.560 834.810 3367.840 ;
      LAYER met3 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2916.710 3372.990 2924.800 3373.290 ;
        RECT 917.510 3370.570 917.890 3370.580 ;
        RECT 941.685 3370.570 942.015 3370.585 ;
        RECT 917.510 3370.270 942.015 3370.570 ;
        RECT 917.510 3370.260 917.890 3370.270 ;
        RECT 941.685 3370.255 942.015 3370.270 ;
        RECT 869.465 3369.890 869.795 3369.905 ;
        RECT 836.590 3369.590 869.795 3369.890 ;
        RECT 772.865 3369.210 773.195 3369.225 ;
        RECT 399.590 3368.910 421.050 3369.210 ;
        RECT 399.590 3368.530 399.890 3368.910 ;
        RECT 351.750 3368.230 399.890 3368.530 ;
        RECT 420.750 3368.530 421.050 3368.910 ;
        RECT 469.510 3368.910 517.650 3369.210 ;
        RECT 420.750 3368.230 468.890 3368.530 ;
        RECT 350.790 3367.850 351.170 3367.860 ;
        RECT 351.750 3367.850 352.050 3368.230 ;
        RECT 350.790 3367.550 352.050 3367.850 ;
        RECT 468.590 3367.850 468.890 3368.230 ;
        RECT 469.510 3367.850 469.810 3368.910 ;
        RECT 517.350 3368.530 517.650 3368.910 ;
        RECT 566.110 3368.910 614.250 3369.210 ;
        RECT 517.350 3368.230 565.490 3368.530 ;
        RECT 468.590 3367.550 469.810 3367.850 ;
        RECT 565.190 3367.850 565.490 3368.230 ;
        RECT 566.110 3367.850 566.410 3368.910 ;
        RECT 613.950 3368.530 614.250 3368.910 ;
        RECT 662.710 3368.910 710.850 3369.210 ;
        RECT 613.950 3368.230 662.090 3368.530 ;
        RECT 565.190 3367.550 566.410 3367.850 ;
        RECT 661.790 3367.850 662.090 3368.230 ;
        RECT 662.710 3367.850 663.010 3368.910 ;
        RECT 710.550 3368.530 710.850 3368.910 ;
        RECT 759.310 3368.910 773.195 3369.210 ;
        RECT 710.550 3368.230 758.690 3368.530 ;
        RECT 661.790 3367.550 663.010 3367.850 ;
        RECT 758.390 3367.850 758.690 3368.230 ;
        RECT 759.310 3367.850 759.610 3368.910 ;
        RECT 772.865 3368.895 773.195 3368.910 ;
        RECT 834.505 3369.210 834.835 3369.225 ;
        RECT 836.590 3369.210 836.890 3369.590 ;
        RECT 869.465 3369.575 869.795 3369.590 ;
        RECT 834.505 3368.910 836.890 3369.210 ;
        RECT 891.545 3369.210 891.875 3369.225 ;
        RECT 917.510 3369.210 917.890 3369.220 ;
        RECT 891.545 3368.910 917.890 3369.210 ;
        RECT 834.505 3368.895 834.835 3368.910 ;
        RECT 891.545 3368.895 891.875 3368.910 ;
        RECT 917.510 3368.900 917.890 3368.910 ;
        RECT 941.685 3369.210 942.015 3369.225 ;
        RECT 941.685 3368.910 1000.650 3369.210 ;
        RECT 941.685 3368.895 942.015 3368.910 ;
        RECT 1000.350 3368.530 1000.650 3368.910 ;
        RECT 1049.110 3368.910 1097.250 3369.210 ;
        RECT 1000.350 3368.230 1048.490 3368.530 ;
        RECT 758.390 3367.550 759.610 3367.850 ;
        RECT 811.045 3367.850 811.375 3367.865 ;
        RECT 834.505 3367.850 834.835 3367.865 ;
        RECT 811.045 3367.550 834.835 3367.850 ;
        RECT 1048.190 3367.850 1048.490 3368.230 ;
        RECT 1049.110 3367.850 1049.410 3368.910 ;
        RECT 1096.950 3368.530 1097.250 3368.910 ;
        RECT 1145.710 3368.910 1193.850 3369.210 ;
        RECT 1096.950 3368.230 1145.090 3368.530 ;
        RECT 1048.190 3367.550 1049.410 3367.850 ;
        RECT 1144.790 3367.850 1145.090 3368.230 ;
        RECT 1145.710 3367.850 1146.010 3368.910 ;
        RECT 1193.550 3368.530 1193.850 3368.910 ;
        RECT 1242.310 3368.910 1290.450 3369.210 ;
        RECT 1193.550 3368.230 1241.690 3368.530 ;
        RECT 1144.790 3367.550 1146.010 3367.850 ;
        RECT 1241.390 3367.850 1241.690 3368.230 ;
        RECT 1242.310 3367.850 1242.610 3368.910 ;
        RECT 1290.150 3368.530 1290.450 3368.910 ;
        RECT 1338.910 3368.910 1387.050 3369.210 ;
        RECT 1290.150 3368.230 1338.290 3368.530 ;
        RECT 1241.390 3367.550 1242.610 3367.850 ;
        RECT 1337.990 3367.850 1338.290 3368.230 ;
        RECT 1338.910 3367.850 1339.210 3368.910 ;
        RECT 1386.750 3368.530 1387.050 3368.910 ;
        RECT 1435.510 3368.910 1483.650 3369.210 ;
        RECT 1386.750 3368.230 1434.890 3368.530 ;
        RECT 1337.990 3367.550 1339.210 3367.850 ;
        RECT 1434.590 3367.850 1434.890 3368.230 ;
        RECT 1435.510 3367.850 1435.810 3368.910 ;
        RECT 1483.350 3368.530 1483.650 3368.910 ;
        RECT 1532.110 3368.910 1580.250 3369.210 ;
        RECT 1483.350 3368.230 1531.490 3368.530 ;
        RECT 1434.590 3367.550 1435.810 3367.850 ;
        RECT 1531.190 3367.850 1531.490 3368.230 ;
        RECT 1532.110 3367.850 1532.410 3368.910 ;
        RECT 1579.950 3368.530 1580.250 3368.910 ;
        RECT 1628.710 3368.910 1676.850 3369.210 ;
        RECT 1579.950 3368.230 1628.090 3368.530 ;
        RECT 1531.190 3367.550 1532.410 3367.850 ;
        RECT 1627.790 3367.850 1628.090 3368.230 ;
        RECT 1628.710 3367.850 1629.010 3368.910 ;
        RECT 1676.550 3368.530 1676.850 3368.910 ;
        RECT 1725.310 3368.910 1773.450 3369.210 ;
        RECT 1676.550 3368.230 1724.690 3368.530 ;
        RECT 1627.790 3367.550 1629.010 3367.850 ;
        RECT 1724.390 3367.850 1724.690 3368.230 ;
        RECT 1725.310 3367.850 1725.610 3368.910 ;
        RECT 1773.150 3368.530 1773.450 3368.910 ;
        RECT 1821.910 3368.910 1870.050 3369.210 ;
        RECT 1773.150 3368.230 1821.290 3368.530 ;
        RECT 1724.390 3367.550 1725.610 3367.850 ;
        RECT 1820.990 3367.850 1821.290 3368.230 ;
        RECT 1821.910 3367.850 1822.210 3368.910 ;
        RECT 1869.750 3368.530 1870.050 3368.910 ;
        RECT 1918.510 3368.910 1966.650 3369.210 ;
        RECT 1869.750 3368.230 1917.890 3368.530 ;
        RECT 1820.990 3367.550 1822.210 3367.850 ;
        RECT 1917.590 3367.850 1917.890 3368.230 ;
        RECT 1918.510 3367.850 1918.810 3368.910 ;
        RECT 1966.350 3368.530 1966.650 3368.910 ;
        RECT 2015.110 3368.910 2063.250 3369.210 ;
        RECT 1966.350 3368.230 2014.490 3368.530 ;
        RECT 1917.590 3367.550 1918.810 3367.850 ;
        RECT 2014.190 3367.850 2014.490 3368.230 ;
        RECT 2015.110 3367.850 2015.410 3368.910 ;
        RECT 2062.950 3368.530 2063.250 3368.910 ;
        RECT 2159.550 3368.910 2207.690 3369.210 ;
        RECT 2062.950 3368.230 2111.090 3368.530 ;
        RECT 2014.190 3367.550 2015.410 3367.850 ;
        RECT 2110.790 3367.850 2111.090 3368.230 ;
        RECT 2159.550 3367.850 2159.850 3368.910 ;
        RECT 2110.790 3367.550 2159.850 3367.850 ;
        RECT 2207.390 3367.850 2207.690 3368.910 ;
        RECT 2208.310 3368.910 2256.450 3369.210 ;
        RECT 2208.310 3367.850 2208.610 3368.910 ;
        RECT 2256.150 3368.530 2256.450 3368.910 ;
        RECT 2304.910 3368.910 2353.050 3369.210 ;
        RECT 2256.150 3368.230 2304.290 3368.530 ;
        RECT 2207.390 3367.550 2208.610 3367.850 ;
        RECT 2303.990 3367.850 2304.290 3368.230 ;
        RECT 2304.910 3367.850 2305.210 3368.910 ;
        RECT 2352.750 3368.530 2353.050 3368.910 ;
        RECT 2401.510 3368.910 2449.650 3369.210 ;
        RECT 2352.750 3368.230 2400.890 3368.530 ;
        RECT 2303.990 3367.550 2305.210 3367.850 ;
        RECT 2400.590 3367.850 2400.890 3368.230 ;
        RECT 2401.510 3367.850 2401.810 3368.910 ;
        RECT 2449.350 3368.530 2449.650 3368.910 ;
        RECT 2498.110 3368.910 2546.250 3369.210 ;
        RECT 2449.350 3368.230 2497.490 3368.530 ;
        RECT 2400.590 3367.550 2401.810 3367.850 ;
        RECT 2497.190 3367.850 2497.490 3368.230 ;
        RECT 2498.110 3367.850 2498.410 3368.910 ;
        RECT 2545.950 3368.530 2546.250 3368.910 ;
        RECT 2594.710 3368.910 2642.850 3369.210 ;
        RECT 2545.950 3368.230 2594.090 3368.530 ;
        RECT 2497.190 3367.550 2498.410 3367.850 ;
        RECT 2593.790 3367.850 2594.090 3368.230 ;
        RECT 2594.710 3367.850 2595.010 3368.910 ;
        RECT 2642.550 3368.530 2642.850 3368.910 ;
        RECT 2691.310 3368.910 2739.450 3369.210 ;
        RECT 2642.550 3368.230 2690.690 3368.530 ;
        RECT 2593.790 3367.550 2595.010 3367.850 ;
        RECT 2690.390 3367.850 2690.690 3368.230 ;
        RECT 2691.310 3367.850 2691.610 3368.910 ;
        RECT 2739.150 3368.530 2739.450 3368.910 ;
        RECT 2787.910 3368.910 2836.050 3369.210 ;
        RECT 2739.150 3368.230 2787.290 3368.530 ;
        RECT 2690.390 3367.550 2691.610 3367.850 ;
        RECT 2786.990 3367.850 2787.290 3368.230 ;
        RECT 2787.910 3367.850 2788.210 3368.910 ;
        RECT 2835.750 3368.530 2836.050 3368.910 ;
        RECT 2916.710 3368.530 2917.010 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2835.750 3368.230 2883.890 3368.530 ;
        RECT 2786.990 3367.550 2788.210 3367.850 ;
        RECT 2883.590 3367.850 2883.890 3368.230 ;
        RECT 2884.510 3368.230 2917.010 3368.530 ;
        RECT 2884.510 3367.850 2884.810 3368.230 ;
        RECT 2883.590 3367.550 2884.810 3367.850 ;
        RECT 350.790 3367.540 351.170 3367.550 ;
        RECT 811.045 3367.535 811.375 3367.550 ;
        RECT 834.505 3367.535 834.835 3367.550 ;
        RECT 350.790 1027.970 351.170 1027.980 ;
        RECT 350.790 1027.670 410.930 1027.970 ;
        RECT 350.790 1027.660 351.170 1027.670 ;
        RECT 410.630 1024.720 410.930 1027.670 ;
        RECT 410.000 1024.120 414.000 1024.720 ;
      LAYER via3 ;
        RECT 917.540 3370.260 917.860 3370.580 ;
        RECT 350.820 3367.540 351.140 3367.860 ;
        RECT 917.540 3368.900 917.860 3369.220 ;
        RECT 350.820 1027.660 351.140 1027.980 ;
      LAYER met4 ;
        RECT 917.535 3370.255 917.865 3370.585 ;
        RECT 917.550 3369.225 917.850 3370.255 ;
        RECT 917.535 3368.895 917.865 3369.225 ;
        RECT 350.815 3367.535 351.145 3367.865 ;
        RECT 350.830 1027.985 351.130 3367.535 ;
        RECT 350.815 1027.655 351.145 1027.985 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2717.750 3501.560 2718.070 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2717.750 3501.420 2798.570 3501.560 ;
        RECT 2717.750 3501.360 2718.070 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 2714.990 3498.500 2715.310 3498.560 ;
        RECT 2717.750 3498.500 2718.070 3498.560 ;
        RECT 2714.990 3498.360 2718.070 3498.500 ;
        RECT 2714.990 3498.300 2715.310 3498.360 ;
        RECT 2717.750 3498.300 2718.070 3498.360 ;
        RECT 641.770 3053.100 642.090 3053.160 ;
        RECT 2714.990 3053.100 2715.310 3053.160 ;
        RECT 641.770 3052.960 2715.310 3053.100 ;
        RECT 641.770 3052.900 642.090 3052.960 ;
        RECT 2714.990 3052.900 2715.310 3052.960 ;
      LAYER via ;
        RECT 2717.780 3501.360 2718.040 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 2715.020 3498.300 2715.280 3498.560 ;
        RECT 2717.780 3498.300 2718.040 3498.560 ;
        RECT 641.800 3052.900 642.060 3053.160 ;
        RECT 2715.020 3052.900 2715.280 3053.160 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2717.780 3501.330 2718.040 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 2717.840 3498.590 2717.980 3501.330 ;
        RECT 2715.020 3498.270 2715.280 3498.590 ;
        RECT 2717.780 3498.270 2718.040 3498.590 ;
        RECT 2715.080 3053.190 2715.220 3498.270 ;
        RECT 641.800 3052.870 642.060 3053.190 ;
        RECT 2715.020 3052.870 2715.280 3053.190 ;
        RECT 641.860 3010.000 642.000 3052.870 ;
        RECT 641.860 3009.340 642.210 3010.000 ;
        RECT 641.930 3006.000 642.210 3009.340 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.845 2474.180 3517.600 ;
        RECT 2473.970 3501.475 2474.250 3501.845 ;
        RECT 857.210 510.340 857.490 514.000 ;
        RECT 857.140 510.000 857.490 510.340 ;
        RECT 857.140 503.725 857.280 510.000 ;
        RECT 857.070 503.355 857.350 503.725 ;
      LAYER via2 ;
        RECT 2473.970 3501.520 2474.250 3501.800 ;
        RECT 857.070 503.400 857.350 503.680 ;
      LAYER met3 ;
        RECT 2431.830 3501.810 2432.210 3501.820 ;
        RECT 2473.945 3501.810 2474.275 3501.825 ;
        RECT 2431.830 3501.510 2474.275 3501.810 ;
        RECT 2431.830 3501.500 2432.210 3501.510 ;
        RECT 2473.945 3501.495 2474.275 3501.510 ;
        RECT 857.045 503.690 857.375 503.705 ;
        RECT 2431.830 503.690 2432.210 503.700 ;
        RECT 857.045 503.390 2432.210 503.690 ;
        RECT 857.045 503.375 857.375 503.390 ;
        RECT 2431.830 503.380 2432.210 503.390 ;
      LAYER via3 ;
        RECT 2431.860 3501.500 2432.180 3501.820 ;
        RECT 2431.860 503.380 2432.180 503.700 ;
      LAYER met4 ;
        RECT 2431.855 3501.495 2432.185 3501.825 ;
        RECT 2431.870 503.705 2432.170 3501.495 ;
        RECT 2431.855 503.375 2432.185 503.705 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.970 3464.160 2146.290 3464.220 ;
        RECT 2149.650 3464.160 2149.970 3464.220 ;
        RECT 2145.970 3464.020 2149.970 3464.160 ;
        RECT 2145.970 3463.960 2146.290 3464.020 ;
        RECT 2149.650 3463.960 2149.970 3464.020 ;
        RECT 2145.970 3367.260 2146.290 3367.320 ;
        RECT 2147.350 3367.260 2147.670 3367.320 ;
        RECT 2145.970 3367.120 2147.670 3367.260 ;
        RECT 2145.970 3367.060 2146.290 3367.120 ;
        RECT 2147.350 3367.060 2147.670 3367.120 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2145.970 3056.840 2146.290 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2145.970 3056.700 2147.670 3056.840 ;
        RECT 2145.970 3056.640 2146.290 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 1642.730 3032.360 1643.050 3032.420 ;
        RECT 2145.970 3032.360 2146.290 3032.420 ;
        RECT 1642.730 3032.220 2146.290 3032.360 ;
        RECT 1642.730 3032.160 1643.050 3032.220 ;
        RECT 2145.970 3032.160 2146.290 3032.220 ;
      LAYER via ;
        RECT 2146.000 3463.960 2146.260 3464.220 ;
        RECT 2149.680 3463.960 2149.940 3464.220 ;
        RECT 2146.000 3367.060 2146.260 3367.320 ;
        RECT 2147.380 3367.060 2147.640 3367.320 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.000 3056.640 2146.260 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 1642.760 3032.160 1643.020 3032.420 ;
        RECT 2146.000 3032.160 2146.260 3032.420 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2149.280 3517.230 2149.880 3517.370 ;
        RECT 2149.740 3464.250 2149.880 3517.230 ;
        RECT 2146.000 3463.930 2146.260 3464.250 ;
        RECT 2149.680 3463.930 2149.940 3464.250 ;
        RECT 2146.060 3367.350 2146.200 3463.930 ;
        RECT 2146.000 3367.030 2146.260 3367.350 ;
        RECT 2147.380 3367.030 2147.640 3367.350 ;
        RECT 2147.440 3236.450 2147.580 3367.030 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.000 3056.610 2146.260 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.060 3032.450 2146.200 3056.610 ;
        RECT 1642.760 3032.130 1643.020 3032.450 ;
        RECT 2146.000 3032.130 2146.260 3032.450 ;
        RECT 1642.820 3010.000 1642.960 3032.130 ;
        RECT 1642.820 3009.340 1643.170 3010.000 ;
        RECT 1642.890 3006.000 1643.170 3009.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3502.240 1825.210 3502.300 ;
        RECT 2549.850 3502.240 2550.170 3502.300 ;
        RECT 1824.890 3502.100 2550.170 3502.240 ;
        RECT 1824.890 3502.040 1825.210 3502.100 ;
        RECT 2549.850 3502.040 2550.170 3502.100 ;
        RECT 2376.890 501.400 2377.210 501.460 ;
        RECT 2549.850 501.400 2550.170 501.460 ;
        RECT 2376.890 501.260 2550.170 501.400 ;
        RECT 2376.890 501.200 2377.210 501.260 ;
        RECT 2549.850 501.200 2550.170 501.260 ;
      LAYER via ;
        RECT 1824.920 3502.040 1825.180 3502.300 ;
        RECT 2549.880 3502.040 2550.140 3502.300 ;
        RECT 2376.920 501.200 2377.180 501.460 ;
        RECT 2549.880 501.200 2550.140 501.460 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.330 1825.120 3517.600 ;
        RECT 1824.920 3502.010 1825.180 3502.330 ;
        RECT 2549.880 3502.010 2550.140 3502.330 ;
        RECT 2377.050 510.340 2377.330 514.000 ;
        RECT 2376.980 510.000 2377.330 510.340 ;
        RECT 2376.980 501.490 2377.120 510.000 ;
        RECT 2549.940 501.490 2550.080 3502.010 ;
        RECT 2376.920 501.170 2377.180 501.490 ;
        RECT 2549.880 501.170 2550.140 501.490 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 3494.760 1297.130 3494.820 ;
        RECT 1500.590 3494.760 1500.910 3494.820 ;
        RECT 1296.810 3494.620 1500.910 3494.760 ;
        RECT 1296.810 3494.560 1297.130 3494.620 ;
        RECT 1500.590 3494.560 1500.910 3494.620 ;
      LAYER via ;
        RECT 1296.840 3494.560 1297.100 3494.820 ;
        RECT 1500.620 3494.560 1500.880 3494.820 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3494.850 1500.820 3517.600 ;
        RECT 1296.840 3494.530 1297.100 3494.850 ;
        RECT 1500.620 3494.530 1500.880 3494.850 ;
        RECT 1296.900 3010.000 1297.040 3494.530 ;
        RECT 1296.900 3009.340 1297.250 3010.000 ;
        RECT 1296.970 3006.000 1297.250 3009.340 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1159.300 2520.730 1159.360 ;
        RECT 2597.690 1159.300 2598.010 1159.360 ;
        RECT 2520.410 1159.160 2598.010 1159.300 ;
        RECT 2520.410 1159.100 2520.730 1159.160 ;
        RECT 2597.690 1159.100 2598.010 1159.160 ;
        RECT 2597.690 324.260 2598.010 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2597.690 324.120 2899.310 324.260 ;
        RECT 2597.690 324.060 2598.010 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2520.440 1159.100 2520.700 1159.360 ;
        RECT 2597.720 1159.100 2597.980 1159.360 ;
        RECT 2597.720 324.060 2597.980 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2520.430 1160.235 2520.710 1160.605 ;
        RECT 2520.500 1159.390 2520.640 1160.235 ;
        RECT 2520.440 1159.070 2520.700 1159.390 ;
        RECT 2597.720 1159.070 2597.980 1159.390 ;
        RECT 2597.780 324.350 2597.920 1159.070 ;
        RECT 2597.720 324.030 2597.980 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2520.430 1160.280 2520.710 1160.560 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2506.000 1160.570 2510.000 1160.720 ;
        RECT 2520.405 1160.570 2520.735 1160.585 ;
        RECT 2506.000 1160.270 2520.735 1160.570 ;
        RECT 2506.000 1160.120 2510.000 1160.270 ;
        RECT 2520.405 1160.255 2520.735 1160.270 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 379.110 3502.580 379.430 3502.640 ;
        RECT 1175.830 3502.580 1176.150 3502.640 ;
        RECT 379.110 3502.440 1176.150 3502.580 ;
        RECT 379.110 3502.380 379.430 3502.440 ;
        RECT 1175.830 3502.380 1176.150 3502.440 ;
        RECT 379.110 501.060 379.430 501.120 ;
        RECT 560.810 501.060 561.130 501.120 ;
        RECT 379.110 500.920 561.130 501.060 ;
        RECT 379.110 500.860 379.430 500.920 ;
        RECT 560.810 500.860 561.130 500.920 ;
      LAYER via ;
        RECT 379.140 3502.380 379.400 3502.640 ;
        RECT 1175.860 3502.380 1176.120 3502.640 ;
        RECT 379.140 500.860 379.400 501.120 ;
        RECT 560.840 500.860 561.100 501.120 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3502.670 1176.060 3517.600 ;
        RECT 379.140 3502.350 379.400 3502.670 ;
        RECT 1175.860 3502.350 1176.120 3502.670 ;
        RECT 379.200 501.150 379.340 3502.350 ;
        RECT 560.970 510.340 561.250 514.000 ;
        RECT 560.900 510.000 561.250 510.340 ;
        RECT 560.900 501.150 561.040 510.000 ;
        RECT 379.140 500.830 379.400 501.150 ;
        RECT 560.840 500.830 561.100 501.150 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 850.685 3332.765 850.855 3415.555 ;
      LAYER mcon ;
        RECT 850.685 3415.385 850.855 3415.555 ;
      LAYER met1 ;
        RECT 849.690 3477.420 850.010 3477.480 ;
        RECT 851.530 3477.420 851.850 3477.480 ;
        RECT 849.690 3477.280 851.850 3477.420 ;
        RECT 849.690 3477.220 850.010 3477.280 ;
        RECT 851.530 3477.220 851.850 3477.280 ;
        RECT 849.690 3439.680 850.010 3439.740 ;
        RECT 850.610 3439.680 850.930 3439.740 ;
        RECT 849.690 3439.540 850.930 3439.680 ;
        RECT 849.690 3439.480 850.010 3439.540 ;
        RECT 850.610 3439.480 850.930 3439.540 ;
        RECT 848.770 3415.540 849.090 3415.600 ;
        RECT 850.625 3415.540 850.915 3415.585 ;
        RECT 848.770 3415.400 850.915 3415.540 ;
        RECT 848.770 3415.340 849.090 3415.400 ;
        RECT 850.625 3415.355 850.915 3415.400 ;
        RECT 850.625 3332.920 850.915 3332.965 ;
        RECT 851.070 3332.920 851.390 3332.980 ;
        RECT 850.625 3332.780 851.390 3332.920 ;
        RECT 850.625 3332.735 850.915 3332.780 ;
        RECT 851.070 3332.720 851.390 3332.780 ;
        RECT 849.690 3236.360 850.010 3236.420 ;
        RECT 850.150 3236.360 850.470 3236.420 ;
        RECT 849.690 3236.220 850.470 3236.360 ;
        RECT 849.690 3236.160 850.010 3236.220 ;
        RECT 850.150 3236.160 850.470 3236.220 ;
        RECT 849.690 3202.020 850.010 3202.080 ;
        RECT 850.150 3202.020 850.470 3202.080 ;
        RECT 849.690 3201.880 850.470 3202.020 ;
        RECT 849.690 3201.820 850.010 3201.880 ;
        RECT 850.150 3201.820 850.470 3201.880 ;
        RECT 849.230 3153.400 849.550 3153.460 ;
        RECT 850.150 3153.400 850.470 3153.460 ;
        RECT 849.230 3153.260 850.470 3153.400 ;
        RECT 849.230 3153.200 849.550 3153.260 ;
        RECT 850.150 3153.200 850.470 3153.260 ;
        RECT 848.770 3056.840 849.090 3056.900 ;
        RECT 850.150 3056.840 850.470 3056.900 ;
        RECT 848.770 3056.700 850.470 3056.840 ;
        RECT 848.770 3056.640 849.090 3056.700 ;
        RECT 850.150 3056.640 850.470 3056.700 ;
        RECT 408.090 3039.500 408.410 3039.560 ;
        RECT 848.770 3039.500 849.090 3039.560 ;
        RECT 408.090 3039.360 849.090 3039.500 ;
        RECT 408.090 3039.300 408.410 3039.360 ;
        RECT 848.770 3039.300 849.090 3039.360 ;
      LAYER via ;
        RECT 849.720 3477.220 849.980 3477.480 ;
        RECT 851.560 3477.220 851.820 3477.480 ;
        RECT 849.720 3439.480 849.980 3439.740 ;
        RECT 850.640 3439.480 850.900 3439.740 ;
        RECT 848.800 3415.340 849.060 3415.600 ;
        RECT 851.100 3332.720 851.360 3332.980 ;
        RECT 849.720 3236.160 849.980 3236.420 ;
        RECT 850.180 3236.160 850.440 3236.420 ;
        RECT 849.720 3201.820 849.980 3202.080 ;
        RECT 850.180 3201.820 850.440 3202.080 ;
        RECT 849.260 3153.200 849.520 3153.460 ;
        RECT 850.180 3153.200 850.440 3153.460 ;
        RECT 848.800 3056.640 849.060 3056.900 ;
        RECT 850.180 3056.640 850.440 3056.900 ;
        RECT 408.120 3039.300 408.380 3039.560 ;
        RECT 848.800 3039.300 849.060 3039.560 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3477.510 851.760 3517.600 ;
        RECT 849.720 3477.190 849.980 3477.510 ;
        RECT 851.560 3477.190 851.820 3477.510 ;
        RECT 849.780 3439.770 849.920 3477.190 ;
        RECT 849.720 3439.450 849.980 3439.770 ;
        RECT 850.640 3439.450 850.900 3439.770 ;
        RECT 850.700 3416.165 850.840 3439.450 ;
        RECT 848.790 3415.795 849.070 3416.165 ;
        RECT 850.630 3415.795 850.910 3416.165 ;
        RECT 848.860 3415.630 849.000 3415.795 ;
        RECT 848.800 3415.310 849.060 3415.630 ;
        RECT 851.100 3332.690 851.360 3333.010 ;
        RECT 851.160 3298.410 851.300 3332.690 ;
        RECT 850.240 3298.270 851.300 3298.410 ;
        RECT 850.240 3236.450 850.380 3298.270 ;
        RECT 849.720 3236.130 849.980 3236.450 ;
        RECT 850.180 3236.130 850.440 3236.450 ;
        RECT 849.780 3202.110 849.920 3236.130 ;
        RECT 849.720 3201.790 849.980 3202.110 ;
        RECT 850.180 3201.790 850.440 3202.110 ;
        RECT 850.240 3153.490 850.380 3201.790 ;
        RECT 849.260 3153.170 849.520 3153.490 ;
        RECT 850.180 3153.170 850.440 3153.490 ;
        RECT 849.320 3152.890 849.460 3153.170 ;
        RECT 849.320 3152.750 849.920 3152.890 ;
        RECT 849.780 3105.290 849.920 3152.750 ;
        RECT 849.780 3105.150 850.380 3105.290 ;
        RECT 850.240 3056.930 850.380 3105.150 ;
        RECT 848.800 3056.610 849.060 3056.930 ;
        RECT 850.180 3056.610 850.440 3056.930 ;
        RECT 848.860 3039.590 849.000 3056.610 ;
        RECT 408.120 3039.270 408.380 3039.590 ;
        RECT 848.800 3039.270 849.060 3039.590 ;
        RECT 408.180 1572.685 408.320 3039.270 ;
        RECT 408.110 1572.315 408.390 1572.685 ;
      LAYER via2 ;
        RECT 848.790 3415.840 849.070 3416.120 ;
        RECT 850.630 3415.840 850.910 3416.120 ;
        RECT 408.110 1572.360 408.390 1572.640 ;
      LAYER met3 ;
        RECT 848.765 3416.130 849.095 3416.145 ;
        RECT 850.605 3416.130 850.935 3416.145 ;
        RECT 848.765 3415.830 850.935 3416.130 ;
        RECT 848.765 3415.815 849.095 3415.830 ;
        RECT 850.605 3415.815 850.935 3415.830 ;
        RECT 408.085 1572.650 408.415 1572.665 ;
        RECT 410.000 1572.650 414.000 1572.800 ;
        RECT 408.085 1572.350 414.000 1572.650 ;
        RECT 408.085 1572.335 408.415 1572.350 ;
        RECT 410.000 1572.200 414.000 1572.350 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.470 3498.500 524.790 3498.560 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 524.470 3498.360 527.550 3498.500 ;
        RECT 524.470 3498.300 524.790 3498.360 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 357.490 3011.960 357.810 3012.020 ;
        RECT 524.010 3011.960 524.330 3012.020 ;
        RECT 357.490 3011.820 524.330 3011.960 ;
        RECT 357.490 3011.760 357.810 3011.820 ;
        RECT 524.010 3011.760 524.330 3011.820 ;
        RECT 357.490 501.740 357.810 501.800 ;
        RECT 820.250 501.740 820.570 501.800 ;
        RECT 357.490 501.600 820.570 501.740 ;
        RECT 357.490 501.540 357.810 501.600 ;
        RECT 820.250 501.540 820.570 501.600 ;
      LAYER via ;
        RECT 524.500 3498.300 524.760 3498.560 ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 357.520 3011.760 357.780 3012.020 ;
        RECT 524.040 3011.760 524.300 3012.020 ;
        RECT 357.520 501.540 357.780 501.800 ;
        RECT 820.280 501.540 820.540 501.800 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 524.500 3498.270 524.760 3498.590 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 524.560 3012.130 524.700 3498.270 ;
        RECT 524.100 3012.050 524.700 3012.130 ;
        RECT 357.520 3011.730 357.780 3012.050 ;
        RECT 524.040 3011.990 524.700 3012.050 ;
        RECT 524.040 3011.730 524.300 3011.990 ;
        RECT 357.580 501.830 357.720 3011.730 ;
        RECT 820.410 510.340 820.690 514.000 ;
        RECT 820.340 510.000 820.690 510.340 ;
        RECT 820.340 501.830 820.480 510.000 ;
        RECT 357.520 501.510 357.780 501.830 ;
        RECT 820.280 501.510 820.540 501.830 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3498.500 202.790 3498.560 ;
        RECT 217.190 3498.500 217.510 3498.560 ;
        RECT 202.470 3498.360 217.510 3498.500 ;
        RECT 202.470 3498.300 202.790 3498.360 ;
        RECT 217.190 3498.300 217.510 3498.360 ;
        RECT 217.190 3080.640 217.510 3080.700 ;
        RECT 1994.170 3080.640 1994.490 3080.700 ;
        RECT 217.190 3080.500 1994.490 3080.640 ;
        RECT 217.190 3080.440 217.510 3080.500 ;
        RECT 1994.170 3080.440 1994.490 3080.500 ;
      LAYER via ;
        RECT 202.500 3498.300 202.760 3498.560 ;
        RECT 217.220 3498.300 217.480 3498.560 ;
        RECT 217.220 3080.440 217.480 3080.700 ;
        RECT 1994.200 3080.440 1994.460 3080.700 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3498.590 202.700 3517.600 ;
        RECT 202.500 3498.270 202.760 3498.590 ;
        RECT 217.220 3498.270 217.480 3498.590 ;
        RECT 217.280 3080.730 217.420 3498.270 ;
        RECT 217.220 3080.410 217.480 3080.730 ;
        RECT 1994.200 3080.410 1994.460 3080.730 ;
        RECT 1994.260 3020.970 1994.400 3080.410 ;
        RECT 1994.260 3020.830 1999.460 3020.970 ;
        RECT 1999.320 3009.410 1999.460 3020.830 ;
        RECT 2000.770 3009.410 2001.050 3010.000 ;
        RECT 1999.320 3009.270 2001.050 3009.410 ;
        RECT 2000.770 3006.000 2001.050 3009.270 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT -4.800 3411.070 3.370 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 3.070 3409.330 3.370 3411.070 ;
        RECT 2563.390 3409.330 2563.770 3409.340 ;
        RECT 3.070 3409.030 2563.770 3409.330 ;
        RECT 2563.390 3409.020 2563.770 3409.030 ;
        RECT 2506.000 576.680 2510.000 577.280 ;
        RECT 2509.150 574.410 2509.450 576.680 ;
        RECT 2509.150 574.110 2510.370 574.410 ;
        RECT 2510.070 573.050 2510.370 574.110 ;
        RECT 2563.390 573.050 2563.770 573.060 ;
        RECT 2510.070 572.750 2563.770 573.050 ;
        RECT 2563.390 572.740 2563.770 572.750 ;
      LAYER via3 ;
        RECT 2563.420 3409.020 2563.740 3409.340 ;
        RECT 2563.420 572.740 2563.740 573.060 ;
      LAYER met4 ;
        RECT 2563.415 3409.015 2563.745 3409.345 ;
        RECT 2563.430 573.065 2563.730 3409.015 ;
        RECT 2563.415 572.735 2563.745 573.065 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 279.290 3119.060 279.610 3119.120 ;
        RECT 17.090 3118.920 279.610 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 279.290 3118.860 279.610 3118.920 ;
        RECT 279.290 1317.740 279.610 1317.800 ;
        RECT 393.370 1317.740 393.690 1317.800 ;
        RECT 279.290 1317.600 393.690 1317.740 ;
        RECT 279.290 1317.540 279.610 1317.600 ;
        RECT 393.370 1317.540 393.690 1317.600 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 279.320 3118.860 279.580 3119.120 ;
        RECT 279.320 1317.540 279.580 1317.800 ;
        RECT 393.400 1317.540 393.660 1317.800 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 279.320 3118.830 279.580 3119.150 ;
        RECT 279.380 1317.830 279.520 3118.830 ;
        RECT 279.320 1317.510 279.580 1317.830 ;
        RECT 393.400 1317.510 393.660 1317.830 ;
        RECT 393.460 1317.005 393.600 1317.510 ;
        RECT 393.390 1316.635 393.670 1317.005 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
        RECT 393.390 1316.680 393.670 1316.960 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
        RECT 393.365 1316.970 393.695 1316.985 ;
        RECT 410.000 1316.970 414.000 1317.120 ;
        RECT 393.365 1316.670 414.000 1316.970 ;
        RECT 393.365 1316.655 393.695 1316.670 ;
        RECT 410.000 1316.520 414.000 1316.670 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 127.490 2836.180 127.810 2836.240 ;
        RECT 17.090 2836.040 127.810 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 127.490 2835.980 127.810 2836.040 ;
        RECT 127.490 489.840 127.810 489.900 ;
        RECT 647.290 489.840 647.610 489.900 ;
        RECT 127.490 489.700 647.610 489.840 ;
        RECT 127.490 489.640 127.810 489.700 ;
        RECT 647.290 489.640 647.610 489.700 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 127.520 2835.980 127.780 2836.240 ;
        RECT 127.520 489.640 127.780 489.900 ;
        RECT 647.320 489.640 647.580 489.900 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 127.520 2835.950 127.780 2836.270 ;
        RECT 127.580 489.930 127.720 2835.950 ;
        RECT 647.450 510.340 647.730 514.000 ;
        RECT 647.380 510.000 647.730 510.340 ;
        RECT 647.380 489.930 647.520 510.000 ;
        RECT 127.520 489.610 127.780 489.930 ;
        RECT 647.320 489.610 647.580 489.930 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 2546.500 16.030 2546.560 ;
        RECT 45.610 2546.500 45.930 2546.560 ;
        RECT 15.710 2546.360 45.930 2546.500 ;
        RECT 15.710 2546.300 16.030 2546.360 ;
        RECT 45.610 2546.300 45.930 2546.360 ;
        RECT 45.610 1614.560 45.930 1614.620 ;
        RECT 393.370 1614.560 393.690 1614.620 ;
        RECT 45.610 1614.420 393.690 1614.560 ;
        RECT 45.610 1614.360 45.930 1614.420 ;
        RECT 393.370 1614.360 393.690 1614.420 ;
      LAYER via ;
        RECT 15.740 2546.300 16.000 2546.560 ;
        RECT 45.640 2546.300 45.900 2546.560 ;
        RECT 45.640 1614.360 45.900 1614.620 ;
        RECT 393.400 1614.360 393.660 1614.620 ;
      LAYER met2 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
        RECT 15.800 2546.590 15.940 2549.475 ;
        RECT 15.740 2546.270 16.000 2546.590 ;
        RECT 45.640 2546.270 45.900 2546.590 ;
        RECT 45.700 1614.650 45.840 2546.270 ;
        RECT 45.640 1614.330 45.900 1614.650 ;
        RECT 393.400 1614.330 393.660 1614.650 ;
        RECT 393.460 1609.405 393.600 1614.330 ;
        RECT 393.390 1609.035 393.670 1609.405 ;
      LAYER via2 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
        RECT 393.390 1609.080 393.670 1609.360 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
        RECT 393.365 1609.370 393.695 1609.385 ;
        RECT 410.000 1609.370 414.000 1609.520 ;
        RECT 393.365 1609.070 414.000 1609.370 ;
        RECT 393.365 1609.055 393.695 1609.070 ;
        RECT 410.000 1608.920 414.000 1609.070 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2506.000 2457.560 2510.000 2458.160 ;
        RECT 2507.310 2455.300 2507.610 2457.560 ;
        RECT 2507.270 2454.980 2507.650 2455.300 ;
        RECT 168.630 2436.250 169.010 2436.260 ;
        RECT 233.950 2436.250 234.330 2436.260 ;
        RECT 168.630 2435.950 234.330 2436.250 ;
        RECT 168.630 2435.940 169.010 2435.950 ;
        RECT 233.950 2435.940 234.330 2435.950 ;
        RECT 89.510 2429.450 89.890 2429.460 ;
        RECT 137.350 2429.450 137.730 2429.460 ;
        RECT 89.510 2429.150 137.730 2429.450 ;
        RECT 89.510 2429.140 89.890 2429.150 ;
        RECT 137.350 2429.140 137.730 2429.150 ;
        RECT 50.870 2262.850 51.250 2262.860 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 3.070 2262.550 51.250 2262.850 ;
        RECT 3.070 2262.170 3.370 2262.550 ;
        RECT 50.870 2262.540 51.250 2262.550 ;
        RECT -4.800 2261.870 3.370 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
      LAYER via3 ;
        RECT 2507.300 2454.980 2507.620 2455.300 ;
        RECT 168.660 2435.940 168.980 2436.260 ;
        RECT 233.980 2435.940 234.300 2436.260 ;
        RECT 89.540 2429.140 89.860 2429.460 ;
        RECT 137.380 2429.140 137.700 2429.460 ;
        RECT 50.900 2262.540 51.220 2262.860 ;
      LAYER met4 ;
        RECT 2507.295 2454.975 2507.625 2455.305 ;
        RECT 2507.310 2436.690 2507.610 2454.975 ;
        RECT 136.950 2435.510 138.130 2436.690 ;
        RECT 168.230 2435.510 169.410 2436.690 ;
        RECT 233.975 2435.935 234.305 2436.265 ;
        RECT 50.470 2428.710 51.650 2429.890 ;
        RECT 89.110 2428.710 90.290 2429.890 ;
        RECT 137.390 2429.465 137.690 2435.510 ;
        RECT 137.375 2429.135 137.705 2429.465 ;
        RECT 50.910 2262.865 51.210 2428.710 ;
        RECT 233.990 2423.090 234.290 2435.935 ;
        RECT 2506.870 2435.510 2508.050 2436.690 ;
        RECT 233.550 2421.910 234.730 2423.090 ;
        RECT 50.895 2262.535 51.225 2262.865 ;
      LAYER met5 ;
        RECT 136.740 2435.300 169.620 2436.900 ;
        RECT 2447.780 2435.300 2477.900 2436.900 ;
        RECT 288.540 2431.900 302.100 2433.500 ;
        RECT 288.540 2430.100 290.140 2431.900 ;
        RECT 50.260 2428.500 90.500 2430.100 ;
        RECT 264.620 2428.500 290.140 2430.100 ;
        RECT 300.500 2430.100 302.100 2431.900 ;
        RECT 304.180 2431.900 314.980 2433.500 ;
        RECT 304.180 2430.100 305.780 2431.900 ;
        RECT 300.500 2428.500 305.780 2430.100 ;
        RECT 313.380 2430.100 314.980 2431.900 ;
        RECT 476.220 2431.900 491.620 2433.500 ;
        RECT 313.380 2428.500 424.460 2430.100 ;
        RECT 264.620 2423.300 266.220 2428.500 ;
        RECT 233.340 2421.700 266.220 2423.300 ;
        RECT 422.860 2423.300 424.460 2428.500 ;
        RECT 476.220 2423.300 477.820 2431.900 ;
        RECT 422.860 2421.700 477.820 2423.300 ;
        RECT 490.020 2423.300 491.620 2431.900 ;
        RECT 2447.780 2423.300 2449.380 2435.300 ;
        RECT 2476.300 2433.500 2477.900 2435.300 ;
        RECT 2497.460 2435.300 2508.260 2436.900 ;
        RECT 2497.460 2433.500 2499.060 2435.300 ;
        RECT 2476.300 2431.900 2499.060 2433.500 ;
        RECT 490.020 2421.700 524.740 2423.300 ;
        RECT 523.140 2419.900 524.740 2421.700 ;
        RECT 2441.340 2421.700 2449.380 2423.300 ;
        RECT 2441.340 2419.900 2442.940 2421.700 ;
        RECT 523.140 2418.300 542.220 2419.900 ;
        RECT 540.620 2413.100 542.220 2418.300 ;
        RECT 545.220 2418.300 573.500 2419.900 ;
        RECT 545.220 2413.100 546.820 2418.300 ;
        RECT 540.620 2411.500 546.820 2413.100 ;
        RECT 571.900 2413.100 573.500 2418.300 ;
        RECT 575.580 2418.300 638.820 2419.900 ;
        RECT 575.580 2413.100 577.180 2418.300 ;
        RECT 571.900 2411.500 577.180 2413.100 ;
        RECT 637.220 2413.100 638.820 2418.300 ;
        RECT 641.820 2418.300 670.100 2419.900 ;
        RECT 641.820 2413.100 643.420 2418.300 ;
        RECT 637.220 2411.500 643.420 2413.100 ;
        RECT 668.500 2413.100 670.100 2418.300 ;
        RECT 672.180 2418.300 735.420 2419.900 ;
        RECT 672.180 2413.100 673.780 2418.300 ;
        RECT 668.500 2411.500 673.780 2413.100 ;
        RECT 733.820 2413.100 735.420 2418.300 ;
        RECT 738.420 2418.300 766.700 2419.900 ;
        RECT 738.420 2413.100 740.020 2418.300 ;
        RECT 733.820 2411.500 740.020 2413.100 ;
        RECT 765.100 2413.100 766.700 2418.300 ;
        RECT 768.780 2418.300 832.020 2419.900 ;
        RECT 768.780 2413.100 770.380 2418.300 ;
        RECT 765.100 2411.500 770.380 2413.100 ;
        RECT 830.420 2413.100 832.020 2418.300 ;
        RECT 835.020 2418.300 863.300 2419.900 ;
        RECT 835.020 2413.100 836.620 2418.300 ;
        RECT 830.420 2411.500 836.620 2413.100 ;
        RECT 861.700 2413.100 863.300 2418.300 ;
        RECT 865.380 2418.300 928.620 2419.900 ;
        RECT 865.380 2413.100 866.980 2418.300 ;
        RECT 861.700 2411.500 866.980 2413.100 ;
        RECT 927.020 2413.100 928.620 2418.300 ;
        RECT 931.620 2418.300 959.900 2419.900 ;
        RECT 931.620 2413.100 933.220 2418.300 ;
        RECT 927.020 2411.500 933.220 2413.100 ;
        RECT 958.300 2413.100 959.900 2418.300 ;
        RECT 961.980 2418.300 1025.220 2419.900 ;
        RECT 961.980 2413.100 963.580 2418.300 ;
        RECT 958.300 2411.500 963.580 2413.100 ;
        RECT 1023.620 2413.100 1025.220 2418.300 ;
        RECT 1028.220 2418.300 1056.500 2419.900 ;
        RECT 1028.220 2413.100 1029.820 2418.300 ;
        RECT 1023.620 2411.500 1029.820 2413.100 ;
        RECT 1054.900 2413.100 1056.500 2418.300 ;
        RECT 1058.580 2418.300 1121.820 2419.900 ;
        RECT 1058.580 2413.100 1060.180 2418.300 ;
        RECT 1054.900 2411.500 1060.180 2413.100 ;
        RECT 1120.220 2413.100 1121.820 2418.300 ;
        RECT 1124.820 2418.300 1153.100 2419.900 ;
        RECT 1124.820 2413.100 1126.420 2418.300 ;
        RECT 1120.220 2411.500 1126.420 2413.100 ;
        RECT 1151.500 2413.100 1153.100 2418.300 ;
        RECT 1155.180 2418.300 1218.420 2419.900 ;
        RECT 1155.180 2413.100 1156.780 2418.300 ;
        RECT 1151.500 2411.500 1156.780 2413.100 ;
        RECT 1216.820 2413.100 1218.420 2418.300 ;
        RECT 1221.420 2418.300 1249.700 2419.900 ;
        RECT 1221.420 2413.100 1223.020 2418.300 ;
        RECT 1216.820 2411.500 1223.020 2413.100 ;
        RECT 1248.100 2413.100 1249.700 2418.300 ;
        RECT 1251.780 2418.300 1315.020 2419.900 ;
        RECT 1251.780 2413.100 1253.380 2418.300 ;
        RECT 1248.100 2411.500 1253.380 2413.100 ;
        RECT 1313.420 2413.100 1315.020 2418.300 ;
        RECT 1318.020 2418.300 1346.300 2419.900 ;
        RECT 1318.020 2413.100 1319.620 2418.300 ;
        RECT 1313.420 2411.500 1319.620 2413.100 ;
        RECT 1344.700 2413.100 1346.300 2418.300 ;
        RECT 1348.380 2418.300 1411.620 2419.900 ;
        RECT 1348.380 2413.100 1349.980 2418.300 ;
        RECT 1344.700 2411.500 1349.980 2413.100 ;
        RECT 1410.020 2413.100 1411.620 2418.300 ;
        RECT 1414.620 2418.300 1442.900 2419.900 ;
        RECT 1414.620 2413.100 1416.220 2418.300 ;
        RECT 1410.020 2411.500 1416.220 2413.100 ;
        RECT 1441.300 2413.100 1442.900 2418.300 ;
        RECT 1444.980 2418.300 1508.220 2419.900 ;
        RECT 1444.980 2413.100 1446.580 2418.300 ;
        RECT 1441.300 2411.500 1446.580 2413.100 ;
        RECT 1506.620 2413.100 1508.220 2418.300 ;
        RECT 1511.220 2418.300 1539.500 2419.900 ;
        RECT 1511.220 2413.100 1512.820 2418.300 ;
        RECT 1506.620 2411.500 1512.820 2413.100 ;
        RECT 1537.900 2413.100 1539.500 2418.300 ;
        RECT 1541.580 2418.300 1604.820 2419.900 ;
        RECT 1541.580 2413.100 1543.180 2418.300 ;
        RECT 1537.900 2411.500 1543.180 2413.100 ;
        RECT 1603.220 2413.100 1604.820 2418.300 ;
        RECT 1607.820 2418.300 1636.100 2419.900 ;
        RECT 1607.820 2413.100 1609.420 2418.300 ;
        RECT 1603.220 2411.500 1609.420 2413.100 ;
        RECT 1634.500 2413.100 1636.100 2418.300 ;
        RECT 1638.180 2418.300 1701.420 2419.900 ;
        RECT 1638.180 2413.100 1639.780 2418.300 ;
        RECT 1634.500 2411.500 1639.780 2413.100 ;
        RECT 1699.820 2413.100 1701.420 2418.300 ;
        RECT 1704.420 2418.300 1732.700 2419.900 ;
        RECT 1704.420 2413.100 1706.020 2418.300 ;
        RECT 1699.820 2411.500 1706.020 2413.100 ;
        RECT 1731.100 2413.100 1732.700 2418.300 ;
        RECT 1734.780 2418.300 1798.020 2419.900 ;
        RECT 1734.780 2413.100 1736.380 2418.300 ;
        RECT 1731.100 2411.500 1736.380 2413.100 ;
        RECT 1796.420 2413.100 1798.020 2418.300 ;
        RECT 1801.020 2418.300 1829.300 2419.900 ;
        RECT 1801.020 2413.100 1802.620 2418.300 ;
        RECT 1796.420 2411.500 1802.620 2413.100 ;
        RECT 1827.700 2413.100 1829.300 2418.300 ;
        RECT 1831.380 2418.300 1894.620 2419.900 ;
        RECT 1831.380 2413.100 1832.980 2418.300 ;
        RECT 1827.700 2411.500 1832.980 2413.100 ;
        RECT 1893.020 2413.100 1894.620 2418.300 ;
        RECT 1897.620 2418.300 1925.900 2419.900 ;
        RECT 1897.620 2413.100 1899.220 2418.300 ;
        RECT 1893.020 2411.500 1899.220 2413.100 ;
        RECT 1924.300 2413.100 1925.900 2418.300 ;
        RECT 1927.980 2418.300 1991.220 2419.900 ;
        RECT 1927.980 2413.100 1929.580 2418.300 ;
        RECT 1924.300 2411.500 1929.580 2413.100 ;
        RECT 1989.620 2413.100 1991.220 2418.300 ;
        RECT 1994.220 2418.300 2022.500 2419.900 ;
        RECT 1994.220 2413.100 1995.820 2418.300 ;
        RECT 1989.620 2411.500 1995.820 2413.100 ;
        RECT 2020.900 2413.100 2022.500 2418.300 ;
        RECT 2024.580 2418.300 2087.820 2419.900 ;
        RECT 2024.580 2413.100 2026.180 2418.300 ;
        RECT 2020.900 2411.500 2026.180 2413.100 ;
        RECT 2086.220 2413.100 2087.820 2418.300 ;
        RECT 2090.820 2418.300 2119.100 2419.900 ;
        RECT 2090.820 2413.100 2092.420 2418.300 ;
        RECT 2086.220 2411.500 2092.420 2413.100 ;
        RECT 2117.500 2413.100 2119.100 2418.300 ;
        RECT 2121.180 2418.300 2184.420 2419.900 ;
        RECT 2121.180 2413.100 2122.780 2418.300 ;
        RECT 2117.500 2411.500 2122.780 2413.100 ;
        RECT 2182.820 2413.100 2184.420 2418.300 ;
        RECT 2187.420 2418.300 2215.700 2419.900 ;
        RECT 2187.420 2413.100 2189.020 2418.300 ;
        RECT 2182.820 2411.500 2189.020 2413.100 ;
        RECT 2214.100 2413.100 2215.700 2418.300 ;
        RECT 2217.780 2418.300 2281.020 2419.900 ;
        RECT 2217.780 2413.100 2219.380 2418.300 ;
        RECT 2214.100 2411.500 2219.380 2413.100 ;
        RECT 2279.420 2413.100 2281.020 2418.300 ;
        RECT 2284.020 2418.300 2312.300 2419.900 ;
        RECT 2284.020 2413.100 2285.620 2418.300 ;
        RECT 2279.420 2411.500 2285.620 2413.100 ;
        RECT 2310.700 2413.100 2312.300 2418.300 ;
        RECT 2314.380 2418.300 2377.620 2419.900 ;
        RECT 2314.380 2413.100 2315.980 2418.300 ;
        RECT 2376.020 2416.500 2377.620 2418.300 ;
        RECT 2393.500 2418.300 2442.940 2419.900 ;
        RECT 2393.500 2416.500 2395.100 2418.300 ;
        RECT 2376.020 2414.900 2395.100 2416.500 ;
        RECT 2310.700 2411.500 2315.980 2413.100 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 1973.600 16.950 1973.660 ;
        RECT 349.210 1973.600 349.530 1973.660 ;
        RECT 16.630 1973.460 349.530 1973.600 ;
        RECT 16.630 1973.400 16.950 1973.460 ;
        RECT 349.210 1973.400 349.530 1973.460 ;
        RECT 349.210 489.160 349.530 489.220 ;
        RECT 893.850 489.160 894.170 489.220 ;
        RECT 349.210 489.020 894.170 489.160 ;
        RECT 349.210 488.960 349.530 489.020 ;
        RECT 893.850 488.960 894.170 489.020 ;
      LAYER via ;
        RECT 16.660 1973.400 16.920 1973.660 ;
        RECT 349.240 1973.400 349.500 1973.660 ;
        RECT 349.240 488.960 349.500 489.220 ;
        RECT 893.880 488.960 894.140 489.220 ;
      LAYER met2 ;
        RECT 16.650 1974.875 16.930 1975.245 ;
        RECT 16.720 1973.690 16.860 1974.875 ;
        RECT 16.660 1973.370 16.920 1973.690 ;
        RECT 349.240 1973.370 349.500 1973.690 ;
        RECT 349.300 489.250 349.440 1973.370 ;
        RECT 894.010 510.340 894.290 514.000 ;
        RECT 893.940 510.000 894.290 510.340 ;
        RECT 893.940 489.250 894.080 510.000 ;
        RECT 349.240 488.930 349.500 489.250 ;
        RECT 893.880 488.930 894.140 489.250 ;
      LAYER via2 ;
        RECT 16.650 1974.920 16.930 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.625 1975.210 16.955 1975.225 ;
        RECT -4.800 1974.910 16.955 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.625 1974.895 16.955 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 384.630 2863.720 384.950 2863.780 ;
        RECT 393.830 2863.720 394.150 2863.780 ;
        RECT 384.630 2863.580 394.150 2863.720 ;
        RECT 384.630 2863.520 384.950 2863.580 ;
        RECT 393.830 2863.520 394.150 2863.580 ;
        RECT 427.870 507.180 428.190 507.240 ;
        RECT 2476.250 507.180 2476.570 507.240 ;
        RECT 427.870 507.040 2476.570 507.180 ;
        RECT 427.870 506.980 428.190 507.040 ;
        RECT 2476.250 506.980 2476.570 507.040 ;
      LAYER via ;
        RECT 384.660 2863.520 384.920 2863.780 ;
        RECT 393.860 2863.520 394.120 2863.780 ;
        RECT 427.900 506.980 428.160 507.240 ;
        RECT 2476.280 506.980 2476.540 507.240 ;
      LAYER met2 ;
        RECT 393.850 2869.755 394.130 2870.125 ;
        RECT 393.920 2863.810 394.060 2869.755 ;
        RECT 384.660 2863.490 384.920 2863.810 ;
        RECT 393.860 2863.490 394.120 2863.810 ;
        RECT 384.720 509.845 384.860 2863.490 ;
        RECT 2901.310 557.075 2901.590 557.445 ;
        RECT 2901.380 510.525 2901.520 557.075 ;
        RECT 2476.270 510.155 2476.550 510.525 ;
        RECT 2901.310 510.155 2901.590 510.525 ;
        RECT 384.650 509.475 384.930 509.845 ;
        RECT 427.890 509.475 428.170 509.845 ;
        RECT 427.960 507.270 428.100 509.475 ;
        RECT 2476.340 507.270 2476.480 510.155 ;
        RECT 427.900 506.950 428.160 507.270 ;
        RECT 2476.280 506.950 2476.540 507.270 ;
      LAYER via2 ;
        RECT 393.850 2869.800 394.130 2870.080 ;
        RECT 2901.310 557.120 2901.590 557.400 ;
        RECT 2476.270 510.200 2476.550 510.480 ;
        RECT 2901.310 510.200 2901.590 510.480 ;
        RECT 384.650 509.520 384.930 509.800 ;
        RECT 427.890 509.520 428.170 509.800 ;
      LAYER met3 ;
        RECT 393.825 2870.090 394.155 2870.105 ;
        RECT 410.000 2870.090 414.000 2870.240 ;
        RECT 393.825 2869.790 414.000 2870.090 ;
        RECT 393.825 2869.775 394.155 2869.790 ;
        RECT 410.000 2869.640 414.000 2869.790 ;
        RECT 2901.285 557.410 2901.615 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2901.285 557.110 2924.800 557.410 ;
        RECT 2901.285 557.095 2901.615 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2476.245 510.490 2476.575 510.505 ;
        RECT 2901.285 510.490 2901.615 510.505 ;
        RECT 2476.245 510.190 2901.615 510.490 ;
        RECT 2476.245 510.175 2476.575 510.190 ;
        RECT 2901.285 510.175 2901.615 510.190 ;
        RECT 384.625 509.810 384.955 509.825 ;
        RECT 427.865 509.810 428.195 509.825 ;
        RECT 384.625 509.510 428.195 509.810 ;
        RECT 384.625 509.495 384.955 509.510 ;
        RECT 427.865 509.495 428.195 509.510 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1683.920 17.410 1683.980 ;
        RECT 363.010 1683.920 363.330 1683.980 ;
        RECT 17.090 1683.780 363.330 1683.920 ;
        RECT 17.090 1683.720 17.410 1683.780 ;
        RECT 363.010 1683.720 363.330 1683.780 ;
        RECT 363.010 503.780 363.330 503.840 ;
        RECT 2339.170 503.780 2339.490 503.840 ;
        RECT 363.010 503.640 2339.490 503.780 ;
        RECT 363.010 503.580 363.330 503.640 ;
        RECT 2339.170 503.580 2339.490 503.640 ;
      LAYER via ;
        RECT 17.120 1683.720 17.380 1683.980 ;
        RECT 363.040 1683.720 363.300 1683.980 ;
        RECT 363.040 503.580 363.300 503.840 ;
        RECT 2339.200 503.580 2339.460 503.840 ;
      LAYER met2 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
        RECT 17.180 1684.010 17.320 1687.235 ;
        RECT 17.120 1683.690 17.380 1684.010 ;
        RECT 363.040 1683.690 363.300 1684.010 ;
        RECT 363.100 503.870 363.240 1683.690 ;
        RECT 2339.330 510.340 2339.610 514.000 ;
        RECT 2339.260 510.000 2339.610 510.340 ;
        RECT 2339.260 503.870 2339.400 510.000 ;
        RECT 363.040 503.550 363.300 503.870 ;
        RECT 2339.200 503.550 2339.460 503.870 ;
      LAYER via2 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 106.790 3024.200 107.110 3024.260 ;
        RECT 1283.930 3024.200 1284.250 3024.260 ;
        RECT 106.790 3024.060 1284.250 3024.200 ;
        RECT 106.790 3024.000 107.110 3024.060 ;
        RECT 1283.930 3024.000 1284.250 3024.060 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 106.790 1476.520 107.110 1476.580 ;
        RECT 17.090 1476.380 107.110 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 106.790 1476.320 107.110 1476.380 ;
      LAYER via ;
        RECT 106.820 3024.000 107.080 3024.260 ;
        RECT 1283.960 3024.000 1284.220 3024.260 ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 106.820 1476.320 107.080 1476.580 ;
      LAYER met2 ;
        RECT 106.820 3023.970 107.080 3024.290 ;
        RECT 1283.960 3023.970 1284.220 3024.290 ;
        RECT 106.880 1476.610 107.020 3023.970 ;
        RECT 1284.020 3010.000 1284.160 3023.970 ;
        RECT 1284.020 3009.340 1284.370 3010.000 ;
        RECT 1284.090 3006.000 1284.370 3009.340 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 106.820 1476.290 107.080 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1256.200 17.410 1256.260 ;
        RECT 342.310 1256.200 342.630 1256.260 ;
        RECT 17.090 1256.060 342.630 1256.200 ;
        RECT 17.090 1256.000 17.410 1256.060 ;
        RECT 342.310 1256.000 342.630 1256.060 ;
        RECT 342.310 827.460 342.630 827.520 ;
        RECT 393.370 827.460 393.690 827.520 ;
        RECT 342.310 827.320 393.690 827.460 ;
        RECT 342.310 827.260 342.630 827.320 ;
        RECT 393.370 827.260 393.690 827.320 ;
      LAYER via ;
        RECT 17.120 1256.000 17.380 1256.260 ;
        RECT 342.340 1256.000 342.600 1256.260 ;
        RECT 342.340 827.260 342.600 827.520 ;
        RECT 393.400 827.260 393.660 827.520 ;
      LAYER met2 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
        RECT 17.120 1255.970 17.380 1256.115 ;
        RECT 342.340 1255.970 342.600 1256.290 ;
        RECT 342.400 827.550 342.540 1255.970 ;
        RECT 342.340 827.230 342.600 827.550 ;
        RECT 393.400 827.230 393.660 827.550 ;
        RECT 393.460 824.685 393.600 827.230 ;
        RECT 393.390 824.315 393.670 824.685 ;
      LAYER via2 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
        RECT 393.390 824.360 393.670 824.640 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
        RECT 393.365 824.650 393.695 824.665 ;
        RECT 410.000 824.650 414.000 824.800 ;
        RECT 393.365 824.350 414.000 824.650 ;
        RECT 393.365 824.335 393.695 824.350 ;
        RECT 410.000 824.200 414.000 824.350 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 3024.540 286.510 3024.600 ;
        RECT 1383.290 3024.540 1383.610 3024.600 ;
        RECT 286.190 3024.400 1383.610 3024.540 ;
        RECT 286.190 3024.340 286.510 3024.400 ;
        RECT 1383.290 3024.340 1383.610 3024.400 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 286.190 1041.660 286.510 1041.720 ;
        RECT 17.090 1041.520 286.510 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 286.190 1041.460 286.510 1041.520 ;
      LAYER via ;
        RECT 286.220 3024.340 286.480 3024.600 ;
        RECT 1383.320 3024.340 1383.580 3024.600 ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 286.220 1041.460 286.480 1041.720 ;
      LAYER met2 ;
        RECT 286.220 3024.310 286.480 3024.630 ;
        RECT 1383.320 3024.310 1383.580 3024.630 ;
        RECT 286.280 1041.750 286.420 3024.310 ;
        RECT 1383.380 3010.000 1383.520 3024.310 ;
        RECT 1383.380 3009.340 1383.730 3010.000 ;
        RECT 1383.450 3006.000 1383.730 3009.340 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 286.220 1041.430 286.480 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 362.090 3026.580 362.410 3026.640 ;
        RECT 1234.250 3026.580 1234.570 3026.640 ;
        RECT 362.090 3026.440 1234.570 3026.580 ;
        RECT 362.090 3026.380 362.410 3026.440 ;
        RECT 1234.250 3026.380 1234.570 3026.440 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 362.090 827.800 362.410 827.860 ;
        RECT 17.550 827.660 362.410 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 362.090 827.600 362.410 827.660 ;
      LAYER via ;
        RECT 362.120 3026.380 362.380 3026.640 ;
        RECT 1234.280 3026.380 1234.540 3026.640 ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 362.120 827.600 362.380 827.860 ;
      LAYER met2 ;
        RECT 362.120 3026.350 362.380 3026.670 ;
        RECT 1234.280 3026.350 1234.540 3026.670 ;
        RECT 362.180 827.890 362.320 3026.350 ;
        RECT 1234.340 3010.000 1234.480 3026.350 ;
        RECT 1234.340 3009.340 1234.690 3010.000 ;
        RECT 1234.410 3006.000 1234.690 3009.340 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 362.120 827.570 362.380 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 607.480 17.410 607.540 ;
        RECT 58.490 607.480 58.810 607.540 ;
        RECT 17.090 607.340 58.810 607.480 ;
        RECT 17.090 607.280 17.410 607.340 ;
        RECT 58.490 607.280 58.810 607.340 ;
        RECT 58.490 503.440 58.810 503.500 ;
        RECT 1425.610 503.440 1425.930 503.500 ;
        RECT 58.490 503.300 1425.930 503.440 ;
        RECT 58.490 503.240 58.810 503.300 ;
        RECT 1425.610 503.240 1425.930 503.300 ;
      LAYER via ;
        RECT 17.120 607.280 17.380 607.540 ;
        RECT 58.520 607.280 58.780 607.540 ;
        RECT 58.520 503.240 58.780 503.500 ;
        RECT 1425.640 503.240 1425.900 503.500 ;
      LAYER met2 ;
        RECT 17.110 610.115 17.390 610.485 ;
        RECT 17.180 607.570 17.320 610.115 ;
        RECT 17.120 607.250 17.380 607.570 ;
        RECT 58.520 607.250 58.780 607.570 ;
        RECT 58.580 503.530 58.720 607.250 ;
        RECT 1425.770 510.340 1426.050 514.000 ;
        RECT 1425.700 510.000 1426.050 510.340 ;
        RECT 1425.700 503.530 1425.840 510.000 ;
        RECT 58.520 503.210 58.780 503.530 ;
        RECT 1425.640 503.210 1425.900 503.530 ;
      LAYER via2 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 399.995 17.390 400.365 ;
        RECT 17.180 394.925 17.320 399.995 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 17.110 400.040 17.390 400.320 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 2506.000 2512.410 2510.000 2512.560 ;
        RECT 2553.270 2512.410 2553.650 2512.420 ;
        RECT 2506.000 2512.110 2553.650 2512.410 ;
        RECT 2506.000 2511.960 2510.000 2512.110 ;
        RECT 2553.270 2512.100 2553.650 2512.110 ;
        RECT 17.085 400.330 17.415 400.345 ;
        RECT 2553.270 400.330 2553.650 400.340 ;
        RECT 17.085 400.030 2553.650 400.330 ;
        RECT 17.085 400.015 17.415 400.030 ;
        RECT 2553.270 400.020 2553.650 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
      LAYER via3 ;
        RECT 2553.300 2512.100 2553.620 2512.420 ;
        RECT 2553.300 400.020 2553.620 400.340 ;
      LAYER met4 ;
        RECT 2553.295 2512.095 2553.625 2512.425 ;
        RECT 2553.310 400.345 2553.610 2512.095 ;
        RECT 2553.295 400.015 2553.625 400.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2444.990 3020.035 2445.270 3020.405 ;
        RECT 2445.060 3010.000 2445.200 3020.035 ;
        RECT 2445.060 3009.340 2445.410 3010.000 ;
        RECT 2445.130 3006.000 2445.410 3009.340 ;
      LAYER via2 ;
        RECT 2444.990 3020.080 2445.270 3020.360 ;
      LAYER met3 ;
        RECT 2141.110 3033.290 2141.490 3033.300 ;
        RECT 1946.110 3032.990 2141.490 3033.290 ;
        RECT 1946.110 3032.610 1946.410 3032.990 ;
        RECT 2141.110 3032.980 2141.490 3032.990 ;
        RECT 2188.950 3033.290 2189.330 3033.300 ;
        RECT 2293.830 3033.290 2294.210 3033.300 ;
        RECT 2188.950 3032.990 2294.210 3033.290 ;
        RECT 2188.950 3032.980 2189.330 3032.990 ;
        RECT 2293.830 3032.980 2294.210 3032.990 ;
        RECT 1901.030 3032.310 1946.410 3032.610 ;
        RECT 1901.030 3031.930 1901.330 3032.310 ;
        RECT 1656.310 3031.630 1901.330 3031.930 ;
        RECT 1179.710 3031.250 1180.090 3031.260 ;
        RECT 1222.030 3031.250 1222.410 3031.260 ;
        RECT 1179.710 3030.950 1222.410 3031.250 ;
        RECT 1179.710 3030.940 1180.090 3030.950 ;
        RECT 1222.030 3030.940 1222.410 3030.950 ;
        RECT 1269.870 3031.250 1270.250 3031.260 ;
        RECT 1364.630 3031.250 1365.010 3031.260 ;
        RECT 1269.870 3030.950 1365.010 3031.250 ;
        RECT 1269.870 3030.940 1270.250 3030.950 ;
        RECT 1364.630 3030.940 1365.010 3030.950 ;
        RECT 1366.470 3031.250 1366.850 3031.260 ;
        RECT 1656.310 3031.250 1656.610 3031.630 ;
        RECT 1366.470 3030.950 1656.610 3031.250 ;
        RECT 1366.470 3030.940 1366.850 3030.950 ;
        RECT 594.590 3030.570 594.970 3030.580 ;
        RECT 643.350 3030.570 643.730 3030.580 ;
        RECT 594.590 3030.270 643.730 3030.570 ;
        RECT 594.590 3030.260 594.970 3030.270 ;
        RECT 643.350 3030.260 643.730 3030.270 ;
        RECT 692.110 3030.570 692.490 3030.580 ;
        RECT 785.950 3030.570 786.330 3030.580 ;
        RECT 692.110 3030.270 786.330 3030.570 ;
        RECT 692.110 3030.260 692.490 3030.270 ;
        RECT 785.950 3030.260 786.330 3030.270 ;
        RECT 884.390 3030.570 884.770 3030.580 ;
        RECT 979.150 3030.570 979.530 3030.580 ;
        RECT 884.390 3030.270 979.530 3030.570 ;
        RECT 884.390 3030.260 884.770 3030.270 ;
        RECT 979.150 3030.260 979.530 3030.270 ;
        RECT 982.830 3030.570 983.210 3030.580 ;
        RECT 1035.270 3030.570 1035.650 3030.580 ;
        RECT 982.830 3030.270 1035.650 3030.570 ;
        RECT 982.830 3030.260 983.210 3030.270 ;
        RECT 1035.270 3030.260 1035.650 3030.270 ;
        RECT 445.550 3027.850 445.930 3027.860 ;
        RECT 451.070 3027.850 451.450 3027.860 ;
        RECT 445.550 3027.550 451.450 3027.850 ;
        RECT 445.550 3027.540 445.930 3027.550 ;
        RECT 451.070 3027.540 451.450 3027.550 ;
        RECT 548.590 3027.850 548.970 3027.860 ;
        RECT 592.750 3027.850 593.130 3027.860 ;
        RECT 548.590 3027.550 593.130 3027.850 ;
        RECT 548.590 3027.540 548.970 3027.550 ;
        RECT 592.750 3027.540 593.130 3027.550 ;
        RECT 788.710 3027.850 789.090 3027.860 ;
        RECT 882.550 3027.850 882.930 3027.860 ;
        RECT 788.710 3027.550 882.930 3027.850 ;
        RECT 788.710 3027.540 789.090 3027.550 ;
        RECT 882.550 3027.540 882.930 3027.550 ;
        RECT 2442.870 3020.370 2443.250 3020.380 ;
        RECT 2444.965 3020.370 2445.295 3020.385 ;
        RECT 2442.870 3020.070 2445.295 3020.370 ;
        RECT 2442.870 3020.060 2443.250 3020.070 ;
        RECT 2444.965 3020.055 2445.295 3020.070 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 320.430 179.330 320.810 179.340 ;
        RECT -4.800 179.030 320.810 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 320.430 179.020 320.810 179.030 ;
      LAYER via3 ;
        RECT 2141.140 3032.980 2141.460 3033.300 ;
        RECT 2188.980 3032.980 2189.300 3033.300 ;
        RECT 2293.860 3032.980 2294.180 3033.300 ;
        RECT 1179.740 3030.940 1180.060 3031.260 ;
        RECT 1222.060 3030.940 1222.380 3031.260 ;
        RECT 1269.900 3030.940 1270.220 3031.260 ;
        RECT 1364.660 3030.940 1364.980 3031.260 ;
        RECT 1366.500 3030.940 1366.820 3031.260 ;
        RECT 594.620 3030.260 594.940 3030.580 ;
        RECT 643.380 3030.260 643.700 3030.580 ;
        RECT 692.140 3030.260 692.460 3030.580 ;
        RECT 785.980 3030.260 786.300 3030.580 ;
        RECT 884.420 3030.260 884.740 3030.580 ;
        RECT 979.180 3030.260 979.500 3030.580 ;
        RECT 982.860 3030.260 983.180 3030.580 ;
        RECT 1035.300 3030.260 1035.620 3030.580 ;
        RECT 445.580 3027.540 445.900 3027.860 ;
        RECT 451.100 3027.540 451.420 3027.860 ;
        RECT 548.620 3027.540 548.940 3027.860 ;
        RECT 592.780 3027.540 593.100 3027.860 ;
        RECT 788.740 3027.540 789.060 3027.860 ;
        RECT 882.580 3027.540 882.900 3027.860 ;
        RECT 2442.900 3020.060 2443.220 3020.380 ;
        RECT 320.460 179.020 320.780 179.340 ;
      LAYER met4 ;
        RECT 2141.135 3032.975 2141.465 3033.305 ;
        RECT 2188.975 3032.975 2189.305 3033.305 ;
        RECT 2293.855 3032.975 2294.185 3033.305 ;
        RECT 1179.735 3030.935 1180.065 3031.265 ;
        RECT 1222.055 3030.935 1222.385 3031.265 ;
        RECT 1269.895 3030.935 1270.225 3031.265 ;
        RECT 1364.655 3030.935 1364.985 3031.265 ;
        RECT 1366.495 3030.935 1366.825 3031.265 ;
        RECT 594.615 3030.255 594.945 3030.585 ;
        RECT 643.375 3030.255 643.705 3030.585 ;
        RECT 692.135 3030.255 692.465 3030.585 ;
        RECT 785.975 3030.255 786.305 3030.585 ;
        RECT 884.415 3030.255 884.745 3030.585 ;
        RECT 979.175 3030.255 979.505 3030.585 ;
        RECT 982.855 3030.255 983.185 3030.585 ;
        RECT 1035.295 3030.255 1035.625 3030.585 ;
        RECT 594.630 3028.290 594.930 3030.255 ;
        RECT 643.390 3028.290 643.690 3030.255 ;
        RECT 692.150 3028.290 692.450 3030.255 ;
        RECT 785.990 3028.290 786.290 3030.255 ;
        RECT 884.430 3028.290 884.730 3030.255 ;
        RECT 979.190 3028.290 979.490 3030.255 ;
        RECT 982.870 3028.290 983.170 3030.255 ;
        RECT 320.030 3027.110 321.210 3028.290 ;
        RECT 445.150 3027.110 446.330 3028.290 ;
        RECT 450.670 3027.110 451.850 3028.290 ;
        RECT 548.615 3027.535 548.945 3027.865 ;
        RECT 320.470 179.345 320.770 3027.110 ;
        RECT 548.630 3024.890 548.930 3027.535 ;
        RECT 592.350 3027.110 593.530 3028.290 ;
        RECT 594.190 3027.110 595.370 3028.290 ;
        RECT 642.950 3027.110 644.130 3028.290 ;
        RECT 691.710 3027.110 692.890 3028.290 ;
        RECT 785.550 3027.110 786.730 3028.290 ;
        RECT 788.310 3027.110 789.490 3028.290 ;
        RECT 882.150 3027.110 883.330 3028.290 ;
        RECT 883.990 3027.110 885.170 3028.290 ;
        RECT 978.750 3027.110 979.930 3028.290 ;
        RECT 982.430 3027.110 983.610 3028.290 ;
        RECT 1035.310 3024.890 1035.610 3030.255 ;
        RECT 1179.750 3028.290 1180.050 3030.935 ;
        RECT 1222.070 3028.290 1222.370 3030.935 ;
        RECT 1269.910 3028.290 1270.210 3030.935 ;
        RECT 1364.670 3028.290 1364.970 3030.935 ;
        RECT 1366.510 3028.290 1366.810 3030.935 ;
        RECT 1179.310 3027.110 1180.490 3028.290 ;
        RECT 1221.630 3027.110 1222.810 3028.290 ;
        RECT 1269.470 3027.110 1270.650 3028.290 ;
        RECT 1364.230 3027.110 1365.410 3028.290 ;
        RECT 1366.070 3027.110 1367.250 3028.290 ;
        RECT 2141.150 3024.890 2141.450 3032.975 ;
        RECT 2188.990 3024.890 2189.290 3032.975 ;
        RECT 2293.870 3024.890 2294.170 3032.975 ;
        RECT 548.190 3023.710 549.370 3024.890 ;
        RECT 1034.870 3023.710 1036.050 3024.890 ;
        RECT 2140.710 3023.710 2141.890 3024.890 ;
        RECT 2188.550 3023.710 2189.730 3024.890 ;
        RECT 2293.430 3023.710 2294.610 3024.890 ;
        RECT 2442.470 3020.310 2443.650 3021.490 ;
        RECT 2442.895 3020.055 2443.225 3020.310 ;
        RECT 320.455 179.015 320.785 179.345 ;
      LAYER via4 ;
        RECT 2442.470 3020.310 2443.650 3021.490 ;
      LAYER met5 ;
        RECT 319.820 3026.900 446.540 3028.500 ;
        RECT 450.460 3026.900 498.060 3028.500 ;
        RECT 592.140 3026.900 595.580 3028.500 ;
        RECT 642.740 3026.900 693.100 3028.500 ;
        RECT 785.340 3026.900 789.700 3028.500 ;
        RECT 881.940 3026.900 885.380 3028.500 ;
        RECT 978.540 3026.900 983.820 3028.500 ;
        RECT 1124.820 3026.900 1180.700 3028.500 ;
        RECT 1221.420 3026.900 1270.860 3028.500 ;
        RECT 1364.020 3026.900 1367.460 3028.500 ;
        RECT 496.460 3025.100 498.060 3026.900 ;
        RECT 1124.820 3025.100 1126.420 3026.900 ;
        RECT 496.460 3023.500 549.580 3025.100 ;
        RECT 1034.660 3023.500 1126.420 3025.100 ;
        RECT 2140.500 3023.500 2189.940 3025.100 ;
        RECT 2293.220 3023.500 2382.220 3025.100 ;
        RECT 2380.620 3021.700 2382.220 3023.500 ;
        RECT 2380.620 3020.100 2443.860 3021.700 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1946.060 2519.810 1946.120 ;
        RECT 2867.250 1946.060 2867.570 1946.120 ;
        RECT 2519.490 1945.920 2867.570 1946.060 ;
        RECT 2519.490 1945.860 2519.810 1945.920 ;
        RECT 2867.250 1945.860 2867.570 1945.920 ;
        RECT 2867.250 793.460 2867.570 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2867.250 793.320 2899.310 793.460 ;
        RECT 2867.250 793.260 2867.570 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2519.520 1945.860 2519.780 1946.120 ;
        RECT 2867.280 1945.860 2867.540 1946.120 ;
        RECT 2867.280 793.260 2867.540 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2519.510 1946.315 2519.790 1946.685 ;
        RECT 2519.580 1946.150 2519.720 1946.315 ;
        RECT 2519.520 1945.830 2519.780 1946.150 ;
        RECT 2867.280 1945.830 2867.540 1946.150 ;
        RECT 2867.340 793.550 2867.480 1945.830 ;
        RECT 2867.280 793.230 2867.540 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2519.510 1946.360 2519.790 1946.640 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2506.000 1946.650 2510.000 1946.800 ;
        RECT 2519.485 1946.650 2519.815 1946.665 ;
        RECT 2506.000 1946.350 2519.815 1946.650 ;
        RECT 2506.000 1946.200 2510.000 1946.350 ;
        RECT 2519.485 1946.335 2519.815 1946.350 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2557.210 1021.600 2557.530 1021.660 ;
        RECT 2900.830 1021.600 2901.150 1021.660 ;
        RECT 2557.210 1021.460 2901.150 1021.600 ;
        RECT 2557.210 1021.400 2557.530 1021.460 ;
        RECT 2900.830 1021.400 2901.150 1021.460 ;
        RECT 1227.810 504.120 1228.130 504.180 ;
        RECT 2557.210 504.120 2557.530 504.180 ;
        RECT 1227.810 503.980 2557.530 504.120 ;
        RECT 1227.810 503.920 1228.130 503.980 ;
        RECT 2557.210 503.920 2557.530 503.980 ;
      LAYER via ;
        RECT 2557.240 1021.400 2557.500 1021.660 ;
        RECT 2900.860 1021.400 2901.120 1021.660 ;
        RECT 1227.840 503.920 1228.100 504.180 ;
        RECT 2557.240 503.920 2557.500 504.180 ;
      LAYER met2 ;
        RECT 2900.850 1026.275 2901.130 1026.645 ;
        RECT 2900.920 1021.690 2901.060 1026.275 ;
        RECT 2557.240 1021.370 2557.500 1021.690 ;
        RECT 2900.860 1021.370 2901.120 1021.690 ;
        RECT 1227.970 510.340 1228.250 514.000 ;
        RECT 1227.900 510.000 1228.250 510.340 ;
        RECT 1227.900 504.210 1228.040 510.000 ;
        RECT 2557.300 504.210 2557.440 1021.370 ;
        RECT 1227.840 503.890 1228.100 504.210 ;
        RECT 2557.240 503.890 2557.500 504.210 ;
      LAYER via2 ;
        RECT 2900.850 1026.320 2901.130 1026.600 ;
      LAYER met3 ;
        RECT 2900.825 1026.610 2901.155 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.825 1026.310 2924.800 1026.610 ;
        RECT 2900.825 1026.295 2901.155 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2839.190 1256.200 2839.510 1256.260 ;
        RECT 2900.830 1256.200 2901.150 1256.260 ;
        RECT 2839.190 1256.060 2901.150 1256.200 ;
        RECT 2839.190 1256.000 2839.510 1256.060 ;
        RECT 2900.830 1256.000 2901.150 1256.060 ;
        RECT 733.770 489.840 734.090 489.900 ;
        RECT 2839.190 489.840 2839.510 489.900 ;
        RECT 733.770 489.700 2839.510 489.840 ;
        RECT 733.770 489.640 734.090 489.700 ;
        RECT 2839.190 489.640 2839.510 489.700 ;
      LAYER via ;
        RECT 2839.220 1256.000 2839.480 1256.260 ;
        RECT 2900.860 1256.000 2901.120 1256.260 ;
        RECT 733.800 489.640 734.060 489.900 ;
        RECT 2839.220 489.640 2839.480 489.900 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 1256.290 2901.060 1260.875 ;
        RECT 2839.220 1255.970 2839.480 1256.290 ;
        RECT 2900.860 1255.970 2901.120 1256.290 ;
        RECT 733.930 510.340 734.210 514.000 ;
        RECT 733.860 510.000 734.210 510.340 ;
        RECT 733.860 489.930 734.000 510.000 ;
        RECT 2839.280 489.930 2839.420 1255.970 ;
        RECT 733.800 489.610 734.060 489.930 ;
        RECT 2839.220 489.610 2839.480 489.930 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2932.740 2519.810 2932.800 ;
        RECT 2701.190 2932.740 2701.510 2932.800 ;
        RECT 2519.490 2932.600 2701.510 2932.740 ;
        RECT 2519.490 2932.540 2519.810 2932.600 ;
        RECT 2701.190 2932.540 2701.510 2932.600 ;
        RECT 2701.190 1497.260 2701.510 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 2701.190 1497.120 2899.310 1497.260 ;
        RECT 2701.190 1497.060 2701.510 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 2519.520 2932.540 2519.780 2932.800 ;
        RECT 2701.220 2932.540 2701.480 2932.800 ;
        RECT 2701.220 1497.060 2701.480 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 2519.520 2932.685 2519.780 2932.830 ;
        RECT 2519.510 2932.315 2519.790 2932.685 ;
        RECT 2701.220 2932.510 2701.480 2932.830 ;
        RECT 2701.280 1497.350 2701.420 2932.510 ;
        RECT 2701.220 1497.030 2701.480 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2519.510 2932.360 2519.790 2932.640 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2506.000 2932.650 2510.000 2932.800 ;
        RECT 2519.485 2932.650 2519.815 2932.665 ;
        RECT 2506.000 2932.350 2519.815 2932.650 ;
        RECT 2506.000 2932.200 2510.000 2932.350 ;
        RECT 2519.485 2932.335 2519.815 2932.350 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1605.010 3017.740 1605.330 3017.800 ;
        RECT 1907.230 3017.740 1907.550 3017.800 ;
        RECT 1605.010 3017.600 1907.550 3017.740 ;
        RECT 1605.010 3017.540 1605.330 3017.600 ;
        RECT 1907.230 3017.540 1907.550 3017.600 ;
        RECT 1907.230 3011.960 1907.550 3012.020 ;
        RECT 2901.290 3011.960 2901.610 3012.020 ;
        RECT 1907.230 3011.820 2901.610 3011.960 ;
        RECT 1907.230 3011.760 1907.550 3011.820 ;
        RECT 2901.290 3011.760 2901.610 3011.820 ;
      LAYER via ;
        RECT 1605.040 3017.540 1605.300 3017.800 ;
        RECT 1907.260 3017.540 1907.520 3017.800 ;
        RECT 1907.260 3011.760 1907.520 3012.020 ;
        RECT 2901.320 3011.760 2901.580 3012.020 ;
      LAYER met2 ;
        RECT 1605.040 3017.510 1605.300 3017.830 ;
        RECT 1907.260 3017.510 1907.520 3017.830 ;
        RECT 1605.100 3010.000 1605.240 3017.510 ;
        RECT 1907.320 3012.050 1907.460 3017.510 ;
        RECT 1907.260 3011.730 1907.520 3012.050 ;
        RECT 2901.320 3011.730 2901.580 3012.050 ;
        RECT 1605.100 3009.340 1605.450 3010.000 ;
        RECT 1605.170 3006.000 1605.450 3009.340 ;
        RECT 2901.380 1730.445 2901.520 3011.730 ;
        RECT 2901.310 1730.075 2901.590 1730.445 ;
      LAYER via2 ;
        RECT 2901.310 1730.120 2901.590 1730.400 ;
      LAYER met3 ;
        RECT 2901.285 1730.410 2901.615 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2901.285 1730.110 2924.800 1730.410 ;
        RECT 2901.285 1730.095 2901.615 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 3008.560 593.330 3008.620 ;
        RECT 2535.590 3008.560 2535.910 3008.620 ;
        RECT 593.010 3008.420 2535.910 3008.560 ;
        RECT 593.010 3008.360 593.330 3008.420 ;
        RECT 2535.590 3008.360 2535.910 3008.420 ;
        RECT 2535.590 1966.460 2535.910 1966.520 ;
        RECT 2900.830 1966.460 2901.150 1966.520 ;
        RECT 2535.590 1966.320 2901.150 1966.460 ;
        RECT 2535.590 1966.260 2535.910 1966.320 ;
        RECT 2900.830 1966.260 2901.150 1966.320 ;
      LAYER via ;
        RECT 593.040 3008.360 593.300 3008.620 ;
        RECT 2535.620 3008.360 2535.880 3008.620 ;
        RECT 2535.620 1966.260 2535.880 1966.520 ;
        RECT 2900.860 1966.260 2901.120 1966.520 ;
      LAYER met2 ;
        RECT 592.250 3008.730 592.530 3010.000 ;
        RECT 592.250 3008.650 593.240 3008.730 ;
        RECT 592.250 3008.590 593.300 3008.650 ;
        RECT 592.250 3006.000 592.530 3008.590 ;
        RECT 593.040 3008.330 593.300 3008.590 ;
        RECT 2535.620 3008.330 2535.880 3008.650 ;
        RECT 2535.680 1966.550 2535.820 3008.330 ;
        RECT 2535.620 1966.230 2535.880 1966.550 ;
        RECT 2900.860 1966.230 2901.120 1966.550 ;
        RECT 2900.920 1965.045 2901.060 1966.230 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 864.410 3022.840 864.730 3022.900 ;
        RECT 2570.550 3022.840 2570.870 3022.900 ;
        RECT 864.410 3022.700 2570.870 3022.840 ;
        RECT 864.410 3022.640 864.730 3022.700 ;
        RECT 2570.550 3022.640 2570.870 3022.700 ;
        RECT 2570.550 2201.060 2570.870 2201.120 ;
        RECT 2898.070 2201.060 2898.390 2201.120 ;
        RECT 2570.550 2200.920 2898.390 2201.060 ;
        RECT 2570.550 2200.860 2570.870 2200.920 ;
        RECT 2898.070 2200.860 2898.390 2200.920 ;
      LAYER via ;
        RECT 864.440 3022.640 864.700 3022.900 ;
        RECT 2570.580 3022.640 2570.840 3022.900 ;
        RECT 2570.580 2200.860 2570.840 2201.120 ;
        RECT 2898.100 2200.860 2898.360 2201.120 ;
      LAYER met2 ;
        RECT 864.440 3022.610 864.700 3022.930 ;
        RECT 2570.580 3022.610 2570.840 3022.930 ;
        RECT 864.500 3010.000 864.640 3022.610 ;
        RECT 864.500 3009.340 864.850 3010.000 ;
        RECT 864.570 3006.000 864.850 3009.340 ;
        RECT 2570.640 2201.150 2570.780 3022.610 ;
        RECT 2570.580 2200.830 2570.840 2201.150 ;
        RECT 2898.100 2200.830 2898.360 2201.150 ;
        RECT 2898.160 2199.645 2898.300 2200.830 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
      LAYER via2 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
      LAYER met3 ;
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1925.320 2519.810 1925.380 ;
        RECT 2749.490 1925.320 2749.810 1925.380 ;
        RECT 2519.490 1925.180 2749.810 1925.320 ;
        RECT 2519.490 1925.120 2519.810 1925.180 ;
        RECT 2749.490 1925.120 2749.810 1925.180 ;
        RECT 2749.490 206.960 2749.810 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2749.490 206.820 2901.150 206.960 ;
        RECT 2749.490 206.760 2749.810 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2519.520 1925.120 2519.780 1925.380 ;
        RECT 2749.520 1925.120 2749.780 1925.380 ;
        RECT 2749.520 206.760 2749.780 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2519.510 1927.275 2519.790 1927.645 ;
        RECT 2519.580 1925.410 2519.720 1927.275 ;
        RECT 2519.520 1925.090 2519.780 1925.410 ;
        RECT 2749.520 1925.090 2749.780 1925.410 ;
        RECT 2749.580 207.050 2749.720 1925.090 ;
        RECT 2749.520 206.730 2749.780 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2519.510 1927.320 2519.790 1927.600 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2506.000 1927.610 2510.000 1927.760 ;
        RECT 2519.485 1927.610 2519.815 1927.625 ;
        RECT 2506.000 1927.310 2519.815 1927.610 ;
        RECT 2506.000 1927.160 2510.000 1927.310 ;
        RECT 2519.485 1927.295 2519.815 1927.310 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2708.340 2519.810 2708.400 ;
        RECT 2825.390 2708.340 2825.710 2708.400 ;
        RECT 2519.490 2708.200 2825.710 2708.340 ;
        RECT 2519.490 2708.140 2519.810 2708.200 ;
        RECT 2825.390 2708.140 2825.710 2708.200 ;
        RECT 2825.390 2552.960 2825.710 2553.020 ;
        RECT 2900.830 2552.960 2901.150 2553.020 ;
        RECT 2825.390 2552.820 2901.150 2552.960 ;
        RECT 2825.390 2552.760 2825.710 2552.820 ;
        RECT 2900.830 2552.760 2901.150 2552.820 ;
      LAYER via ;
        RECT 2519.520 2708.140 2519.780 2708.400 ;
        RECT 2825.420 2708.140 2825.680 2708.400 ;
        RECT 2825.420 2552.760 2825.680 2553.020 ;
        RECT 2900.860 2552.760 2901.120 2553.020 ;
      LAYER met2 ;
        RECT 2519.510 2713.355 2519.790 2713.725 ;
        RECT 2519.580 2708.430 2519.720 2713.355 ;
        RECT 2519.520 2708.110 2519.780 2708.430 ;
        RECT 2825.420 2708.110 2825.680 2708.430 ;
        RECT 2825.480 2553.050 2825.620 2708.110 ;
        RECT 2825.420 2552.730 2825.680 2553.050 ;
        RECT 2900.860 2552.730 2901.120 2553.050 ;
        RECT 2900.920 2551.885 2901.060 2552.730 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
      LAYER via2 ;
        RECT 2519.510 2713.400 2519.790 2713.680 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
      LAYER met3 ;
        RECT 2506.000 2713.690 2510.000 2713.840 ;
        RECT 2519.485 2713.690 2519.815 2713.705 ;
        RECT 2506.000 2713.390 2519.815 2713.690 ;
        RECT 2506.000 2713.240 2510.000 2713.390 ;
        RECT 2519.485 2713.375 2519.815 2713.390 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2846.550 2781.100 2846.870 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2846.550 2780.960 2901.150 2781.100 ;
        RECT 2846.550 2780.900 2846.870 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2520.410 1676.440 2520.730 1676.500 ;
        RECT 2846.550 1676.440 2846.870 1676.500 ;
        RECT 2520.410 1676.300 2846.870 1676.440 ;
        RECT 2520.410 1676.240 2520.730 1676.300 ;
        RECT 2846.550 1676.240 2846.870 1676.300 ;
      LAYER via ;
        RECT 2846.580 2780.900 2846.840 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2520.440 1676.240 2520.700 1676.500 ;
        RECT 2846.580 1676.240 2846.840 1676.500 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2846.580 2780.870 2846.840 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2846.640 1676.530 2846.780 2780.870 ;
        RECT 2520.440 1676.210 2520.700 1676.530 ;
        RECT 2846.580 1676.210 2846.840 1676.530 ;
        RECT 2520.500 1671.965 2520.640 1676.210 ;
        RECT 2520.430 1671.595 2520.710 1671.965 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2520.430 1671.640 2520.710 1671.920 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2506.000 1671.930 2510.000 1672.080 ;
        RECT 2520.405 1671.930 2520.735 1671.945 ;
        RECT 2506.000 1671.630 2520.735 1671.930 ;
        RECT 2506.000 1671.480 2510.000 1671.630 ;
        RECT 2520.405 1671.615 2520.735 1671.630 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.070 3020.460 1449.390 3020.520 ;
        RECT 1496.910 3020.460 1497.230 3020.520 ;
        RECT 1449.070 3020.320 1497.230 3020.460 ;
        RECT 1449.070 3020.260 1449.390 3020.320 ;
        RECT 1496.910 3020.260 1497.230 3020.320 ;
        RECT 1642.270 3020.460 1642.590 3020.520 ;
        RECT 1690.110 3020.460 1690.430 3020.520 ;
        RECT 1642.270 3020.320 1690.430 3020.460 ;
        RECT 1642.270 3020.260 1642.590 3020.320 ;
        RECT 1690.110 3020.260 1690.430 3020.320 ;
        RECT 1738.870 3020.460 1739.190 3020.520 ;
        RECT 1786.710 3020.460 1787.030 3020.520 ;
        RECT 1738.870 3020.320 1787.030 3020.460 ;
        RECT 1738.870 3020.260 1739.190 3020.320 ;
        RECT 1786.710 3020.260 1787.030 3020.320 ;
        RECT 2415.070 3019.440 2415.390 3019.500 ;
        RECT 2463.830 3019.440 2464.150 3019.500 ;
        RECT 2415.070 3019.300 2464.150 3019.440 ;
        RECT 2415.070 3019.240 2415.390 3019.300 ;
        RECT 2463.830 3019.240 2464.150 3019.300 ;
        RECT 2222.330 3018.760 2222.650 3018.820 ;
        RECT 2245.790 3018.760 2246.110 3018.820 ;
        RECT 2222.330 3018.620 2246.110 3018.760 ;
        RECT 2222.330 3018.560 2222.650 3018.620 ;
        RECT 2245.790 3018.560 2246.110 3018.620 ;
        RECT 2584.350 3018.760 2584.670 3018.820 ;
        RECT 2628.510 3018.760 2628.830 3018.820 ;
        RECT 2584.350 3018.620 2628.830 3018.760 ;
        RECT 2584.350 3018.560 2584.670 3018.620 ;
        RECT 2628.510 3018.560 2628.830 3018.620 ;
        RECT 1546.130 3018.420 1546.450 3018.480 ;
        RECT 1593.510 3018.420 1593.830 3018.480 ;
        RECT 1546.130 3018.280 1593.830 3018.420 ;
        RECT 1546.130 3018.220 1546.450 3018.280 ;
        RECT 1593.510 3018.220 1593.830 3018.280 ;
        RECT 2669.910 3018.420 2670.230 3018.480 ;
        RECT 2704.410 3018.420 2704.730 3018.480 ;
        RECT 2669.910 3018.280 2704.730 3018.420 ;
        RECT 2669.910 3018.220 2670.230 3018.280 ;
        RECT 2704.410 3018.220 2704.730 3018.280 ;
        RECT 335.410 1248.720 335.730 1248.780 ;
        RECT 393.370 1248.720 393.690 1248.780 ;
        RECT 335.410 1248.580 393.690 1248.720 ;
        RECT 335.410 1248.520 335.730 1248.580 ;
        RECT 393.370 1248.520 393.690 1248.580 ;
      LAYER via ;
        RECT 1449.100 3020.260 1449.360 3020.520 ;
        RECT 1496.940 3020.260 1497.200 3020.520 ;
        RECT 1642.300 3020.260 1642.560 3020.520 ;
        RECT 1690.140 3020.260 1690.400 3020.520 ;
        RECT 1738.900 3020.260 1739.160 3020.520 ;
        RECT 1786.740 3020.260 1787.000 3020.520 ;
        RECT 2415.100 3019.240 2415.360 3019.500 ;
        RECT 2463.860 3019.240 2464.120 3019.500 ;
        RECT 2222.360 3018.560 2222.620 3018.820 ;
        RECT 2245.820 3018.560 2246.080 3018.820 ;
        RECT 2584.380 3018.560 2584.640 3018.820 ;
        RECT 2628.540 3018.560 2628.800 3018.820 ;
        RECT 1546.160 3018.220 1546.420 3018.480 ;
        RECT 1593.540 3018.220 1593.800 3018.480 ;
        RECT 2669.940 3018.220 2670.200 3018.480 ;
        RECT 2704.440 3018.220 2704.700 3018.480 ;
        RECT 335.440 1248.520 335.700 1248.780 ;
        RECT 393.400 1248.520 393.660 1248.780 ;
      LAYER met2 ;
        RECT 1545.760 3020.830 1546.360 3020.970 ;
        RECT 1449.100 3020.405 1449.360 3020.550 ;
        RECT 335.430 3020.035 335.710 3020.405 ;
        RECT 980.350 3020.035 980.630 3020.405 ;
        RECT 1449.090 3020.035 1449.370 3020.405 ;
        RECT 1496.940 3020.230 1497.200 3020.550 ;
        RECT 1545.760 3020.405 1545.900 3020.830 ;
        RECT 335.500 1248.810 335.640 3020.035 ;
        RECT 593.950 3019.610 594.230 3019.725 ;
        RECT 593.100 3019.470 594.230 3019.610 ;
        RECT 593.100 3019.045 593.240 3019.470 ;
        RECT 593.950 3019.355 594.230 3019.470 ;
        RECT 690.550 3019.355 690.830 3019.725 ;
        RECT 748.050 3019.610 748.330 3019.725 ;
        RECT 748.050 3019.470 748.720 3019.610 ;
        RECT 748.050 3019.355 748.330 3019.470 ;
        RECT 593.030 3018.675 593.310 3019.045 ;
        RECT 689.630 3018.930 689.910 3019.045 ;
        RECT 690.620 3018.930 690.760 3019.355 ;
        RECT 748.580 3019.045 748.720 3019.470 ;
        RECT 689.630 3018.790 690.760 3018.930 ;
        RECT 689.630 3018.675 689.910 3018.790 ;
        RECT 748.510 3018.675 748.790 3019.045 ;
        RECT 979.430 3018.930 979.710 3019.045 ;
        RECT 980.420 3018.930 980.560 3020.035 ;
        RECT 1497.000 3019.045 1497.140 3020.230 ;
        RECT 1545.690 3020.035 1545.970 3020.405 ;
        RECT 979.430 3018.790 980.560 3018.930 ;
        RECT 979.430 3018.675 979.710 3018.790 ;
        RECT 1496.930 3018.675 1497.210 3019.045 ;
        RECT 1546.220 3018.510 1546.360 3020.830 ;
        RECT 2318.030 3020.715 2318.310 3021.085 ;
        RECT 1642.300 3020.405 1642.560 3020.550 ;
        RECT 1642.290 3020.035 1642.570 3020.405 ;
        RECT 1690.140 3020.230 1690.400 3020.550 ;
        RECT 1738.900 3020.405 1739.160 3020.550 ;
        RECT 1690.200 3019.045 1690.340 3020.230 ;
        RECT 1738.890 3020.035 1739.170 3020.405 ;
        RECT 1786.740 3020.230 1787.000 3020.550 ;
        RECT 1786.800 3019.725 1786.940 3020.230 ;
        RECT 2318.100 3019.725 2318.240 3020.715 ;
        RECT 1786.730 3019.355 1787.010 3019.725 ;
        RECT 2318.030 3019.355 2318.310 3019.725 ;
        RECT 2415.090 3019.355 2415.370 3019.725 ;
        RECT 2463.850 3019.355 2464.130 3019.725 ;
        RECT 2584.370 3019.355 2584.650 3019.725 ;
        RECT 2415.100 3019.210 2415.360 3019.355 ;
        RECT 2463.860 3019.210 2464.120 3019.355 ;
        RECT 1593.530 3018.675 1593.810 3019.045 ;
        RECT 1690.130 3018.675 1690.410 3019.045 ;
        RECT 1848.370 3018.930 1848.650 3019.045 ;
        RECT 1849.750 3018.930 1850.030 3019.045 ;
        RECT 1848.370 3018.790 1850.030 3018.930 ;
        RECT 1848.370 3018.675 1848.650 3018.790 ;
        RECT 1849.750 3018.675 1850.030 3018.790 ;
        RECT 1897.130 3018.675 1897.410 3019.045 ;
        RECT 1593.600 3018.510 1593.740 3018.675 ;
        RECT 1546.160 3018.190 1546.420 3018.510 ;
        RECT 1593.540 3018.190 1593.800 3018.510 ;
        RECT 1897.200 3018.250 1897.340 3018.675 ;
        RECT 2222.360 3018.530 2222.620 3018.850 ;
        RECT 2245.810 3018.675 2246.090 3019.045 ;
        RECT 2366.330 3018.675 2366.610 3019.045 ;
        RECT 2584.440 3018.850 2584.580 3019.355 ;
        RECT 2245.820 3018.530 2246.080 3018.675 ;
        RECT 1898.050 3018.250 1898.330 3018.365 ;
        RECT 1897.200 3018.110 1898.330 3018.250 ;
        RECT 1898.050 3017.995 1898.330 3018.110 ;
        RECT 2221.890 3017.995 2222.170 3018.365 ;
        RECT 2221.960 3017.570 2222.100 3017.995 ;
        RECT 2222.420 3017.570 2222.560 3018.530 ;
        RECT 2366.400 3018.365 2366.540 3018.675 ;
        RECT 2584.380 3018.530 2584.640 3018.850 ;
        RECT 2628.540 3018.530 2628.800 3018.850 ;
        RECT 2704.430 3018.675 2704.710 3019.045 ;
        RECT 2863.130 3018.930 2863.410 3019.045 ;
        RECT 2864.050 3018.930 2864.330 3019.045 ;
        RECT 2863.130 3018.790 2864.330 3018.930 ;
        RECT 2863.130 3018.675 2863.410 3018.790 ;
        RECT 2864.050 3018.675 2864.330 3018.790 ;
        RECT 2628.600 3018.365 2628.740 3018.530 ;
        RECT 2704.500 3018.510 2704.640 3018.675 ;
        RECT 2669.940 3018.365 2670.200 3018.510 ;
        RECT 2366.330 3017.995 2366.610 3018.365 ;
        RECT 2628.530 3017.995 2628.810 3018.365 ;
        RECT 2669.930 3017.995 2670.210 3018.365 ;
        RECT 2704.440 3018.190 2704.700 3018.510 ;
        RECT 2221.960 3017.430 2222.560 3017.570 ;
        RECT 335.440 1248.490 335.700 1248.810 ;
        RECT 393.400 1248.490 393.660 1248.810 ;
        RECT 393.460 1244.925 393.600 1248.490 ;
        RECT 393.390 1244.555 393.670 1244.925 ;
      LAYER via2 ;
        RECT 335.430 3020.080 335.710 3020.360 ;
        RECT 980.350 3020.080 980.630 3020.360 ;
        RECT 1449.090 3020.080 1449.370 3020.360 ;
        RECT 593.950 3019.400 594.230 3019.680 ;
        RECT 690.550 3019.400 690.830 3019.680 ;
        RECT 748.050 3019.400 748.330 3019.680 ;
        RECT 593.030 3018.720 593.310 3019.000 ;
        RECT 689.630 3018.720 689.910 3019.000 ;
        RECT 748.510 3018.720 748.790 3019.000 ;
        RECT 979.430 3018.720 979.710 3019.000 ;
        RECT 1545.690 3020.080 1545.970 3020.360 ;
        RECT 1496.930 3018.720 1497.210 3019.000 ;
        RECT 2318.030 3020.760 2318.310 3021.040 ;
        RECT 1642.290 3020.080 1642.570 3020.360 ;
        RECT 1738.890 3020.080 1739.170 3020.360 ;
        RECT 1786.730 3019.400 1787.010 3019.680 ;
        RECT 2318.030 3019.400 2318.310 3019.680 ;
        RECT 2415.090 3019.400 2415.370 3019.680 ;
        RECT 2463.850 3019.400 2464.130 3019.680 ;
        RECT 2584.370 3019.400 2584.650 3019.680 ;
        RECT 1593.530 3018.720 1593.810 3019.000 ;
        RECT 1690.130 3018.720 1690.410 3019.000 ;
        RECT 1848.370 3018.720 1848.650 3019.000 ;
        RECT 1849.750 3018.720 1850.030 3019.000 ;
        RECT 1897.130 3018.720 1897.410 3019.000 ;
        RECT 2245.810 3018.720 2246.090 3019.000 ;
        RECT 2366.330 3018.720 2366.610 3019.000 ;
        RECT 1898.050 3018.040 1898.330 3018.320 ;
        RECT 2221.890 3018.040 2222.170 3018.320 ;
        RECT 2704.430 3018.720 2704.710 3019.000 ;
        RECT 2863.130 3018.720 2863.410 3019.000 ;
        RECT 2864.050 3018.720 2864.330 3019.000 ;
        RECT 2366.330 3018.040 2366.610 3018.320 ;
        RECT 2628.530 3018.040 2628.810 3018.320 ;
        RECT 2669.930 3018.040 2670.210 3018.320 ;
        RECT 393.390 1244.600 393.670 1244.880 ;
      LAYER met3 ;
        RECT 2269.910 3021.050 2270.290 3021.060 ;
        RECT 2318.005 3021.050 2318.335 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2269.910 3020.750 2318.335 3021.050 ;
        RECT 2269.910 3020.740 2270.290 3020.750 ;
        RECT 2318.005 3020.735 2318.335 3020.750 ;
        RECT 2916.710 3020.750 2924.800 3021.050 ;
        RECT 335.405 3020.370 335.735 3020.385 ;
        RECT 434.510 3020.370 434.890 3020.380 ;
        RECT 765.710 3020.370 766.090 3020.380 ;
        RECT 980.325 3020.370 980.655 3020.385 ;
        RECT 1449.065 3020.370 1449.395 3020.385 ;
        RECT 1545.665 3020.370 1545.995 3020.385 ;
        RECT 1642.265 3020.370 1642.595 3020.385 ;
        RECT 1738.865 3020.370 1739.195 3020.385 ;
        RECT 335.405 3020.070 352.970 3020.370 ;
        RECT 335.405 3020.055 335.735 3020.070 ;
        RECT 352.670 3019.690 352.970 3020.070 ;
        RECT 434.510 3020.070 436.690 3020.370 ;
        RECT 434.510 3020.060 434.890 3020.070 ;
        RECT 436.390 3019.690 436.690 3020.070 ;
        RECT 499.870 3020.070 546.170 3020.370 ;
        RECT 499.870 3019.690 500.170 3020.070 ;
        RECT 352.670 3019.390 379.650 3019.690 ;
        RECT 436.390 3019.390 500.170 3019.690 ;
        RECT 379.350 3019.180 379.650 3019.390 ;
        RECT 379.350 3019.010 380.570 3019.180 ;
        RECT 434.510 3019.010 434.890 3019.020 ;
        RECT 379.350 3018.880 434.890 3019.010 ;
        RECT 380.270 3018.710 434.890 3018.880 ;
        RECT 545.870 3019.010 546.170 3020.070 ;
        RECT 765.710 3020.070 790.890 3020.370 ;
        RECT 765.710 3020.060 766.090 3020.070 ;
        RECT 593.925 3019.690 594.255 3019.705 ;
        RECT 690.525 3019.690 690.855 3019.705 ;
        RECT 748.025 3019.690 748.355 3019.705 ;
        RECT 593.925 3019.390 645.530 3019.690 ;
        RECT 593.925 3019.375 594.255 3019.390 ;
        RECT 593.005 3019.010 593.335 3019.025 ;
        RECT 545.870 3018.710 593.335 3019.010 ;
        RECT 645.230 3019.010 645.530 3019.390 ;
        RECT 690.525 3019.390 748.355 3019.690 ;
        RECT 790.590 3019.690 790.890 3020.070 ;
        RECT 861.430 3020.070 932.570 3020.370 ;
        RECT 861.430 3019.690 861.730 3020.070 ;
        RECT 790.590 3019.390 861.730 3019.690 ;
        RECT 690.525 3019.375 690.855 3019.390 ;
        RECT 748.025 3019.375 748.355 3019.390 ;
        RECT 689.605 3019.010 689.935 3019.025 ;
        RECT 645.230 3018.710 689.935 3019.010 ;
        RECT 434.510 3018.700 434.890 3018.710 ;
        RECT 593.005 3018.695 593.335 3018.710 ;
        RECT 689.605 3018.695 689.935 3018.710 ;
        RECT 748.485 3019.010 748.815 3019.025 ;
        RECT 765.710 3019.010 766.090 3019.020 ;
        RECT 748.485 3018.710 766.090 3019.010 ;
        RECT 932.270 3019.010 932.570 3020.070 ;
        RECT 980.325 3020.070 1029.170 3020.370 ;
        RECT 980.325 3020.055 980.655 3020.070 ;
        RECT 979.405 3019.010 979.735 3019.025 ;
        RECT 932.270 3018.710 979.735 3019.010 ;
        RECT 1028.870 3019.010 1029.170 3020.070 ;
        RECT 1075.790 3020.070 1125.770 3020.370 ;
        RECT 1075.790 3019.010 1076.090 3020.070 ;
        RECT 1028.870 3018.710 1076.090 3019.010 ;
        RECT 1125.470 3019.010 1125.770 3020.070 ;
        RECT 1172.390 3020.070 1222.370 3020.370 ;
        RECT 1172.390 3019.010 1172.690 3020.070 ;
        RECT 1125.470 3018.710 1172.690 3019.010 ;
        RECT 1222.070 3019.010 1222.370 3020.070 ;
        RECT 1268.990 3020.070 1318.970 3020.370 ;
        RECT 1268.990 3019.010 1269.290 3020.070 ;
        RECT 1222.070 3018.710 1269.290 3019.010 ;
        RECT 1318.670 3019.010 1318.970 3020.070 ;
        RECT 1414.350 3020.070 1449.395 3020.370 ;
        RECT 1414.350 3019.010 1414.650 3020.070 ;
        RECT 1449.065 3020.055 1449.395 3020.070 ;
        RECT 1510.950 3020.070 1545.995 3020.370 ;
        RECT 1318.670 3018.710 1414.650 3019.010 ;
        RECT 1496.905 3019.010 1497.235 3019.025 ;
        RECT 1510.950 3019.010 1511.250 3020.070 ;
        RECT 1545.665 3020.055 1545.995 3020.070 ;
        RECT 1607.550 3020.070 1642.595 3020.370 ;
        RECT 1496.905 3018.710 1511.250 3019.010 ;
        RECT 1593.505 3019.010 1593.835 3019.025 ;
        RECT 1607.550 3019.010 1607.850 3020.070 ;
        RECT 1642.265 3020.055 1642.595 3020.070 ;
        RECT 1704.150 3020.070 1739.195 3020.370 ;
        RECT 1593.505 3018.710 1607.850 3019.010 ;
        RECT 1690.105 3019.010 1690.435 3019.025 ;
        RECT 1704.150 3019.010 1704.450 3020.070 ;
        RECT 1738.865 3020.055 1739.195 3020.070 ;
        RECT 2766.750 3020.070 2815.810 3020.370 ;
        RECT 1786.705 3019.690 1787.035 3019.705 ;
        RECT 1924.910 3019.690 1925.290 3019.700 ;
        RECT 2318.005 3019.690 2318.335 3019.705 ;
        RECT 2415.065 3019.690 2415.395 3019.705 ;
        RECT 1786.705 3019.390 1801.050 3019.690 ;
        RECT 1786.705 3019.375 1787.035 3019.390 ;
        RECT 1690.105 3018.710 1704.450 3019.010 ;
        RECT 1800.750 3019.010 1801.050 3019.390 ;
        RECT 1924.910 3019.390 1995.170 3019.690 ;
        RECT 1924.910 3019.380 1925.290 3019.390 ;
        RECT 1848.345 3019.010 1848.675 3019.025 ;
        RECT 1800.750 3018.710 1848.675 3019.010 ;
        RECT 748.485 3018.695 748.815 3018.710 ;
        RECT 765.710 3018.700 766.090 3018.710 ;
        RECT 979.405 3018.695 979.735 3018.710 ;
        RECT 1496.905 3018.695 1497.235 3018.710 ;
        RECT 1593.505 3018.695 1593.835 3018.710 ;
        RECT 1690.105 3018.695 1690.435 3018.710 ;
        RECT 1848.345 3018.695 1848.675 3018.710 ;
        RECT 1849.725 3019.010 1850.055 3019.025 ;
        RECT 1897.105 3019.010 1897.435 3019.025 ;
        RECT 1849.725 3018.710 1897.435 3019.010 ;
        RECT 1849.725 3018.695 1850.055 3018.710 ;
        RECT 1897.105 3018.695 1897.435 3018.710 ;
        RECT 1898.025 3018.330 1898.355 3018.345 ;
        RECT 1924.910 3018.330 1925.290 3018.340 ;
        RECT 1898.025 3018.030 1925.290 3018.330 ;
        RECT 1994.870 3018.330 1995.170 3019.390 ;
        RECT 2022.470 3019.390 2188.370 3019.690 ;
        RECT 2022.470 3019.010 2022.770 3019.390 ;
        RECT 2021.550 3018.710 2022.770 3019.010 ;
        RECT 2021.550 3018.330 2021.850 3018.710 ;
        RECT 1994.870 3018.030 2021.850 3018.330 ;
        RECT 2188.070 3018.330 2188.370 3019.390 ;
        RECT 2318.005 3019.390 2330.970 3019.690 ;
        RECT 2318.005 3019.375 2318.335 3019.390 ;
        RECT 2245.785 3019.010 2246.115 3019.025 ;
        RECT 2269.910 3019.010 2270.290 3019.020 ;
        RECT 2245.785 3018.710 2270.290 3019.010 ;
        RECT 2330.670 3019.010 2330.970 3019.390 ;
        RECT 2381.270 3019.390 2415.395 3019.690 ;
        RECT 2366.305 3019.010 2366.635 3019.025 ;
        RECT 2381.270 3019.010 2381.570 3019.390 ;
        RECT 2415.065 3019.375 2415.395 3019.390 ;
        RECT 2463.825 3019.690 2464.155 3019.705 ;
        RECT 2584.345 3019.690 2584.675 3019.705 ;
        RECT 2463.825 3019.390 2584.675 3019.690 ;
        RECT 2463.825 3019.375 2464.155 3019.390 ;
        RECT 2584.345 3019.375 2584.675 3019.390 ;
        RECT 2330.670 3018.710 2366.635 3019.010 ;
        RECT 2245.785 3018.695 2246.115 3018.710 ;
        RECT 2269.910 3018.700 2270.290 3018.710 ;
        RECT 2366.305 3018.695 2366.635 3018.710 ;
        RECT 2380.350 3018.710 2381.570 3019.010 ;
        RECT 2704.405 3019.010 2704.735 3019.025 ;
        RECT 2766.750 3019.010 2767.050 3020.070 ;
        RECT 2704.405 3018.710 2767.050 3019.010 ;
        RECT 2815.510 3019.010 2815.810 3020.070 ;
        RECT 2916.710 3019.690 2917.010 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2911.190 3019.390 2917.010 3019.690 ;
        RECT 2863.105 3019.010 2863.435 3019.025 ;
        RECT 2815.510 3018.710 2863.435 3019.010 ;
        RECT 2221.865 3018.330 2222.195 3018.345 ;
        RECT 2188.070 3018.030 2222.195 3018.330 ;
        RECT 1898.025 3018.015 1898.355 3018.030 ;
        RECT 1924.910 3018.020 1925.290 3018.030 ;
        RECT 2221.865 3018.015 2222.195 3018.030 ;
        RECT 2366.305 3018.330 2366.635 3018.345 ;
        RECT 2380.350 3018.330 2380.650 3018.710 ;
        RECT 2704.405 3018.695 2704.735 3018.710 ;
        RECT 2863.105 3018.695 2863.435 3018.710 ;
        RECT 2864.025 3019.010 2864.355 3019.025 ;
        RECT 2911.190 3019.010 2911.490 3019.390 ;
        RECT 2864.025 3018.710 2911.490 3019.010 ;
        RECT 2864.025 3018.695 2864.355 3018.710 ;
        RECT 2366.305 3018.030 2380.650 3018.330 ;
        RECT 2628.505 3018.330 2628.835 3018.345 ;
        RECT 2669.905 3018.330 2670.235 3018.345 ;
        RECT 2628.505 3018.030 2670.235 3018.330 ;
        RECT 2366.305 3018.015 2366.635 3018.030 ;
        RECT 2628.505 3018.015 2628.835 3018.030 ;
        RECT 2669.905 3018.015 2670.235 3018.030 ;
        RECT 393.365 1244.890 393.695 1244.905 ;
        RECT 410.000 1244.890 414.000 1245.040 ;
        RECT 393.365 1244.590 414.000 1244.890 ;
        RECT 393.365 1244.575 393.695 1244.590 ;
        RECT 410.000 1244.440 414.000 1244.590 ;
      LAYER via3 ;
        RECT 2269.940 3020.740 2270.260 3021.060 ;
        RECT 434.540 3020.060 434.860 3020.380 ;
        RECT 434.540 3018.700 434.860 3019.020 ;
        RECT 765.740 3020.060 766.060 3020.380 ;
        RECT 765.740 3018.700 766.060 3019.020 ;
        RECT 1924.940 3019.380 1925.260 3019.700 ;
        RECT 1924.940 3018.020 1925.260 3018.340 ;
        RECT 2269.940 3018.700 2270.260 3019.020 ;
      LAYER met4 ;
        RECT 2269.935 3020.735 2270.265 3021.065 ;
        RECT 434.535 3020.055 434.865 3020.385 ;
        RECT 765.735 3020.055 766.065 3020.385 ;
        RECT 434.550 3019.025 434.850 3020.055 ;
        RECT 765.750 3019.025 766.050 3020.055 ;
        RECT 1924.935 3019.375 1925.265 3019.705 ;
        RECT 434.535 3018.695 434.865 3019.025 ;
        RECT 765.735 3018.695 766.065 3019.025 ;
        RECT 1924.950 3018.345 1925.250 3019.375 ;
        RECT 2269.950 3019.025 2270.250 3020.735 ;
        RECT 2269.935 3018.695 2270.265 3019.025 ;
        RECT 1924.935 3018.015 1925.265 3018.345 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 889.710 3250.300 890.030 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 889.710 3250.160 2901.150 3250.300 ;
        RECT 889.710 3250.100 890.030 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 889.740 3250.100 890.000 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 889.740 3250.070 890.000 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 888.490 3009.410 888.770 3010.000 ;
        RECT 889.800 3009.410 889.940 3250.070 ;
        RECT 888.490 3009.270 889.940 3009.410 ;
        RECT 888.490 3006.000 888.770 3009.270 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 807.530 510.340 807.810 514.000 ;
        RECT 807.460 510.000 807.810 510.340 ;
        RECT 807.460 489.445 807.600 510.000 ;
        RECT 807.390 489.075 807.670 489.445 ;
      LAYER via2 ;
        RECT 807.390 489.120 807.670 489.400 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2916.710 3489.950 2924.800 3490.250 ;
        RECT 2597.430 3486.170 2597.810 3486.180 ;
        RECT 2597.430 3485.870 2642.850 3486.170 ;
        RECT 2597.430 3485.860 2597.810 3485.870 ;
        RECT 2642.550 3485.490 2642.850 3485.870 ;
        RECT 2691.310 3485.870 2739.450 3486.170 ;
        RECT 2642.550 3485.190 2690.690 3485.490 ;
        RECT 2690.390 3484.810 2690.690 3485.190 ;
        RECT 2691.310 3484.810 2691.610 3485.870 ;
        RECT 2739.150 3485.490 2739.450 3485.870 ;
        RECT 2787.910 3485.870 2836.050 3486.170 ;
        RECT 2739.150 3485.190 2787.290 3485.490 ;
        RECT 2690.390 3484.510 2691.610 3484.810 ;
        RECT 2786.990 3484.810 2787.290 3485.190 ;
        RECT 2787.910 3484.810 2788.210 3485.870 ;
        RECT 2835.750 3485.490 2836.050 3485.870 ;
        RECT 2835.750 3485.190 2883.890 3485.490 ;
        RECT 2786.990 3484.510 2788.210 3484.810 ;
        RECT 2883.590 3484.810 2883.890 3485.190 ;
        RECT 2916.710 3484.810 2917.010 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2883.590 3484.510 2917.010 3484.810 ;
        RECT 807.365 489.410 807.695 489.425 ;
        RECT 2597.430 489.410 2597.810 489.420 ;
        RECT 807.365 489.110 2597.810 489.410 ;
        RECT 807.365 489.095 807.695 489.110 ;
        RECT 2597.430 489.100 2597.810 489.110 ;
      LAYER via3 ;
        RECT 2597.460 3485.860 2597.780 3486.180 ;
        RECT 2597.460 489.100 2597.780 489.420 ;
      LAYER met4 ;
        RECT 2597.455 3485.855 2597.785 3486.185 ;
        RECT 2597.470 489.425 2597.770 3485.855 ;
        RECT 2597.455 489.095 2597.785 489.425 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2546.170 859.080 2546.490 859.140 ;
        RECT 2635.870 859.080 2636.190 859.140 ;
        RECT 2546.170 858.940 2636.190 859.080 ;
        RECT 2546.170 858.880 2546.490 858.940 ;
        RECT 2635.870 858.880 2636.190 858.940 ;
        RECT 2518.570 853.980 2518.890 854.040 ;
        RECT 2546.170 853.980 2546.490 854.040 ;
        RECT 2518.570 853.840 2546.490 853.980 ;
        RECT 2518.570 853.780 2518.890 853.840 ;
        RECT 2546.170 853.780 2546.490 853.840 ;
      LAYER via ;
        RECT 2546.200 858.880 2546.460 859.140 ;
        RECT 2635.900 858.880 2636.160 859.140 ;
        RECT 2518.600 853.780 2518.860 854.040 ;
        RECT 2546.200 853.780 2546.460 854.040 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 859.170 2636.100 3517.600 ;
        RECT 2546.200 858.850 2546.460 859.170 ;
        RECT 2635.900 858.850 2636.160 859.170 ;
        RECT 2546.260 854.070 2546.400 858.850 ;
        RECT 2518.600 853.750 2518.860 854.070 ;
        RECT 2546.200 853.750 2546.460 854.070 ;
        RECT 2518.660 850.525 2518.800 853.750 ;
        RECT 2518.590 850.155 2518.870 850.525 ;
      LAYER via2 ;
        RECT 2518.590 850.200 2518.870 850.480 ;
      LAYER met3 ;
        RECT 2506.000 850.490 2510.000 850.640 ;
        RECT 2518.565 850.490 2518.895 850.505 ;
        RECT 2506.000 850.190 2518.895 850.490 ;
        RECT 2506.000 850.040 2510.000 850.190 ;
        RECT 2518.565 850.175 2518.895 850.190 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 343.690 3501.560 344.010 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 343.690 3501.420 2311.890 3501.560 ;
        RECT 343.690 3501.360 344.010 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
        RECT 343.690 1117.480 344.010 1117.540 ;
        RECT 393.370 1117.480 393.690 1117.540 ;
        RECT 343.690 1117.340 393.690 1117.480 ;
        RECT 343.690 1117.280 344.010 1117.340 ;
        RECT 393.370 1117.280 393.690 1117.340 ;
      LAYER via ;
        RECT 343.720 3501.360 343.980 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
        RECT 343.720 1117.280 343.980 1117.540 ;
        RECT 393.400 1117.280 393.660 1117.540 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 343.720 3501.330 343.980 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 343.780 1117.570 343.920 3501.330 ;
        RECT 343.720 1117.250 343.980 1117.570 ;
        RECT 393.400 1117.250 393.660 1117.570 ;
        RECT 393.460 1117.085 393.600 1117.250 ;
        RECT 393.390 1116.715 393.670 1117.085 ;
      LAYER via2 ;
        RECT 393.390 1116.760 393.670 1117.040 ;
      LAYER met3 ;
        RECT 393.365 1117.050 393.695 1117.065 ;
        RECT 410.000 1117.050 414.000 1117.200 ;
        RECT 393.365 1116.750 414.000 1117.050 ;
        RECT 393.365 1116.735 393.695 1116.750 ;
        RECT 410.000 1116.600 414.000 1116.750 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2508.065 2553.145 2508.235 2601.255 ;
        RECT 2508.065 2490.925 2508.235 2539.035 ;
      LAYER mcon ;
        RECT 2508.065 2601.085 2508.235 2601.255 ;
        RECT 2508.065 2538.865 2508.235 2539.035 ;
      LAYER met1 ;
        RECT 1987.270 3499.860 1987.590 3499.920 ;
        RECT 1993.710 3499.860 1994.030 3499.920 ;
        RECT 1987.270 3499.720 1994.030 3499.860 ;
        RECT 1987.270 3499.660 1987.590 3499.720 ;
        RECT 1993.710 3499.660 1994.030 3499.720 ;
        RECT 1993.710 3142.860 1994.030 3142.920 ;
        RECT 2507.990 3142.860 2508.310 3142.920 ;
        RECT 1993.710 3142.720 2508.310 3142.860 ;
        RECT 1993.710 3142.660 1994.030 3142.720 ;
        RECT 2507.990 3142.660 2508.310 3142.720 ;
        RECT 2508.910 3042.900 2509.230 3042.960 ;
        RECT 2509.830 3042.900 2510.150 3042.960 ;
        RECT 2508.910 3042.760 2510.150 3042.900 ;
        RECT 2508.910 3042.700 2509.230 3042.760 ;
        RECT 2509.830 3042.700 2510.150 3042.760 ;
        RECT 2508.450 2870.520 2508.770 2870.580 ;
        RECT 2509.830 2870.520 2510.150 2870.580 ;
        RECT 2508.450 2870.380 2510.150 2870.520 ;
        RECT 2508.450 2870.320 2508.770 2870.380 ;
        RECT 2509.830 2870.320 2510.150 2870.380 ;
        RECT 2508.450 2774.300 2508.770 2774.360 ;
        RECT 2508.080 2774.160 2508.770 2774.300 ;
        RECT 2508.080 2774.020 2508.220 2774.160 ;
        RECT 2508.450 2774.100 2508.770 2774.160 ;
        RECT 2507.990 2773.760 2508.310 2774.020 ;
        RECT 2507.990 2684.000 2508.310 2684.260 ;
        RECT 2508.080 2683.520 2508.220 2684.000 ;
        RECT 2508.450 2683.520 2508.770 2683.580 ;
        RECT 2508.080 2683.380 2508.770 2683.520 ;
        RECT 2508.450 2683.320 2508.770 2683.380 ;
        RECT 2508.005 2601.240 2508.295 2601.285 ;
        RECT 2508.450 2601.240 2508.770 2601.300 ;
        RECT 2508.005 2601.100 2508.770 2601.240 ;
        RECT 2508.005 2601.055 2508.295 2601.100 ;
        RECT 2508.450 2601.040 2508.770 2601.100 ;
        RECT 2507.990 2553.300 2508.310 2553.360 ;
        RECT 2507.795 2553.160 2508.310 2553.300 ;
        RECT 2507.990 2553.100 2508.310 2553.160 ;
        RECT 2507.990 2539.020 2508.310 2539.080 ;
        RECT 2507.795 2538.880 2508.310 2539.020 ;
        RECT 2507.990 2538.820 2508.310 2538.880 ;
        RECT 2508.005 2491.080 2508.295 2491.125 ;
        RECT 2508.450 2491.080 2508.770 2491.140 ;
        RECT 2508.005 2490.940 2508.770 2491.080 ;
        RECT 2508.005 2490.895 2508.295 2490.940 ;
        RECT 2508.450 2490.880 2508.770 2490.940 ;
        RECT 2507.990 2401.320 2508.310 2401.380 ;
        RECT 2508.450 2401.320 2508.770 2401.380 ;
        RECT 2507.990 2401.180 2508.770 2401.320 ;
        RECT 2507.990 2401.120 2508.310 2401.180 ;
        RECT 2508.450 2401.120 2508.770 2401.180 ;
        RECT 2507.990 2339.100 2508.310 2339.160 ;
        RECT 2508.450 2339.100 2508.770 2339.160 ;
        RECT 2507.990 2338.960 2508.770 2339.100 ;
        RECT 2507.990 2338.900 2508.310 2338.960 ;
        RECT 2508.450 2338.900 2508.770 2338.960 ;
        RECT 2507.990 2249.680 2508.310 2249.740 ;
        RECT 2508.450 2249.680 2508.770 2249.740 ;
        RECT 2507.990 2249.540 2508.770 2249.680 ;
        RECT 2507.990 2249.480 2508.310 2249.540 ;
        RECT 2508.450 2249.480 2508.770 2249.540 ;
        RECT 2507.990 2242.540 2508.310 2242.600 ;
        RECT 2508.450 2242.540 2508.770 2242.600 ;
        RECT 2507.990 2242.400 2508.770 2242.540 ;
        RECT 2507.990 2242.340 2508.310 2242.400 ;
        RECT 2508.450 2242.340 2508.770 2242.400 ;
        RECT 2507.990 2056.560 2508.310 2056.620 ;
        RECT 2508.910 2056.560 2509.230 2056.620 ;
        RECT 2507.990 2056.420 2509.230 2056.560 ;
        RECT 2507.990 2056.360 2508.310 2056.420 ;
        RECT 2508.910 2056.360 2509.230 2056.420 ;
        RECT 2508.450 1959.660 2508.770 1959.720 ;
        RECT 2508.910 1959.660 2509.230 1959.720 ;
        RECT 2508.450 1959.520 2509.230 1959.660 ;
        RECT 2508.450 1959.460 2508.770 1959.520 ;
        RECT 2508.910 1959.460 2509.230 1959.520 ;
        RECT 2508.450 1883.500 2508.770 1883.560 ;
        RECT 2508.910 1883.500 2509.230 1883.560 ;
        RECT 2508.450 1883.360 2509.230 1883.500 ;
        RECT 2508.450 1883.300 2508.770 1883.360 ;
        RECT 2508.910 1883.300 2509.230 1883.360 ;
        RECT 2508.450 1794.080 2508.770 1794.140 ;
        RECT 2508.910 1794.080 2509.230 1794.140 ;
        RECT 2508.450 1793.940 2509.230 1794.080 ;
        RECT 2508.450 1793.880 2508.770 1793.940 ;
        RECT 2508.910 1793.880 2509.230 1793.940 ;
        RECT 2507.990 1786.940 2508.310 1787.000 ;
        RECT 2508.450 1786.940 2508.770 1787.000 ;
        RECT 2507.990 1786.800 2508.770 1786.940 ;
        RECT 2507.990 1786.740 2508.310 1786.800 ;
        RECT 2508.450 1786.740 2508.770 1786.800 ;
        RECT 2507.990 1697.180 2508.310 1697.240 ;
        RECT 2508.450 1697.180 2508.770 1697.240 ;
        RECT 2507.990 1697.040 2508.770 1697.180 ;
        RECT 2507.990 1696.980 2508.310 1697.040 ;
        RECT 2508.450 1696.980 2508.770 1697.040 ;
      LAYER via ;
        RECT 1987.300 3499.660 1987.560 3499.920 ;
        RECT 1993.740 3499.660 1994.000 3499.920 ;
        RECT 1993.740 3142.660 1994.000 3142.920 ;
        RECT 2508.020 3142.660 2508.280 3142.920 ;
        RECT 2508.940 3042.700 2509.200 3042.960 ;
        RECT 2509.860 3042.700 2510.120 3042.960 ;
        RECT 2508.480 2870.320 2508.740 2870.580 ;
        RECT 2509.860 2870.320 2510.120 2870.580 ;
        RECT 2508.480 2774.100 2508.740 2774.360 ;
        RECT 2508.020 2773.760 2508.280 2774.020 ;
        RECT 2508.020 2684.000 2508.280 2684.260 ;
        RECT 2508.480 2683.320 2508.740 2683.580 ;
        RECT 2508.480 2601.040 2508.740 2601.300 ;
        RECT 2508.020 2553.100 2508.280 2553.360 ;
        RECT 2508.020 2538.820 2508.280 2539.080 ;
        RECT 2508.480 2490.880 2508.740 2491.140 ;
        RECT 2508.020 2401.120 2508.280 2401.380 ;
        RECT 2508.480 2401.120 2508.740 2401.380 ;
        RECT 2508.020 2338.900 2508.280 2339.160 ;
        RECT 2508.480 2338.900 2508.740 2339.160 ;
        RECT 2508.020 2249.480 2508.280 2249.740 ;
        RECT 2508.480 2249.480 2508.740 2249.740 ;
        RECT 2508.020 2242.340 2508.280 2242.600 ;
        RECT 2508.480 2242.340 2508.740 2242.600 ;
        RECT 2508.020 2056.360 2508.280 2056.620 ;
        RECT 2508.940 2056.360 2509.200 2056.620 ;
        RECT 2508.480 1959.460 2508.740 1959.720 ;
        RECT 2508.940 1959.460 2509.200 1959.720 ;
        RECT 2508.480 1883.300 2508.740 1883.560 ;
        RECT 2508.940 1883.300 2509.200 1883.560 ;
        RECT 2508.480 1793.880 2508.740 1794.140 ;
        RECT 2508.940 1793.880 2509.200 1794.140 ;
        RECT 2508.020 1786.740 2508.280 1787.000 ;
        RECT 2508.480 1786.740 2508.740 1787.000 ;
        RECT 2508.020 1696.980 2508.280 1697.240 ;
        RECT 2508.480 1696.980 2508.740 1697.240 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3499.950 1987.500 3517.600 ;
        RECT 1987.300 3499.630 1987.560 3499.950 ;
        RECT 1993.740 3499.630 1994.000 3499.950 ;
        RECT 1993.800 3142.950 1993.940 3499.630 ;
        RECT 1993.740 3142.630 1994.000 3142.950 ;
        RECT 2508.020 3142.630 2508.280 3142.950 ;
        RECT 2508.080 3104.610 2508.220 3142.630 ;
        RECT 2508.080 3104.470 2508.680 3104.610 ;
        RECT 2508.540 3057.010 2508.680 3104.470 ;
        RECT 2508.540 3056.870 2509.140 3057.010 ;
        RECT 2509.000 3042.990 2509.140 3056.870 ;
        RECT 2508.940 3042.670 2509.200 3042.990 ;
        RECT 2509.860 3042.670 2510.120 3042.990 ;
        RECT 2509.920 2870.610 2510.060 3042.670 ;
        RECT 2508.480 2870.290 2508.740 2870.610 ;
        RECT 2509.860 2870.290 2510.120 2870.610 ;
        RECT 2508.540 2774.390 2508.680 2870.290 ;
        RECT 2508.480 2774.070 2508.740 2774.390 ;
        RECT 2508.020 2773.730 2508.280 2774.050 ;
        RECT 2508.080 2684.290 2508.220 2773.730 ;
        RECT 2508.020 2683.970 2508.280 2684.290 ;
        RECT 2508.480 2683.290 2508.740 2683.610 ;
        RECT 2508.540 2622.490 2508.680 2683.290 ;
        RECT 2508.080 2622.350 2508.680 2622.490 ;
        RECT 2508.080 2621.810 2508.220 2622.350 ;
        RECT 2508.080 2621.670 2508.680 2621.810 ;
        RECT 2508.540 2601.330 2508.680 2621.670 ;
        RECT 2508.480 2601.010 2508.740 2601.330 ;
        RECT 2508.020 2553.070 2508.280 2553.390 ;
        RECT 2508.080 2539.110 2508.220 2553.070 ;
        RECT 2508.020 2538.790 2508.280 2539.110 ;
        RECT 2508.480 2490.850 2508.740 2491.170 ;
        RECT 2508.540 2401.410 2508.680 2490.850 ;
        RECT 2508.020 2401.090 2508.280 2401.410 ;
        RECT 2508.480 2401.090 2508.740 2401.410 ;
        RECT 2508.080 2339.190 2508.220 2401.090 ;
        RECT 2508.020 2338.870 2508.280 2339.190 ;
        RECT 2508.480 2338.870 2508.740 2339.190 ;
        RECT 2508.540 2249.770 2508.680 2338.870 ;
        RECT 2508.020 2249.450 2508.280 2249.770 ;
        RECT 2508.480 2249.450 2508.740 2249.770 ;
        RECT 2508.080 2242.630 2508.220 2249.450 ;
        RECT 2508.020 2242.310 2508.280 2242.630 ;
        RECT 2508.480 2242.310 2508.740 2242.630 ;
        RECT 2508.540 2153.405 2508.680 2242.310 ;
        RECT 2508.470 2153.035 2508.750 2153.405 ;
        RECT 2509.390 2152.355 2509.670 2152.725 ;
        RECT 2509.460 2104.840 2509.600 2152.355 ;
        RECT 2509.000 2104.700 2509.600 2104.840 ;
        RECT 2509.000 2056.650 2509.140 2104.700 ;
        RECT 2508.020 2056.330 2508.280 2056.650 ;
        RECT 2508.940 2056.330 2509.200 2056.650 ;
        RECT 2508.080 2026.130 2508.220 2056.330 ;
        RECT 2508.080 2025.990 2509.140 2026.130 ;
        RECT 2509.000 1959.750 2509.140 2025.990 ;
        RECT 2508.480 1959.430 2508.740 1959.750 ;
        RECT 2508.940 1959.430 2509.200 1959.750 ;
        RECT 2508.540 1883.590 2508.680 1959.430 ;
        RECT 2508.480 1883.270 2508.740 1883.590 ;
        RECT 2508.940 1883.270 2509.200 1883.590 ;
        RECT 2509.000 1794.170 2509.140 1883.270 ;
        RECT 2508.480 1793.850 2508.740 1794.170 ;
        RECT 2508.940 1793.850 2509.200 1794.170 ;
        RECT 2508.540 1787.030 2508.680 1793.850 ;
        RECT 2508.020 1786.710 2508.280 1787.030 ;
        RECT 2508.480 1786.710 2508.740 1787.030 ;
        RECT 2508.080 1697.270 2508.220 1786.710 ;
        RECT 2508.020 1696.950 2508.280 1697.270 ;
        RECT 2508.480 1696.950 2508.740 1697.270 ;
        RECT 2508.540 1637.965 2508.680 1696.950 ;
        RECT 2508.470 1637.595 2508.750 1637.965 ;
      LAYER via2 ;
        RECT 2508.470 2153.080 2508.750 2153.360 ;
        RECT 2509.390 2152.400 2509.670 2152.680 ;
        RECT 2508.470 1637.640 2508.750 1637.920 ;
      LAYER met3 ;
        RECT 2508.445 2153.370 2508.775 2153.385 ;
        RECT 2508.230 2153.055 2508.775 2153.370 ;
        RECT 2508.230 2152.690 2508.530 2153.055 ;
        RECT 2509.365 2152.690 2509.695 2152.705 ;
        RECT 2508.230 2152.390 2509.695 2152.690 ;
        RECT 2509.365 2152.375 2509.695 2152.390 ;
        RECT 2508.445 1637.930 2508.775 1637.945 ;
        RECT 2508.230 1637.615 2508.775 1637.930 ;
        RECT 2508.230 1635.360 2508.530 1637.615 ;
        RECT 2506.000 1634.760 2510.000 1635.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3502.580 1662.830 3502.640 ;
        RECT 2602.290 3502.580 2602.610 3502.640 ;
        RECT 1662.510 3502.440 2602.610 3502.580 ;
        RECT 1662.510 3502.380 1662.830 3502.440 ;
        RECT 2602.290 3502.380 2602.610 3502.440 ;
        RECT 2006.130 502.080 2006.450 502.140 ;
        RECT 2602.290 502.080 2602.610 502.140 ;
        RECT 2006.130 501.940 2602.610 502.080 ;
        RECT 2006.130 501.880 2006.450 501.940 ;
        RECT 2602.290 501.880 2602.610 501.940 ;
      LAYER via ;
        RECT 1662.540 3502.380 1662.800 3502.640 ;
        RECT 2602.320 3502.380 2602.580 3502.640 ;
        RECT 2006.160 501.880 2006.420 502.140 ;
        RECT 2602.320 501.880 2602.580 502.140 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3502.670 1662.740 3517.600 ;
        RECT 1662.540 3502.350 1662.800 3502.670 ;
        RECT 2602.320 3502.350 2602.580 3502.670 ;
        RECT 2006.290 510.340 2006.570 514.000 ;
        RECT 2006.220 510.000 2006.570 510.340 ;
        RECT 2006.220 502.170 2006.360 510.000 ;
        RECT 2602.380 502.170 2602.520 3502.350 ;
        RECT 2006.160 501.850 2006.420 502.170 ;
        RECT 2602.320 501.850 2602.580 502.170 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3501.845 1338.440 3517.600 ;
        RECT 1338.230 3501.475 1338.510 3501.845 ;
        RECT 709.090 510.340 709.370 514.000 ;
        RECT 709.020 510.000 709.370 510.340 ;
        RECT 709.020 503.725 709.160 510.000 ;
        RECT 708.950 503.355 709.230 503.725 ;
      LAYER via2 ;
        RECT 1338.230 3501.520 1338.510 3501.800 ;
        RECT 708.950 503.400 709.230 503.680 ;
      LAYER met3 ;
        RECT 344.350 3501.810 344.730 3501.820 ;
        RECT 1338.205 3501.810 1338.535 3501.825 ;
        RECT 344.350 3501.510 1338.535 3501.810 ;
        RECT 344.350 3501.500 344.730 3501.510 ;
        RECT 1338.205 3501.495 1338.535 3501.510 ;
        RECT 344.350 503.690 344.730 503.700 ;
        RECT 708.925 503.690 709.255 503.705 ;
        RECT 344.350 503.390 709.255 503.690 ;
        RECT 344.350 503.380 344.730 503.390 ;
        RECT 708.925 503.375 709.255 503.390 ;
      LAYER via3 ;
        RECT 344.380 3501.500 344.700 3501.820 ;
        RECT 344.380 503.380 344.700 503.700 ;
      LAYER met4 ;
        RECT 344.375 3501.495 344.705 3501.825 ;
        RECT 344.390 503.705 344.690 3501.495 ;
        RECT 344.375 503.375 344.705 503.705 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.970 3006.690 975.250 3010.000 ;
        RECT 976.670 3006.690 976.950 3006.805 ;
        RECT 974.970 3006.550 976.950 3006.690 ;
        RECT 974.970 3006.000 975.250 3006.550 ;
        RECT 976.670 3006.435 976.950 3006.550 ;
      LAYER via2 ;
        RECT 976.670 3006.480 976.950 3006.760 ;
      LAYER met3 ;
        RECT 976.645 3006.770 976.975 3006.785 ;
        RECT 1003.070 3006.770 1003.450 3006.780 ;
        RECT 976.645 3006.470 1003.450 3006.770 ;
        RECT 976.645 3006.455 976.975 3006.470 ;
        RECT 1003.070 3006.460 1003.450 3006.470 ;
        RECT 1003.070 3002.010 1003.450 3002.020 ;
        RECT 2556.030 3002.010 2556.410 3002.020 ;
        RECT 1003.070 3001.710 2556.410 3002.010 ;
        RECT 1003.070 3001.700 1003.450 3001.710 ;
        RECT 2556.030 3001.700 2556.410 3001.710 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 2573.550 436.070 2670.450 436.370 ;
        RECT 2556.030 435.010 2556.410 435.020 ;
        RECT 2573.550 435.010 2573.850 436.070 ;
        RECT 2670.150 435.690 2670.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2670.150 435.390 2718.290 435.690 ;
        RECT 2556.030 434.710 2573.850 435.010 ;
        RECT 2717.990 435.010 2718.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2717.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 2556.030 434.700 2556.410 434.710 ;
      LAYER via3 ;
        RECT 1003.100 3006.460 1003.420 3006.780 ;
        RECT 1003.100 3001.700 1003.420 3002.020 ;
        RECT 2556.060 3001.700 2556.380 3002.020 ;
        RECT 2556.060 434.700 2556.380 435.020 ;
      LAYER met4 ;
        RECT 1003.095 3006.455 1003.425 3006.785 ;
        RECT 1003.110 3002.025 1003.410 3006.455 ;
        RECT 1003.095 3001.695 1003.425 3002.025 ;
        RECT 2556.055 3001.695 2556.385 3002.025 ;
        RECT 2556.070 435.025 2556.370 3001.695 ;
        RECT 2556.055 434.695 2556.385 435.025 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3487.960 1014.230 3488.020 ;
        RECT 2511.670 3487.960 2511.990 3488.020 ;
        RECT 1013.910 3487.820 2511.990 3487.960 ;
        RECT 1013.910 3487.760 1014.230 3487.820 ;
        RECT 2511.670 3487.760 2511.990 3487.820 ;
      LAYER via ;
        RECT 1013.940 3487.760 1014.200 3488.020 ;
        RECT 2511.700 3487.760 2511.960 3488.020 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3488.050 1014.140 3517.600 ;
        RECT 1013.940 3487.730 1014.200 3488.050 ;
        RECT 2511.700 3487.730 2511.960 3488.050 ;
        RECT 2511.760 2677.005 2511.900 3487.730 ;
        RECT 2511.690 2676.635 2511.970 2677.005 ;
      LAYER via2 ;
        RECT 2511.690 2676.680 2511.970 2676.960 ;
      LAYER met3 ;
        RECT 2506.000 2676.970 2510.000 2677.120 ;
        RECT 2511.665 2676.970 2511.995 2676.985 ;
        RECT 2506.000 2676.670 2511.995 2676.970 ;
        RECT 2506.000 2676.520 2510.000 2676.670 ;
        RECT 2511.665 2676.655 2511.995 2676.670 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.600 689.470 3503.660 ;
        RECT 693.290 3503.600 693.610 3503.660 ;
        RECT 689.150 3503.460 693.610 3503.600 ;
        RECT 689.150 3503.400 689.470 3503.460 ;
        RECT 693.290 3503.400 693.610 3503.460 ;
        RECT 693.290 3073.840 693.610 3073.900 ;
        RECT 1911.370 3073.840 1911.690 3073.900 ;
        RECT 693.290 3073.700 1911.690 3073.840 ;
        RECT 693.290 3073.640 693.610 3073.700 ;
        RECT 1911.370 3073.640 1911.690 3073.700 ;
      LAYER via ;
        RECT 689.180 3503.400 689.440 3503.660 ;
        RECT 693.320 3503.400 693.580 3503.660 ;
        RECT 693.320 3073.640 693.580 3073.900 ;
        RECT 1911.400 3073.640 1911.660 3073.900 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.690 689.380 3517.600 ;
        RECT 689.180 3503.370 689.440 3503.690 ;
        RECT 693.320 3503.370 693.580 3503.690 ;
        RECT 693.380 3073.930 693.520 3503.370 ;
        RECT 693.320 3073.610 693.580 3073.930 ;
        RECT 1911.400 3073.610 1911.660 3073.930 ;
        RECT 1911.460 3010.770 1911.600 3073.610 ;
        RECT 1911.460 3010.630 1912.980 3010.770 ;
        RECT 1912.840 3009.410 1912.980 3010.630 ;
        RECT 1914.290 3009.410 1914.570 3010.000 ;
        RECT 1912.840 3009.270 1914.570 3009.410 ;
        RECT 1914.290 3006.000 1914.570 3009.270 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 362.625 3422.865 362.795 3470.635 ;
        RECT 364.005 3380.365 364.175 3422.355 ;
        RECT 364.925 3236.205 365.095 3284.315 ;
        RECT 364.005 3139.645 364.175 3187.755 ;
        RECT 364.925 3043.425 365.095 3090.855 ;
      LAYER mcon ;
        RECT 362.625 3470.465 362.795 3470.635 ;
        RECT 364.005 3422.185 364.175 3422.355 ;
        RECT 364.925 3284.145 365.095 3284.315 ;
        RECT 364.005 3187.585 364.175 3187.755 ;
        RECT 364.925 3090.685 365.095 3090.855 ;
      LAYER met1 ;
        RECT 362.565 3470.620 362.855 3470.665 ;
        RECT 363.470 3470.620 363.790 3470.680 ;
        RECT 362.565 3470.480 363.790 3470.620 ;
        RECT 362.565 3470.435 362.855 3470.480 ;
        RECT 363.470 3470.420 363.790 3470.480 ;
        RECT 362.550 3423.020 362.870 3423.080 ;
        RECT 362.355 3422.880 362.870 3423.020 ;
        RECT 362.550 3422.820 362.870 3422.880 ;
        RECT 362.550 3422.340 362.870 3422.400 ;
        RECT 363.945 3422.340 364.235 3422.385 ;
        RECT 362.550 3422.200 364.235 3422.340 ;
        RECT 362.550 3422.140 362.870 3422.200 ;
        RECT 363.945 3422.155 364.235 3422.200 ;
        RECT 363.930 3380.520 364.250 3380.580 ;
        RECT 363.735 3380.380 364.250 3380.520 ;
        RECT 363.930 3380.320 364.250 3380.380 ;
        RECT 363.930 3346.660 364.250 3346.920 ;
        RECT 364.020 3346.240 364.160 3346.660 ;
        RECT 363.930 3345.980 364.250 3346.240 ;
        RECT 364.390 3298.240 364.710 3298.300 ;
        RECT 365.310 3298.240 365.630 3298.300 ;
        RECT 364.390 3298.100 365.630 3298.240 ;
        RECT 364.390 3298.040 364.710 3298.100 ;
        RECT 365.310 3298.040 365.630 3298.100 ;
        RECT 364.865 3284.300 365.155 3284.345 ;
        RECT 365.310 3284.300 365.630 3284.360 ;
        RECT 364.865 3284.160 365.630 3284.300 ;
        RECT 364.865 3284.115 365.155 3284.160 ;
        RECT 365.310 3284.100 365.630 3284.160 ;
        RECT 364.850 3236.360 365.170 3236.420 ;
        RECT 364.655 3236.220 365.170 3236.360 ;
        RECT 364.850 3236.160 365.170 3236.220 ;
        RECT 364.850 3202.020 365.170 3202.080 ;
        RECT 364.020 3201.880 365.170 3202.020 ;
        RECT 364.020 3201.400 364.160 3201.880 ;
        RECT 364.850 3201.820 365.170 3201.880 ;
        RECT 363.930 3201.140 364.250 3201.400 ;
        RECT 363.930 3187.740 364.250 3187.800 ;
        RECT 363.735 3187.600 364.250 3187.740 ;
        RECT 363.930 3187.540 364.250 3187.600 ;
        RECT 363.945 3139.800 364.235 3139.845 ;
        RECT 365.310 3139.800 365.630 3139.860 ;
        RECT 363.945 3139.660 365.630 3139.800 ;
        RECT 363.945 3139.615 364.235 3139.660 ;
        RECT 365.310 3139.600 365.630 3139.660 ;
        RECT 364.850 3091.520 365.170 3091.580 ;
        RECT 365.310 3091.520 365.630 3091.580 ;
        RECT 364.850 3091.380 365.630 3091.520 ;
        RECT 364.850 3091.320 365.170 3091.380 ;
        RECT 365.310 3091.320 365.630 3091.380 ;
        RECT 364.850 3090.840 365.170 3090.900 ;
        RECT 364.655 3090.700 365.170 3090.840 ;
        RECT 364.850 3090.640 365.170 3090.700 ;
        RECT 364.865 3043.580 365.155 3043.625 ;
        RECT 365.310 3043.580 365.630 3043.640 ;
        RECT 364.865 3043.440 365.630 3043.580 ;
        RECT 364.865 3043.395 365.155 3043.440 ;
        RECT 365.310 3043.380 365.630 3043.440 ;
        RECT 363.930 2932.400 364.250 2932.460 ;
        RECT 365.310 2932.400 365.630 2932.460 ;
        RECT 363.930 2932.260 365.630 2932.400 ;
        RECT 363.930 2932.200 364.250 2932.260 ;
        RECT 365.310 2932.200 365.630 2932.260 ;
        RECT 363.930 2884.460 364.250 2884.520 ;
        RECT 365.310 2884.460 365.630 2884.520 ;
        RECT 363.930 2884.320 365.630 2884.460 ;
        RECT 363.930 2884.260 364.250 2884.320 ;
        RECT 365.310 2884.260 365.630 2884.320 ;
        RECT 363.930 2739.280 364.250 2739.340 ;
        RECT 365.310 2739.280 365.630 2739.340 ;
        RECT 363.930 2739.140 365.630 2739.280 ;
        RECT 363.930 2739.080 364.250 2739.140 ;
        RECT 365.310 2739.080 365.630 2739.140 ;
        RECT 363.930 2691.340 364.250 2691.400 ;
        RECT 365.310 2691.340 365.630 2691.400 ;
        RECT 363.930 2691.200 365.630 2691.340 ;
        RECT 363.930 2691.140 364.250 2691.200 ;
        RECT 365.310 2691.140 365.630 2691.200 ;
        RECT 363.930 2449.260 364.250 2449.320 ;
        RECT 365.310 2449.260 365.630 2449.320 ;
        RECT 363.930 2449.120 365.630 2449.260 ;
        RECT 363.930 2449.060 364.250 2449.120 ;
        RECT 365.310 2449.060 365.630 2449.120 ;
        RECT 363.930 2401.320 364.250 2401.380 ;
        RECT 365.310 2401.320 365.630 2401.380 ;
        RECT 363.930 2401.180 365.630 2401.320 ;
        RECT 363.930 2401.120 364.250 2401.180 ;
        RECT 365.310 2401.120 365.630 2401.180 ;
        RECT 363.930 2256.140 364.250 2256.200 ;
        RECT 365.310 2256.140 365.630 2256.200 ;
        RECT 363.930 2256.000 365.630 2256.140 ;
        RECT 363.930 2255.940 364.250 2256.000 ;
        RECT 365.310 2255.940 365.630 2256.000 ;
        RECT 363.930 2208.540 364.250 2208.600 ;
        RECT 365.310 2208.540 365.630 2208.600 ;
        RECT 363.930 2208.400 365.630 2208.540 ;
        RECT 363.930 2208.340 364.250 2208.400 ;
        RECT 365.310 2208.340 365.630 2208.400 ;
        RECT 363.930 2159.580 364.250 2159.640 ;
        RECT 365.310 2159.580 365.630 2159.640 ;
        RECT 363.930 2159.440 365.630 2159.580 ;
        RECT 363.930 2159.380 364.250 2159.440 ;
        RECT 365.310 2159.380 365.630 2159.440 ;
        RECT 363.930 2111.640 364.250 2111.700 ;
        RECT 365.310 2111.640 365.630 2111.700 ;
        RECT 363.930 2111.500 365.630 2111.640 ;
        RECT 363.930 2111.440 364.250 2111.500 ;
        RECT 365.310 2111.440 365.630 2111.500 ;
        RECT 363.930 2063.020 364.250 2063.080 ;
        RECT 365.310 2063.020 365.630 2063.080 ;
        RECT 363.930 2062.880 365.630 2063.020 ;
        RECT 363.930 2062.820 364.250 2062.880 ;
        RECT 365.310 2062.820 365.630 2062.880 ;
        RECT 363.930 2015.080 364.250 2015.140 ;
        RECT 365.310 2015.080 365.630 2015.140 ;
        RECT 363.930 2014.940 365.630 2015.080 ;
        RECT 363.930 2014.880 364.250 2014.940 ;
        RECT 365.310 2014.880 365.630 2014.940 ;
        RECT 363.930 1966.460 364.250 1966.520 ;
        RECT 365.310 1966.460 365.630 1966.520 ;
        RECT 363.930 1966.320 365.630 1966.460 ;
        RECT 363.930 1966.260 364.250 1966.320 ;
        RECT 365.310 1966.260 365.630 1966.320 ;
        RECT 363.930 1918.860 364.250 1918.920 ;
        RECT 365.310 1918.860 365.630 1918.920 ;
        RECT 363.930 1918.720 365.630 1918.860 ;
        RECT 363.930 1918.660 364.250 1918.720 ;
        RECT 365.310 1918.660 365.630 1918.720 ;
        RECT 363.930 1869.900 364.250 1869.960 ;
        RECT 365.310 1869.900 365.630 1869.960 ;
        RECT 363.930 1869.760 365.630 1869.900 ;
        RECT 363.930 1869.700 364.250 1869.760 ;
        RECT 365.310 1869.700 365.630 1869.760 ;
        RECT 363.930 1821.960 364.250 1822.020 ;
        RECT 365.310 1821.960 365.630 1822.020 ;
        RECT 363.930 1821.820 365.630 1821.960 ;
        RECT 363.930 1821.760 364.250 1821.820 ;
        RECT 365.310 1821.760 365.630 1821.820 ;
        RECT 363.930 1579.880 364.250 1579.940 ;
        RECT 365.310 1579.880 365.630 1579.940 ;
        RECT 363.930 1579.740 365.630 1579.880 ;
        RECT 363.930 1579.680 364.250 1579.740 ;
        RECT 365.310 1579.680 365.630 1579.740 ;
        RECT 363.930 1531.940 364.250 1532.000 ;
        RECT 365.310 1531.940 365.630 1532.000 ;
        RECT 363.930 1531.800 365.630 1531.940 ;
        RECT 363.930 1531.740 364.250 1531.800 ;
        RECT 365.310 1531.740 365.630 1531.800 ;
        RECT 363.930 1483.320 364.250 1483.380 ;
        RECT 365.310 1483.320 365.630 1483.380 ;
        RECT 363.930 1483.180 365.630 1483.320 ;
        RECT 363.930 1483.120 364.250 1483.180 ;
        RECT 365.310 1483.120 365.630 1483.180 ;
        RECT 363.930 1435.380 364.250 1435.440 ;
        RECT 365.310 1435.380 365.630 1435.440 ;
        RECT 363.930 1435.240 365.630 1435.380 ;
        RECT 363.930 1435.180 364.250 1435.240 ;
        RECT 365.310 1435.180 365.630 1435.240 ;
        RECT 363.470 1386.760 363.790 1386.820 ;
        RECT 365.310 1386.760 365.630 1386.820 ;
        RECT 363.470 1386.620 365.630 1386.760 ;
        RECT 363.470 1386.560 363.790 1386.620 ;
        RECT 365.310 1386.560 365.630 1386.620 ;
        RECT 363.470 1338.820 363.790 1338.880 ;
        RECT 365.310 1338.820 365.630 1338.880 ;
        RECT 363.470 1338.680 365.630 1338.820 ;
        RECT 363.470 1338.620 363.790 1338.680 ;
        RECT 365.310 1338.620 365.630 1338.680 ;
        RECT 363.470 1293.940 363.790 1294.000 ;
        RECT 365.310 1293.940 365.630 1294.000 ;
        RECT 363.470 1293.800 365.630 1293.940 ;
        RECT 363.470 1293.740 363.790 1293.800 ;
        RECT 365.310 1293.740 365.630 1293.800 ;
        RECT 363.470 1245.660 363.790 1245.720 ;
        RECT 365.310 1245.660 365.630 1245.720 ;
        RECT 363.470 1245.520 365.630 1245.660 ;
        RECT 363.470 1245.460 363.790 1245.520 ;
        RECT 365.310 1245.460 365.630 1245.520 ;
        RECT 363.470 1197.380 363.790 1197.440 ;
        RECT 365.310 1197.380 365.630 1197.440 ;
        RECT 363.470 1197.240 365.630 1197.380 ;
        RECT 363.470 1197.180 363.790 1197.240 ;
        RECT 365.310 1197.180 365.630 1197.240 ;
        RECT 363.470 1148.760 363.790 1148.820 ;
        RECT 365.310 1148.760 365.630 1148.820 ;
        RECT 363.470 1148.620 365.630 1148.760 ;
        RECT 363.470 1148.560 363.790 1148.620 ;
        RECT 365.310 1148.560 365.630 1148.620 ;
        RECT 363.470 1084.840 363.790 1084.900 ;
        RECT 365.310 1084.840 365.630 1084.900 ;
        RECT 363.470 1084.700 365.630 1084.840 ;
        RECT 363.470 1084.640 363.790 1084.700 ;
        RECT 365.310 1084.640 365.630 1084.700 ;
        RECT 363.470 1052.200 363.790 1052.260 ;
        RECT 365.310 1052.200 365.630 1052.260 ;
        RECT 363.470 1052.060 365.630 1052.200 ;
        RECT 363.470 1052.000 363.790 1052.060 ;
        RECT 365.310 1052.000 365.630 1052.060 ;
        RECT 361.630 1003.920 361.950 1003.980 ;
        RECT 365.310 1003.920 365.630 1003.980 ;
        RECT 361.630 1003.780 365.630 1003.920 ;
        RECT 361.630 1003.720 361.950 1003.780 ;
        RECT 365.310 1003.720 365.630 1003.780 ;
        RECT 361.630 903.960 361.950 904.020 ;
        RECT 365.310 903.960 365.630 904.020 ;
        RECT 361.630 903.820 365.630 903.960 ;
        RECT 361.630 903.760 361.950 903.820 ;
        RECT 365.310 903.760 365.630 903.820 ;
        RECT 361.630 856.020 361.950 856.080 ;
        RECT 365.310 856.020 365.630 856.080 ;
        RECT 361.630 855.880 365.630 856.020 ;
        RECT 361.630 855.820 361.950 855.880 ;
        RECT 365.310 855.820 365.630 855.880 ;
        RECT 362.090 807.060 362.410 807.120 ;
        RECT 365.310 807.060 365.630 807.120 ;
        RECT 362.090 806.920 365.630 807.060 ;
        RECT 362.090 806.860 362.410 806.920 ;
        RECT 365.310 806.860 365.630 806.920 ;
        RECT 362.090 759.120 362.410 759.180 ;
        RECT 365.310 759.120 365.630 759.180 ;
        RECT 362.090 758.980 365.630 759.120 ;
        RECT 362.090 758.920 362.410 758.980 ;
        RECT 365.310 758.920 365.630 758.980 ;
        RECT 362.090 710.500 362.410 710.560 ;
        RECT 365.310 710.500 365.630 710.560 ;
        RECT 362.090 710.360 365.630 710.500 ;
        RECT 362.090 710.300 362.410 710.360 ;
        RECT 365.310 710.300 365.630 710.360 ;
        RECT 362.090 662.560 362.410 662.620 ;
        RECT 365.310 662.560 365.630 662.620 ;
        RECT 362.090 662.420 365.630 662.560 ;
        RECT 362.090 662.360 362.410 662.420 ;
        RECT 365.310 662.360 365.630 662.420 ;
        RECT 361.630 613.940 361.950 614.000 ;
        RECT 365.310 613.940 365.630 614.000 ;
        RECT 361.630 613.800 365.630 613.940 ;
        RECT 361.630 613.740 361.950 613.800 ;
        RECT 365.310 613.740 365.630 613.800 ;
        RECT 361.630 566.000 361.950 566.060 ;
        RECT 365.310 566.000 365.630 566.060 ;
        RECT 361.630 565.860 365.630 566.000 ;
        RECT 361.630 565.800 361.950 565.860 ;
        RECT 365.310 565.800 365.630 565.860 ;
        RECT 365.310 552.060 365.630 552.120 ;
        RECT 393.370 552.060 393.690 552.120 ;
        RECT 365.310 551.920 393.690 552.060 ;
        RECT 365.310 551.860 365.630 551.920 ;
        RECT 393.370 551.860 393.690 551.920 ;
      LAYER via ;
        RECT 363.500 3470.420 363.760 3470.680 ;
        RECT 362.580 3422.820 362.840 3423.080 ;
        RECT 362.580 3422.140 362.840 3422.400 ;
        RECT 363.960 3380.320 364.220 3380.580 ;
        RECT 363.960 3346.660 364.220 3346.920 ;
        RECT 363.960 3345.980 364.220 3346.240 ;
        RECT 364.420 3298.040 364.680 3298.300 ;
        RECT 365.340 3298.040 365.600 3298.300 ;
        RECT 365.340 3284.100 365.600 3284.360 ;
        RECT 364.880 3236.160 365.140 3236.420 ;
        RECT 364.880 3201.820 365.140 3202.080 ;
        RECT 363.960 3201.140 364.220 3201.400 ;
        RECT 363.960 3187.540 364.220 3187.800 ;
        RECT 365.340 3139.600 365.600 3139.860 ;
        RECT 364.880 3091.320 365.140 3091.580 ;
        RECT 365.340 3091.320 365.600 3091.580 ;
        RECT 364.880 3090.640 365.140 3090.900 ;
        RECT 365.340 3043.380 365.600 3043.640 ;
        RECT 363.960 2932.200 364.220 2932.460 ;
        RECT 365.340 2932.200 365.600 2932.460 ;
        RECT 363.960 2884.260 364.220 2884.520 ;
        RECT 365.340 2884.260 365.600 2884.520 ;
        RECT 363.960 2739.080 364.220 2739.340 ;
        RECT 365.340 2739.080 365.600 2739.340 ;
        RECT 363.960 2691.140 364.220 2691.400 ;
        RECT 365.340 2691.140 365.600 2691.400 ;
        RECT 363.960 2449.060 364.220 2449.320 ;
        RECT 365.340 2449.060 365.600 2449.320 ;
        RECT 363.960 2401.120 364.220 2401.380 ;
        RECT 365.340 2401.120 365.600 2401.380 ;
        RECT 363.960 2255.940 364.220 2256.200 ;
        RECT 365.340 2255.940 365.600 2256.200 ;
        RECT 363.960 2208.340 364.220 2208.600 ;
        RECT 365.340 2208.340 365.600 2208.600 ;
        RECT 363.960 2159.380 364.220 2159.640 ;
        RECT 365.340 2159.380 365.600 2159.640 ;
        RECT 363.960 2111.440 364.220 2111.700 ;
        RECT 365.340 2111.440 365.600 2111.700 ;
        RECT 363.960 2062.820 364.220 2063.080 ;
        RECT 365.340 2062.820 365.600 2063.080 ;
        RECT 363.960 2014.880 364.220 2015.140 ;
        RECT 365.340 2014.880 365.600 2015.140 ;
        RECT 363.960 1966.260 364.220 1966.520 ;
        RECT 365.340 1966.260 365.600 1966.520 ;
        RECT 363.960 1918.660 364.220 1918.920 ;
        RECT 365.340 1918.660 365.600 1918.920 ;
        RECT 363.960 1869.700 364.220 1869.960 ;
        RECT 365.340 1869.700 365.600 1869.960 ;
        RECT 363.960 1821.760 364.220 1822.020 ;
        RECT 365.340 1821.760 365.600 1822.020 ;
        RECT 363.960 1579.680 364.220 1579.940 ;
        RECT 365.340 1579.680 365.600 1579.940 ;
        RECT 363.960 1531.740 364.220 1532.000 ;
        RECT 365.340 1531.740 365.600 1532.000 ;
        RECT 363.960 1483.120 364.220 1483.380 ;
        RECT 365.340 1483.120 365.600 1483.380 ;
        RECT 363.960 1435.180 364.220 1435.440 ;
        RECT 365.340 1435.180 365.600 1435.440 ;
        RECT 363.500 1386.560 363.760 1386.820 ;
        RECT 365.340 1386.560 365.600 1386.820 ;
        RECT 363.500 1338.620 363.760 1338.880 ;
        RECT 365.340 1338.620 365.600 1338.880 ;
        RECT 363.500 1293.740 363.760 1294.000 ;
        RECT 365.340 1293.740 365.600 1294.000 ;
        RECT 363.500 1245.460 363.760 1245.720 ;
        RECT 365.340 1245.460 365.600 1245.720 ;
        RECT 363.500 1197.180 363.760 1197.440 ;
        RECT 365.340 1197.180 365.600 1197.440 ;
        RECT 363.500 1148.560 363.760 1148.820 ;
        RECT 365.340 1148.560 365.600 1148.820 ;
        RECT 363.500 1084.640 363.760 1084.900 ;
        RECT 365.340 1084.640 365.600 1084.900 ;
        RECT 363.500 1052.000 363.760 1052.260 ;
        RECT 365.340 1052.000 365.600 1052.260 ;
        RECT 361.660 1003.720 361.920 1003.980 ;
        RECT 365.340 1003.720 365.600 1003.980 ;
        RECT 361.660 903.760 361.920 904.020 ;
        RECT 365.340 903.760 365.600 904.020 ;
        RECT 361.660 855.820 361.920 856.080 ;
        RECT 365.340 855.820 365.600 856.080 ;
        RECT 362.120 806.860 362.380 807.120 ;
        RECT 365.340 806.860 365.600 807.120 ;
        RECT 362.120 758.920 362.380 759.180 ;
        RECT 365.340 758.920 365.600 759.180 ;
        RECT 362.120 710.300 362.380 710.560 ;
        RECT 365.340 710.300 365.600 710.560 ;
        RECT 362.120 662.360 362.380 662.620 ;
        RECT 365.340 662.360 365.600 662.620 ;
        RECT 361.660 613.740 361.920 614.000 ;
        RECT 365.340 613.740 365.600 614.000 ;
        RECT 361.660 565.800 361.920 566.060 ;
        RECT 365.340 565.800 365.600 566.060 ;
        RECT 365.340 551.860 365.600 552.120 ;
        RECT 393.400 551.860 393.660 552.120 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3517.370 365.080 3517.600 ;
        RECT 364.020 3517.230 365.080 3517.370 ;
        RECT 364.020 3491.530 364.160 3517.230 ;
        RECT 363.560 3491.390 364.160 3491.530 ;
        RECT 363.560 3470.710 363.700 3491.390 ;
        RECT 363.500 3470.390 363.760 3470.710 ;
        RECT 362.580 3422.790 362.840 3423.110 ;
        RECT 362.640 3422.430 362.780 3422.790 ;
        RECT 362.580 3422.110 362.840 3422.430 ;
        RECT 363.960 3380.290 364.220 3380.610 ;
        RECT 364.020 3346.950 364.160 3380.290 ;
        RECT 363.960 3346.630 364.220 3346.950 ;
        RECT 363.960 3345.950 364.220 3346.270 ;
        RECT 364.020 3298.410 364.160 3345.950 ;
        RECT 364.020 3298.330 364.620 3298.410 ;
        RECT 364.020 3298.270 364.680 3298.330 ;
        RECT 364.420 3298.010 364.680 3298.270 ;
        RECT 365.340 3298.010 365.600 3298.330 ;
        RECT 365.400 3284.390 365.540 3298.010 ;
        RECT 365.340 3284.070 365.600 3284.390 ;
        RECT 364.880 3236.130 365.140 3236.450 ;
        RECT 364.940 3202.110 365.080 3236.130 ;
        RECT 364.880 3201.790 365.140 3202.110 ;
        RECT 363.960 3201.110 364.220 3201.430 ;
        RECT 364.020 3187.830 364.160 3201.110 ;
        RECT 363.960 3187.510 364.220 3187.830 ;
        RECT 365.340 3139.570 365.600 3139.890 ;
        RECT 365.400 3091.610 365.540 3139.570 ;
        RECT 364.880 3091.290 365.140 3091.610 ;
        RECT 365.340 3091.290 365.600 3091.610 ;
        RECT 364.940 3090.930 365.080 3091.290 ;
        RECT 364.880 3090.610 365.140 3090.930 ;
        RECT 365.340 3043.350 365.600 3043.670 ;
        RECT 365.400 2932.490 365.540 3043.350 ;
        RECT 363.960 2932.170 364.220 2932.490 ;
        RECT 365.340 2932.170 365.600 2932.490 ;
        RECT 364.020 2884.550 364.160 2932.170 ;
        RECT 363.960 2884.230 364.220 2884.550 ;
        RECT 365.340 2884.230 365.600 2884.550 ;
        RECT 365.400 2739.370 365.540 2884.230 ;
        RECT 363.960 2739.050 364.220 2739.370 ;
        RECT 365.340 2739.050 365.600 2739.370 ;
        RECT 364.020 2691.430 364.160 2739.050 ;
        RECT 363.960 2691.110 364.220 2691.430 ;
        RECT 365.340 2691.110 365.600 2691.430 ;
        RECT 365.400 2449.350 365.540 2691.110 ;
        RECT 363.960 2449.030 364.220 2449.350 ;
        RECT 365.340 2449.030 365.600 2449.350 ;
        RECT 364.020 2401.410 364.160 2449.030 ;
        RECT 363.960 2401.090 364.220 2401.410 ;
        RECT 365.340 2401.090 365.600 2401.410 ;
        RECT 365.400 2256.230 365.540 2401.090 ;
        RECT 363.960 2255.910 364.220 2256.230 ;
        RECT 365.340 2255.910 365.600 2256.230 ;
        RECT 364.020 2208.630 364.160 2255.910 ;
        RECT 363.960 2208.310 364.220 2208.630 ;
        RECT 365.340 2208.310 365.600 2208.630 ;
        RECT 365.400 2159.670 365.540 2208.310 ;
        RECT 363.960 2159.350 364.220 2159.670 ;
        RECT 365.340 2159.350 365.600 2159.670 ;
        RECT 364.020 2111.730 364.160 2159.350 ;
        RECT 363.960 2111.410 364.220 2111.730 ;
        RECT 365.340 2111.410 365.600 2111.730 ;
        RECT 365.400 2063.110 365.540 2111.410 ;
        RECT 363.960 2062.790 364.220 2063.110 ;
        RECT 365.340 2062.790 365.600 2063.110 ;
        RECT 364.020 2015.170 364.160 2062.790 ;
        RECT 363.960 2014.850 364.220 2015.170 ;
        RECT 365.340 2014.850 365.600 2015.170 ;
        RECT 365.400 1966.550 365.540 2014.850 ;
        RECT 363.960 1966.230 364.220 1966.550 ;
        RECT 365.340 1966.230 365.600 1966.550 ;
        RECT 364.020 1918.950 364.160 1966.230 ;
        RECT 363.960 1918.630 364.220 1918.950 ;
        RECT 365.340 1918.630 365.600 1918.950 ;
        RECT 365.400 1869.990 365.540 1918.630 ;
        RECT 363.960 1869.670 364.220 1869.990 ;
        RECT 365.340 1869.670 365.600 1869.990 ;
        RECT 364.020 1822.050 364.160 1869.670 ;
        RECT 363.960 1821.730 364.220 1822.050 ;
        RECT 365.340 1821.730 365.600 1822.050 ;
        RECT 365.400 1579.970 365.540 1821.730 ;
        RECT 363.960 1579.650 364.220 1579.970 ;
        RECT 365.340 1579.650 365.600 1579.970 ;
        RECT 364.020 1532.030 364.160 1579.650 ;
        RECT 363.960 1531.710 364.220 1532.030 ;
        RECT 365.340 1531.710 365.600 1532.030 ;
        RECT 365.400 1483.410 365.540 1531.710 ;
        RECT 363.960 1483.090 364.220 1483.410 ;
        RECT 365.340 1483.090 365.600 1483.410 ;
        RECT 364.020 1435.470 364.160 1483.090 ;
        RECT 363.960 1435.150 364.220 1435.470 ;
        RECT 365.340 1435.150 365.600 1435.470 ;
        RECT 365.400 1386.850 365.540 1435.150 ;
        RECT 363.500 1386.530 363.760 1386.850 ;
        RECT 365.340 1386.530 365.600 1386.850 ;
        RECT 363.560 1338.910 363.700 1386.530 ;
        RECT 363.500 1338.590 363.760 1338.910 ;
        RECT 365.340 1338.590 365.600 1338.910 ;
        RECT 365.400 1294.030 365.540 1338.590 ;
        RECT 363.500 1293.710 363.760 1294.030 ;
        RECT 365.340 1293.710 365.600 1294.030 ;
        RECT 363.560 1245.750 363.700 1293.710 ;
        RECT 363.500 1245.430 363.760 1245.750 ;
        RECT 365.340 1245.430 365.600 1245.750 ;
        RECT 365.400 1197.470 365.540 1245.430 ;
        RECT 363.500 1197.150 363.760 1197.470 ;
        RECT 365.340 1197.150 365.600 1197.470 ;
        RECT 363.560 1148.850 363.700 1197.150 ;
        RECT 363.500 1148.530 363.760 1148.850 ;
        RECT 365.340 1148.530 365.600 1148.850 ;
        RECT 365.400 1084.930 365.540 1148.530 ;
        RECT 363.500 1084.610 363.760 1084.930 ;
        RECT 365.340 1084.610 365.600 1084.930 ;
        RECT 363.560 1052.290 363.700 1084.610 ;
        RECT 363.500 1051.970 363.760 1052.290 ;
        RECT 365.340 1051.970 365.600 1052.290 ;
        RECT 365.400 1004.010 365.540 1051.970 ;
        RECT 361.660 1003.690 361.920 1004.010 ;
        RECT 365.340 1003.690 365.600 1004.010 ;
        RECT 361.720 952.525 361.860 1003.690 ;
        RECT 361.650 952.155 361.930 952.525 ;
        RECT 365.330 952.155 365.610 952.525 ;
        RECT 365.400 904.050 365.540 952.155 ;
        RECT 361.660 903.730 361.920 904.050 ;
        RECT 365.340 903.730 365.600 904.050 ;
        RECT 361.720 856.110 361.860 903.730 ;
        RECT 361.660 855.790 361.920 856.110 ;
        RECT 365.340 855.790 365.600 856.110 ;
        RECT 365.400 807.150 365.540 855.790 ;
        RECT 362.120 806.830 362.380 807.150 ;
        RECT 365.340 806.830 365.600 807.150 ;
        RECT 362.180 759.210 362.320 806.830 ;
        RECT 362.120 758.890 362.380 759.210 ;
        RECT 365.340 758.890 365.600 759.210 ;
        RECT 365.400 710.590 365.540 758.890 ;
        RECT 362.120 710.270 362.380 710.590 ;
        RECT 365.340 710.270 365.600 710.590 ;
        RECT 362.180 662.650 362.320 710.270 ;
        RECT 362.120 662.330 362.380 662.650 ;
        RECT 365.340 662.330 365.600 662.650 ;
        RECT 365.400 614.030 365.540 662.330 ;
        RECT 361.660 613.710 361.920 614.030 ;
        RECT 365.340 613.710 365.600 614.030 ;
        RECT 361.720 566.090 361.860 613.710 ;
        RECT 361.660 565.770 361.920 566.090 ;
        RECT 365.340 565.770 365.600 566.090 ;
        RECT 365.400 552.150 365.540 565.770 ;
        RECT 365.340 551.830 365.600 552.150 ;
        RECT 393.400 551.830 393.660 552.150 ;
        RECT 393.460 549.965 393.600 551.830 ;
        RECT 393.390 549.595 393.670 549.965 ;
      LAYER via2 ;
        RECT 361.650 952.200 361.930 952.480 ;
        RECT 365.330 952.200 365.610 952.480 ;
        RECT 393.390 549.640 393.670 549.920 ;
      LAYER met3 ;
        RECT 361.625 952.490 361.955 952.505 ;
        RECT 365.305 952.490 365.635 952.505 ;
        RECT 361.625 952.190 365.635 952.490 ;
        RECT 361.625 952.175 361.955 952.190 ;
        RECT 365.305 952.175 365.635 952.190 ;
        RECT 393.365 549.930 393.695 549.945 ;
        RECT 410.000 549.930 414.000 550.080 ;
        RECT 393.365 549.630 414.000 549.930 ;
        RECT 393.365 549.615 393.695 549.630 ;
        RECT 410.000 549.480 414.000 549.630 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.220 40.870 3501.280 ;
        RECT 72.290 3501.220 72.610 3501.280 ;
        RECT 40.550 3501.080 72.610 3501.220 ;
        RECT 40.550 3501.020 40.870 3501.080 ;
        RECT 72.290 3501.020 72.610 3501.080 ;
        RECT 72.290 793.460 72.610 793.520 ;
        RECT 393.370 793.460 393.690 793.520 ;
        RECT 72.290 793.320 393.690 793.460 ;
        RECT 72.290 793.260 72.610 793.320 ;
        RECT 393.370 793.260 393.690 793.320 ;
      LAYER via ;
        RECT 40.580 3501.020 40.840 3501.280 ;
        RECT 72.320 3501.020 72.580 3501.280 ;
        RECT 72.320 793.260 72.580 793.520 ;
        RECT 393.400 793.260 393.660 793.520 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.310 40.780 3517.600 ;
        RECT 40.580 3500.990 40.840 3501.310 ;
        RECT 72.320 3500.990 72.580 3501.310 ;
        RECT 72.380 793.550 72.520 3500.990 ;
        RECT 72.320 793.230 72.580 793.550 ;
        RECT 393.400 793.230 393.660 793.550 ;
        RECT 393.460 787.965 393.600 793.230 ;
        RECT 393.390 787.595 393.670 787.965 ;
      LAYER via2 ;
        RECT 393.390 787.640 393.670 787.920 ;
      LAYER met3 ;
        RECT 393.365 787.930 393.695 787.945 ;
        RECT 410.000 787.930 414.000 788.080 ;
        RECT 393.365 787.630 414.000 787.930 ;
        RECT 393.365 787.615 393.695 787.630 ;
        RECT 410.000 787.480 414.000 787.630 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 86.090 3263.900 86.410 3263.960 ;
        RECT 15.250 3263.760 86.410 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 86.090 3263.700 86.410 3263.760 ;
        RECT 86.090 1648.900 86.410 1648.960 ;
        RECT 393.370 1648.900 393.690 1648.960 ;
        RECT 86.090 1648.760 393.690 1648.900 ;
        RECT 86.090 1648.700 86.410 1648.760 ;
        RECT 393.370 1648.700 393.690 1648.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 86.120 3263.700 86.380 3263.960 ;
        RECT 86.120 1648.700 86.380 1648.960 ;
        RECT 393.400 1648.700 393.660 1648.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 86.120 3263.670 86.380 3263.990 ;
        RECT 86.180 1648.990 86.320 3263.670 ;
        RECT 86.120 1648.670 86.380 1648.990 ;
        RECT 393.400 1648.670 393.660 1648.990 ;
        RECT 393.460 1646.125 393.600 1648.670 ;
        RECT 393.390 1645.755 393.670 1646.125 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 393.390 1645.800 393.670 1646.080 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 393.365 1646.090 393.695 1646.105 ;
        RECT 410.000 1646.090 414.000 1646.240 ;
        RECT 393.365 1645.790 414.000 1646.090 ;
        RECT 393.365 1645.775 393.695 1645.790 ;
        RECT 410.000 1645.640 414.000 1645.790 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 882.885 482.545 884.895 482.715 ;
        RECT 1781.725 482.545 1783.735 482.715 ;
      LAYER mcon ;
        RECT 884.725 482.545 884.895 482.715 ;
        RECT 1783.565 482.545 1783.735 482.715 ;
      LAYER met1 ;
        RECT 14.330 2974.220 14.650 2974.280 ;
        RECT 161.990 2974.220 162.310 2974.280 ;
        RECT 14.330 2974.080 162.310 2974.220 ;
        RECT 14.330 2974.020 14.650 2974.080 ;
        RECT 161.990 2974.020 162.310 2974.080 ;
        RECT 161.990 482.700 162.310 482.760 ;
        RECT 882.825 482.700 883.115 482.745 ;
        RECT 161.990 482.560 883.115 482.700 ;
        RECT 161.990 482.500 162.310 482.560 ;
        RECT 882.825 482.515 883.115 482.560 ;
        RECT 884.665 482.700 884.955 482.745 ;
        RECT 1781.665 482.700 1781.955 482.745 ;
        RECT 884.665 482.560 1781.955 482.700 ;
        RECT 884.665 482.515 884.955 482.560 ;
        RECT 1781.665 482.515 1781.955 482.560 ;
        RECT 1783.505 482.700 1783.795 482.745 ;
        RECT 2067.770 482.700 2068.090 482.760 ;
        RECT 1783.505 482.560 2068.090 482.700 ;
        RECT 1783.505 482.515 1783.795 482.560 ;
        RECT 2067.770 482.500 2068.090 482.560 ;
      LAYER via ;
        RECT 14.360 2974.020 14.620 2974.280 ;
        RECT 162.020 2974.020 162.280 2974.280 ;
        RECT 162.020 482.500 162.280 482.760 ;
        RECT 2067.800 482.500 2068.060 482.760 ;
      LAYER met2 ;
        RECT 14.350 2979.915 14.630 2980.285 ;
        RECT 14.420 2974.310 14.560 2979.915 ;
        RECT 14.360 2973.990 14.620 2974.310 ;
        RECT 162.020 2973.990 162.280 2974.310 ;
        RECT 162.080 482.790 162.220 2973.990 ;
        RECT 2067.930 510.340 2068.210 514.000 ;
        RECT 2067.860 510.000 2068.210 510.340 ;
        RECT 2067.860 482.790 2068.000 510.000 ;
        RECT 162.020 482.470 162.280 482.790 ;
        RECT 2067.800 482.470 2068.060 482.790 ;
      LAYER via2 ;
        RECT 14.350 2979.960 14.630 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 14.325 2980.250 14.655 2980.265 ;
        RECT -4.800 2979.950 14.655 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 14.325 2979.935 14.655 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2691.340 17.410 2691.400 ;
        RECT 217.190 2691.340 217.510 2691.400 ;
        RECT 17.090 2691.200 217.510 2691.340 ;
        RECT 17.090 2691.140 17.410 2691.200 ;
        RECT 217.190 2691.140 217.510 2691.200 ;
        RECT 217.190 489.500 217.510 489.560 ;
        RECT 1733.810 489.500 1734.130 489.560 ;
        RECT 217.190 489.360 1734.130 489.500 ;
        RECT 217.190 489.300 217.510 489.360 ;
        RECT 1733.810 489.300 1734.130 489.360 ;
      LAYER via ;
        RECT 17.120 2691.140 17.380 2691.400 ;
        RECT 217.220 2691.140 217.480 2691.400 ;
        RECT 217.220 489.300 217.480 489.560 ;
        RECT 1733.840 489.300 1734.100 489.560 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2691.430 17.320 2692.955 ;
        RECT 17.120 2691.110 17.380 2691.430 ;
        RECT 217.220 2691.110 217.480 2691.430 ;
        RECT 217.280 489.590 217.420 2691.110 ;
        RECT 1733.970 510.340 1734.250 514.000 ;
        RECT 1733.900 510.000 1734.250 510.340 ;
        RECT 1733.900 489.590 1734.040 510.000 ;
        RECT 217.220 489.270 217.480 489.590 ;
        RECT 1733.840 489.270 1734.100 489.590 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.800 2692.990 17.415 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 515.805 3029.145 516.895 3029.315 ;
      LAYER mcon ;
        RECT 516.725 3029.145 516.895 3029.315 ;
      LAYER met1 ;
        RECT 196.950 3029.300 197.270 3029.360 ;
        RECT 515.745 3029.300 516.035 3029.345 ;
        RECT 196.950 3029.160 516.035 3029.300 ;
        RECT 196.950 3029.100 197.270 3029.160 ;
        RECT 515.745 3029.115 516.035 3029.160 ;
        RECT 516.665 3029.300 516.955 3029.345 ;
        RECT 2519.490 3029.300 2519.810 3029.360 ;
        RECT 516.665 3029.160 2519.810 3029.300 ;
        RECT 516.665 3029.115 516.955 3029.160 ;
        RECT 2519.490 3029.100 2519.810 3029.160 ;
        RECT 18.930 2408.120 19.250 2408.180 ;
        RECT 196.950 2408.120 197.270 2408.180 ;
        RECT 18.930 2407.980 197.270 2408.120 ;
        RECT 18.930 2407.920 19.250 2407.980 ;
        RECT 196.950 2407.920 197.270 2407.980 ;
      LAYER via ;
        RECT 196.980 3029.100 197.240 3029.360 ;
        RECT 2519.520 3029.100 2519.780 3029.360 ;
        RECT 18.960 2407.920 19.220 2408.180 ;
        RECT 196.980 2407.920 197.240 2408.180 ;
      LAYER met2 ;
        RECT 196.980 3029.070 197.240 3029.390 ;
        RECT 2519.520 3029.070 2519.780 3029.390 ;
        RECT 197.040 2408.210 197.180 3029.070 ;
        RECT 2519.580 2969.405 2519.720 3029.070 ;
        RECT 2519.510 2969.035 2519.790 2969.405 ;
        RECT 18.960 2407.890 19.220 2408.210 ;
        RECT 196.980 2407.890 197.240 2408.210 ;
        RECT 19.020 2405.685 19.160 2407.890 ;
        RECT 18.950 2405.315 19.230 2405.685 ;
      LAYER via2 ;
        RECT 2519.510 2969.080 2519.790 2969.360 ;
        RECT 18.950 2405.360 19.230 2405.640 ;
      LAYER met3 ;
        RECT 2506.000 2969.370 2510.000 2969.520 ;
        RECT 2519.485 2969.370 2519.815 2969.385 ;
        RECT 2506.000 2969.070 2519.815 2969.370 ;
        RECT 2506.000 2968.920 2510.000 2969.070 ;
        RECT 2519.485 2969.055 2519.815 2969.070 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 18.925 2405.650 19.255 2405.665 ;
        RECT -4.800 2405.350 19.255 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 18.925 2405.335 19.255 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 348.750 3033.040 349.070 3033.100 ;
        RECT 2309.730 3033.040 2310.050 3033.100 ;
        RECT 348.750 3032.900 2310.050 3033.040 ;
        RECT 348.750 3032.840 349.070 3032.900 ;
        RECT 2309.730 3032.840 2310.050 3032.900 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 348.750 2125.240 349.070 2125.300 ;
        RECT 16.170 2125.100 349.070 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 348.750 2125.040 349.070 2125.100 ;
      LAYER via ;
        RECT 348.780 3032.840 349.040 3033.100 ;
        RECT 2309.760 3032.840 2310.020 3033.100 ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 348.780 2125.040 349.040 2125.300 ;
      LAYER met2 ;
        RECT 348.780 3032.810 349.040 3033.130 ;
        RECT 2309.760 3032.810 2310.020 3033.130 ;
        RECT 348.840 2125.330 348.980 3032.810 ;
        RECT 2309.820 3010.000 2309.960 3032.810 ;
        RECT 2309.820 3009.340 2310.170 3010.000 ;
        RECT 2309.890 3006.000 2310.170 3009.340 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 348.780 2125.010 349.040 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2400.970 510.340 2401.250 514.000 ;
        RECT 2400.900 510.000 2401.250 510.340 ;
        RECT 2400.900 482.645 2401.040 510.000 ;
        RECT 2400.830 482.275 2401.110 482.645 ;
      LAYER via2 ;
        RECT 2400.830 482.320 2401.110 482.600 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT -4.800 1830.750 3.370 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 3.070 1829.010 3.370 1830.750 ;
        RECT 355.390 1829.010 355.770 1829.020 ;
        RECT 3.070 1828.710 355.770 1829.010 ;
        RECT 355.390 1828.700 355.770 1828.710 ;
        RECT 355.390 482.610 355.770 482.620 ;
        RECT 2400.805 482.610 2401.135 482.625 ;
        RECT 355.390 482.310 2401.135 482.610 ;
        RECT 355.390 482.300 355.770 482.310 ;
        RECT 2400.805 482.295 2401.135 482.310 ;
      LAYER via3 ;
        RECT 355.420 1828.700 355.740 1829.020 ;
        RECT 355.420 482.300 355.740 482.620 ;
      LAYER met4 ;
        RECT 355.415 1828.695 355.745 1829.025 ;
        RECT 355.430 482.625 355.730 1828.695 ;
        RECT 355.415 482.295 355.745 482.625 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1556.250 3016.040 1556.570 3016.100 ;
        RECT 2763.290 3016.040 2763.610 3016.100 ;
        RECT 1556.250 3015.900 2763.610 3016.040 ;
        RECT 1556.250 3015.840 1556.570 3015.900 ;
        RECT 2763.290 3015.840 2763.610 3015.900 ;
        RECT 2763.290 676.160 2763.610 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2763.290 676.020 2901.150 676.160 ;
        RECT 2763.290 675.960 2763.610 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 1556.280 3015.840 1556.540 3016.100 ;
        RECT 2763.320 3015.840 2763.580 3016.100 ;
        RECT 2763.320 675.960 2763.580 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 1556.280 3015.810 1556.540 3016.130 ;
        RECT 2763.320 3015.810 2763.580 3016.130 ;
        RECT 1556.340 3010.000 1556.480 3015.810 ;
        RECT 1556.340 3009.340 1556.690 3010.000 ;
        RECT 1556.410 3006.000 1556.690 3009.340 ;
        RECT 2763.380 676.250 2763.520 3015.810 ;
        RECT 2763.320 675.930 2763.580 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 45.610 1587.360 45.930 1587.420 ;
        RECT 393.370 1587.360 393.690 1587.420 ;
        RECT 45.610 1587.220 393.690 1587.360 ;
        RECT 45.610 1587.160 45.930 1587.220 ;
        RECT 393.370 1587.160 393.690 1587.220 ;
        RECT 17.090 1544.860 17.410 1544.920 ;
        RECT 45.610 1544.860 45.930 1544.920 ;
        RECT 17.090 1544.720 45.930 1544.860 ;
        RECT 17.090 1544.660 17.410 1544.720 ;
        RECT 45.610 1544.660 45.930 1544.720 ;
      LAYER via ;
        RECT 45.640 1587.160 45.900 1587.420 ;
        RECT 393.400 1587.160 393.660 1587.420 ;
        RECT 17.120 1544.660 17.380 1544.920 ;
        RECT 45.640 1544.660 45.900 1544.920 ;
      LAYER met2 ;
        RECT 393.390 1591.355 393.670 1591.725 ;
        RECT 393.460 1587.450 393.600 1591.355 ;
        RECT 45.640 1587.130 45.900 1587.450 ;
        RECT 393.400 1587.130 393.660 1587.450 ;
        RECT 45.700 1544.950 45.840 1587.130 ;
        RECT 17.120 1544.630 17.380 1544.950 ;
        RECT 45.640 1544.630 45.900 1544.950 ;
        RECT 17.180 1544.125 17.320 1544.630 ;
        RECT 17.110 1543.755 17.390 1544.125 ;
      LAYER via2 ;
        RECT 393.390 1591.400 393.670 1591.680 ;
        RECT 17.110 1543.800 17.390 1544.080 ;
      LAYER met3 ;
        RECT 393.365 1591.690 393.695 1591.705 ;
        RECT 410.000 1591.690 414.000 1591.840 ;
        RECT 393.365 1591.390 414.000 1591.690 ;
        RECT 393.365 1591.375 393.695 1591.390 ;
        RECT 410.000 1591.240 414.000 1591.390 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 17.085 1544.090 17.415 1544.105 ;
        RECT -4.800 1543.790 17.415 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 17.085 1543.775 17.415 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1324.880 17.410 1324.940 ;
        RECT 341.850 1324.880 342.170 1324.940 ;
        RECT 17.090 1324.740 342.170 1324.880 ;
        RECT 17.090 1324.680 17.410 1324.740 ;
        RECT 341.850 1324.680 342.170 1324.740 ;
        RECT 341.850 503.100 342.170 503.160 ;
        RECT 1610.530 503.100 1610.850 503.160 ;
        RECT 341.850 502.960 1610.850 503.100 ;
        RECT 341.850 502.900 342.170 502.960 ;
        RECT 1610.530 502.900 1610.850 502.960 ;
      LAYER via ;
        RECT 17.120 1324.680 17.380 1324.940 ;
        RECT 341.880 1324.680 342.140 1324.940 ;
        RECT 341.880 502.900 342.140 503.160 ;
        RECT 1610.560 502.900 1610.820 503.160 ;
      LAYER met2 ;
        RECT 17.110 1328.195 17.390 1328.565 ;
        RECT 17.180 1324.970 17.320 1328.195 ;
        RECT 17.120 1324.650 17.380 1324.970 ;
        RECT 341.880 1324.650 342.140 1324.970 ;
        RECT 341.940 503.190 342.080 1324.650 ;
        RECT 1610.690 510.340 1610.970 514.000 ;
        RECT 1610.620 510.000 1610.970 510.340 ;
        RECT 1610.620 503.190 1610.760 510.000 ;
        RECT 341.880 502.870 342.140 503.190 ;
        RECT 1610.560 502.870 1610.820 503.190 ;
      LAYER via2 ;
        RECT 17.110 1328.240 17.390 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 17.085 1328.530 17.415 1328.545 ;
        RECT -4.800 1328.230 17.415 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 17.085 1328.215 17.415 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 362.550 3008.900 362.870 3008.960 ;
        RECT 579.670 3008.900 579.990 3008.960 ;
        RECT 362.550 3008.760 579.990 3008.900 ;
        RECT 362.550 3008.700 362.870 3008.760 ;
        RECT 579.670 3008.700 579.990 3008.760 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 362.550 1117.820 362.870 1117.880 ;
        RECT 15.710 1117.680 362.870 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 362.550 1117.620 362.870 1117.680 ;
      LAYER via ;
        RECT 362.580 3008.700 362.840 3008.960 ;
        RECT 579.700 3008.700 579.960 3008.960 ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 362.580 1117.620 362.840 1117.880 ;
      LAYER met2 ;
        RECT 362.580 3008.670 362.840 3008.990 ;
        RECT 579.700 3008.730 579.960 3008.990 ;
        RECT 580.290 3008.730 580.570 3010.000 ;
        RECT 579.700 3008.670 580.570 3008.730 ;
        RECT 362.640 1117.910 362.780 3008.670 ;
        RECT 579.760 3008.590 580.570 3008.670 ;
        RECT 580.290 3006.000 580.570 3008.590 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 362.580 1117.590 362.840 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 100.350 2970.480 100.670 2970.540 ;
        RECT 393.370 2970.480 393.690 2970.540 ;
        RECT 100.350 2970.340 393.690 2970.480 ;
        RECT 100.350 2970.280 100.670 2970.340 ;
        RECT 393.370 2970.280 393.690 2970.340 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 100.350 903.960 100.670 904.020 ;
        RECT 16.170 903.820 100.670 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 100.350 903.760 100.670 903.820 ;
      LAYER via ;
        RECT 100.380 2970.280 100.640 2970.540 ;
        RECT 393.400 2970.280 393.660 2970.540 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 100.380 903.760 100.640 904.020 ;
      LAYER met2 ;
        RECT 393.390 2978.555 393.670 2978.925 ;
        RECT 393.460 2970.570 393.600 2978.555 ;
        RECT 100.380 2970.250 100.640 2970.570 ;
        RECT 393.400 2970.250 393.660 2970.570 ;
        RECT 100.440 904.050 100.580 2970.250 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 100.380 903.730 100.640 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 393.390 2978.600 393.670 2978.880 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 393.365 2978.890 393.695 2978.905 ;
        RECT 410.000 2978.890 414.000 2979.040 ;
        RECT 393.365 2978.590 414.000 2978.890 ;
        RECT 393.365 2978.575 393.695 2978.590 ;
        RECT 410.000 2978.440 414.000 2978.590 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 96.745 514.165 96.915 515.015 ;
        RECT 48.445 512.805 48.615 513.655 ;
        RECT 96.285 512.805 96.455 513.995 ;
        RECT 193.345 513.825 193.515 515.695 ;
        RECT 254.985 515.525 255.615 515.695 ;
        RECT 255.445 515.185 255.615 515.525 ;
        RECT 283.045 513.825 283.215 515.355 ;
        RECT 330.885 513.825 331.055 514.675 ;
        RECT 400.805 512.295 400.975 512.635 ;
        RECT 399.885 512.125 400.975 512.295 ;
        RECT 434.845 511.955 435.015 512.295 ;
        RECT 434.845 511.785 435.475 511.955 ;
        RECT 517.645 511.785 517.815 512.635 ;
        RECT 579.745 510.765 579.915 511.955 ;
        RECT 690.145 511.615 690.315 511.955 ;
        RECT 628.045 510.765 628.215 511.615 ;
        RECT 689.685 511.445 690.315 511.615 ;
      LAYER mcon ;
        RECT 193.345 515.525 193.515 515.695 ;
        RECT 96.745 514.845 96.915 515.015 ;
        RECT 283.045 515.185 283.215 515.355 ;
        RECT 96.285 513.825 96.455 513.995 ;
        RECT 330.885 514.505 331.055 514.675 ;
        RECT 48.445 513.485 48.615 513.655 ;
        RECT 400.805 512.465 400.975 512.635 ;
        RECT 517.645 512.465 517.815 512.635 ;
        RECT 434.845 512.125 435.015 512.295 ;
        RECT 435.305 511.785 435.475 511.955 ;
        RECT 579.745 511.785 579.915 511.955 ;
        RECT 690.145 511.785 690.315 511.955 ;
        RECT 628.045 511.445 628.215 511.615 ;
      LAYER met1 ;
        RECT 17.550 679.220 17.870 679.280 ;
        RECT 45.610 679.220 45.930 679.280 ;
        RECT 17.550 679.080 45.930 679.220 ;
        RECT 17.550 679.020 17.870 679.080 ;
        RECT 45.610 679.020 45.930 679.080 ;
        RECT 193.285 515.680 193.575 515.725 ;
        RECT 254.925 515.680 255.215 515.725 ;
        RECT 193.285 515.540 255.215 515.680 ;
        RECT 193.285 515.495 193.575 515.540 ;
        RECT 254.925 515.495 255.215 515.540 ;
        RECT 255.385 515.340 255.675 515.385 ;
        RECT 282.985 515.340 283.275 515.385 ;
        RECT 255.385 515.200 283.275 515.340 ;
        RECT 255.385 515.155 255.675 515.200 ;
        RECT 282.985 515.155 283.275 515.200 ;
        RECT 96.685 515.000 96.975 515.045 ;
        RECT 96.685 514.860 149.340 515.000 ;
        RECT 96.685 514.815 96.975 514.860 ;
        RECT 96.685 514.320 96.975 514.365 ;
        RECT 96.300 514.180 96.975 514.320 ;
        RECT 96.300 514.025 96.440 514.180 ;
        RECT 96.685 514.135 96.975 514.180 ;
        RECT 96.225 513.795 96.515 514.025 ;
        RECT 149.200 513.980 149.340 514.860 ;
        RECT 330.825 514.660 331.115 514.705 ;
        RECT 330.825 514.520 356.340 514.660 ;
        RECT 330.825 514.475 331.115 514.520 ;
        RECT 193.285 513.980 193.575 514.025 ;
        RECT 149.200 513.840 193.575 513.980 ;
        RECT 193.285 513.795 193.575 513.840 ;
        RECT 282.985 513.980 283.275 514.025 ;
        RECT 330.825 513.980 331.115 514.025 ;
        RECT 282.985 513.840 331.115 513.980 ;
        RECT 282.985 513.795 283.275 513.840 ;
        RECT 330.825 513.795 331.115 513.840 ;
        RECT 45.610 513.640 45.930 513.700 ;
        RECT 48.385 513.640 48.675 513.685 ;
        RECT 45.610 513.500 48.675 513.640 ;
        RECT 45.610 513.440 45.930 513.500 ;
        RECT 48.385 513.455 48.675 513.500 ;
        RECT 48.385 512.960 48.675 513.005 ;
        RECT 96.225 512.960 96.515 513.005 ;
        RECT 48.385 512.820 96.515 512.960 ;
        RECT 48.385 512.775 48.675 512.820 ;
        RECT 96.225 512.775 96.515 512.820 ;
        RECT 356.200 512.280 356.340 514.520 ;
        RECT 400.745 512.620 401.035 512.665 ;
        RECT 517.585 512.620 517.875 512.665 ;
        RECT 400.745 512.480 435.000 512.620 ;
        RECT 400.745 512.435 401.035 512.480 ;
        RECT 434.860 512.325 435.000 512.480 ;
        RECT 517.585 512.480 545.400 512.620 ;
        RECT 517.585 512.435 517.875 512.480 ;
        RECT 399.825 512.280 400.115 512.325 ;
        RECT 356.200 512.140 400.115 512.280 ;
        RECT 399.825 512.095 400.115 512.140 ;
        RECT 434.785 512.095 435.075 512.325 ;
        RECT 435.245 511.940 435.535 511.985 ;
        RECT 435.245 511.800 517.340 511.940 ;
        RECT 435.245 511.755 435.535 511.800 ;
        RECT 517.200 511.600 517.340 511.800 ;
        RECT 517.585 511.755 517.875 511.985 ;
        RECT 545.260 511.940 545.400 512.480 ;
        RECT 745.270 512.280 745.590 512.340 ;
        RECT 714.080 512.140 745.590 512.280 ;
        RECT 579.685 511.940 579.975 511.985 ;
        RECT 545.260 511.800 579.975 511.940 ;
        RECT 579.685 511.755 579.975 511.800 ;
        RECT 690.085 511.940 690.375 511.985 ;
        RECT 714.080 511.940 714.220 512.140 ;
        RECT 745.270 512.080 745.590 512.140 ;
        RECT 690.085 511.800 714.220 511.940 ;
        RECT 690.085 511.755 690.375 511.800 ;
        RECT 517.660 511.600 517.800 511.755 ;
        RECT 517.200 511.460 517.800 511.600 ;
        RECT 627.985 511.600 628.275 511.645 ;
        RECT 689.625 511.600 689.915 511.645 ;
        RECT 627.985 511.460 689.915 511.600 ;
        RECT 627.985 511.415 628.275 511.460 ;
        RECT 689.625 511.415 689.915 511.460 ;
        RECT 579.685 510.920 579.975 510.965 ;
        RECT 627.985 510.920 628.275 510.965 ;
        RECT 579.685 510.780 628.275 510.920 ;
        RECT 579.685 510.735 579.975 510.780 ;
        RECT 627.985 510.735 628.275 510.780 ;
      LAYER via ;
        RECT 17.580 679.020 17.840 679.280 ;
        RECT 45.640 679.020 45.900 679.280 ;
        RECT 45.640 513.440 45.900 513.700 ;
        RECT 745.300 512.080 745.560 512.340 ;
      LAYER met2 ;
        RECT 17.570 681.515 17.850 681.885 ;
        RECT 17.640 679.310 17.780 681.515 ;
        RECT 17.580 678.990 17.840 679.310 ;
        RECT 45.640 678.990 45.900 679.310 ;
        RECT 45.700 513.730 45.840 678.990 ;
        RECT 45.640 513.410 45.900 513.730 ;
        RECT 745.890 512.450 746.170 514.000 ;
        RECT 745.360 512.370 746.170 512.450 ;
        RECT 745.300 512.310 746.170 512.370 ;
        RECT 745.300 512.050 745.560 512.310 ;
        RECT 745.890 510.000 746.170 512.310 ;
      LAYER via2 ;
        RECT 17.570 681.560 17.850 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.545 681.850 17.875 681.865 ;
        RECT -4.800 681.550 17.875 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 17.545 681.535 17.875 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.650 1732.200 79.970 1732.260 ;
        RECT 393.370 1732.200 393.690 1732.260 ;
        RECT 79.650 1732.060 393.690 1732.200 ;
        RECT 79.650 1732.000 79.970 1732.060 ;
        RECT 393.370 1732.000 393.690 1732.060 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 79.650 469.100 79.970 469.160 ;
        RECT 17.090 468.960 79.970 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 79.650 468.900 79.970 468.960 ;
      LAYER via ;
        RECT 79.680 1732.000 79.940 1732.260 ;
        RECT 393.400 1732.000 393.660 1732.260 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 79.680 468.900 79.940 469.160 ;
      LAYER met2 ;
        RECT 393.390 1736.875 393.670 1737.245 ;
        RECT 393.460 1732.290 393.600 1736.875 ;
        RECT 79.680 1731.970 79.940 1732.290 ;
        RECT 393.400 1731.970 393.660 1732.290 ;
        RECT 79.740 469.190 79.880 1731.970 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 79.680 468.870 79.940 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 393.390 1736.920 393.670 1737.200 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 393.365 1737.210 393.695 1737.225 ;
        RECT 410.000 1737.210 414.000 1737.360 ;
        RECT 393.365 1736.910 414.000 1737.210 ;
        RECT 393.365 1736.895 393.695 1736.910 ;
        RECT 410.000 1736.760 414.000 1736.910 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 3018.760 355.510 3018.820 ;
        RECT 480.770 3018.760 481.090 3018.820 ;
        RECT 355.190 3018.620 481.090 3018.760 ;
        RECT 355.190 3018.560 355.510 3018.620 ;
        RECT 480.770 3018.560 481.090 3018.620 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 355.190 255.240 355.510 255.300 ;
        RECT 17.090 255.100 355.510 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 355.190 255.040 355.510 255.100 ;
      LAYER via ;
        RECT 355.220 3018.560 355.480 3018.820 ;
        RECT 480.800 3018.560 481.060 3018.820 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 355.220 255.040 355.480 255.300 ;
      LAYER met2 ;
        RECT 355.220 3018.530 355.480 3018.850 ;
        RECT 480.800 3018.530 481.060 3018.850 ;
        RECT 355.280 255.330 355.420 3018.530 ;
        RECT 480.860 3010.000 481.000 3018.530 ;
        RECT 480.860 3009.340 481.210 3010.000 ;
        RECT 480.930 3006.000 481.210 3009.340 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 355.220 255.010 355.480 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2015.080 2519.810 2015.140 ;
        RECT 2568.710 2015.080 2569.030 2015.140 ;
        RECT 2519.490 2014.940 2569.030 2015.080 ;
        RECT 2519.490 2014.880 2519.810 2014.940 ;
        RECT 2568.710 2014.880 2569.030 2014.940 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 2568.710 41.380 2569.030 41.440 ;
        RECT 17.090 41.240 2569.030 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 2568.710 41.180 2569.030 41.240 ;
      LAYER via ;
        RECT 2519.520 2014.880 2519.780 2015.140 ;
        RECT 2568.740 2014.880 2569.000 2015.140 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 2568.740 41.180 2569.000 41.440 ;
      LAYER met2 ;
        RECT 2519.510 2018.395 2519.790 2018.765 ;
        RECT 2519.580 2015.170 2519.720 2018.395 ;
        RECT 2519.520 2014.850 2519.780 2015.170 ;
        RECT 2568.740 2014.850 2569.000 2015.170 ;
        RECT 2568.800 41.470 2568.940 2014.850 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 2568.740 41.150 2569.000 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 2519.510 2018.440 2519.790 2018.720 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 2506.000 2018.730 2510.000 2018.880 ;
        RECT 2519.485 2018.730 2519.815 2018.745 ;
        RECT 2506.000 2018.430 2519.815 2018.730 ;
        RECT 2506.000 2018.280 2510.000 2018.430 ;
        RECT 2519.485 2018.415 2519.815 2018.430 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2704.430 906.595 2704.710 906.965 ;
        RECT 2704.500 905.605 2704.640 906.595 ;
        RECT 2704.430 905.235 2704.710 905.605 ;
      LAYER via2 ;
        RECT 2704.430 906.640 2704.710 906.920 ;
        RECT 2704.430 905.280 2704.710 905.560 ;
      LAYER met3 ;
        RECT 2509.110 1140.850 2509.490 1140.860 ;
        RECT 2535.790 1140.850 2536.170 1140.860 ;
        RECT 2509.110 1140.550 2536.170 1140.850 ;
        RECT 2509.110 1140.540 2509.490 1140.550 ;
        RECT 2535.790 1140.540 2536.170 1140.550 ;
        RECT 412.430 1137.140 412.810 1137.460 ;
        RECT 2557.870 1137.450 2558.250 1137.460 ;
        RECT 2611.230 1137.450 2611.610 1137.460 ;
        RECT 2557.870 1137.150 2611.610 1137.450 ;
        RECT 2557.870 1137.140 2558.250 1137.150 ;
        RECT 2611.230 1137.140 2611.610 1137.150 ;
        RECT 412.470 1134.880 412.770 1137.140 ;
        RECT 410.000 1134.280 414.000 1134.880 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 2656.310 906.930 2656.690 906.940 ;
        RECT 2704.405 906.930 2704.735 906.945 ;
        RECT 2656.310 906.630 2704.735 906.930 ;
        RECT 2656.310 906.620 2656.690 906.630 ;
        RECT 2704.405 906.615 2704.735 906.630 ;
        RECT 2611.230 905.570 2611.610 905.580 ;
        RECT 2704.405 905.570 2704.735 905.585 ;
        RECT 2916.710 905.570 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2611.230 905.270 2622.610 905.570 ;
        RECT 2611.230 905.260 2611.610 905.270 ;
        RECT 2622.310 904.890 2622.610 905.270 ;
        RECT 2704.405 905.270 2767.050 905.570 ;
        RECT 2704.405 905.255 2704.735 905.270 ;
        RECT 2656.310 904.890 2656.690 904.900 ;
        RECT 2622.310 904.590 2656.690 904.890 ;
        RECT 2766.750 904.890 2767.050 905.270 ;
        RECT 2863.350 905.270 2917.010 905.570 ;
        RECT 2766.750 904.590 2814.890 904.890 ;
        RECT 2656.310 904.580 2656.690 904.590 ;
        RECT 2814.590 904.210 2814.890 904.590 ;
        RECT 2863.350 904.210 2863.650 905.270 ;
        RECT 2814.590 903.910 2863.650 904.210 ;
      LAYER via3 ;
        RECT 2509.140 1140.540 2509.460 1140.860 ;
        RECT 2535.820 1140.540 2536.140 1140.860 ;
        RECT 412.460 1137.140 412.780 1137.460 ;
        RECT 2557.900 1137.140 2558.220 1137.460 ;
        RECT 2611.260 1137.140 2611.580 1137.460 ;
        RECT 2656.340 906.620 2656.660 906.940 ;
        RECT 2611.260 905.260 2611.580 905.580 ;
        RECT 2656.340 904.580 2656.660 904.900 ;
      LAYER met4 ;
        RECT 2508.710 1140.110 2509.890 1141.290 ;
        RECT 2535.815 1140.535 2536.145 1140.865 ;
        RECT 412.030 1136.710 413.210 1137.890 ;
        RECT 2535.830 1134.490 2536.130 1140.535 ;
        RECT 2557.895 1137.135 2558.225 1137.465 ;
        RECT 2611.255 1137.135 2611.585 1137.465 ;
        RECT 2557.910 1134.490 2558.210 1137.135 ;
        RECT 2535.390 1133.310 2536.570 1134.490 ;
        RECT 2557.470 1133.310 2558.650 1134.490 ;
        RECT 2611.270 905.585 2611.570 1137.135 ;
        RECT 2656.335 906.615 2656.665 906.945 ;
        RECT 2611.255 905.255 2611.585 905.585 ;
        RECT 2656.350 904.905 2656.650 906.615 ;
        RECT 2656.335 904.575 2656.665 904.905 ;
      LAYER met5 ;
        RECT 495.540 1139.900 627.780 1141.500 ;
        RECT 411.820 1136.500 483.340 1138.100 ;
        RECT 481.740 1134.700 483.340 1136.500 ;
        RECT 495.540 1134.700 497.140 1139.900 ;
        RECT 481.740 1133.100 497.140 1134.700 ;
        RECT 626.180 1134.700 627.780 1139.900 ;
        RECT 639.980 1139.900 724.380 1141.500 ;
        RECT 639.980 1134.700 641.580 1139.900 ;
        RECT 626.180 1133.100 641.580 1134.700 ;
        RECT 722.780 1134.700 724.380 1139.900 ;
        RECT 736.580 1139.900 820.980 1141.500 ;
        RECT 736.580 1134.700 738.180 1139.900 ;
        RECT 722.780 1133.100 738.180 1134.700 ;
        RECT 819.380 1134.700 820.980 1139.900 ;
        RECT 833.180 1139.900 917.580 1141.500 ;
        RECT 833.180 1134.700 834.780 1139.900 ;
        RECT 819.380 1133.100 834.780 1134.700 ;
        RECT 915.980 1134.700 917.580 1139.900 ;
        RECT 929.780 1139.900 980.140 1141.500 ;
        RECT 929.780 1134.700 931.380 1139.900 ;
        RECT 915.980 1133.100 931.380 1134.700 ;
        RECT 978.540 1134.700 980.140 1139.900 ;
        RECT 999.700 1139.900 1049.140 1141.500 ;
        RECT 999.700 1134.700 1001.300 1139.900 ;
        RECT 978.540 1133.100 1001.300 1134.700 ;
        RECT 1047.540 1134.700 1049.140 1139.900 ;
        RECT 1096.300 1139.900 1145.740 1141.500 ;
        RECT 1096.300 1134.700 1097.900 1139.900 ;
        RECT 1047.540 1133.100 1097.900 1134.700 ;
        RECT 1144.140 1134.700 1145.740 1139.900 ;
        RECT 1192.900 1139.900 1242.340 1141.500 ;
        RECT 1192.900 1134.700 1194.500 1139.900 ;
        RECT 1144.140 1133.100 1194.500 1134.700 ;
        RECT 1240.740 1134.700 1242.340 1139.900 ;
        RECT 1289.500 1139.900 1338.940 1141.500 ;
        RECT 1289.500 1134.700 1291.100 1139.900 ;
        RECT 1240.740 1133.100 1291.100 1134.700 ;
        RECT 1337.340 1134.700 1338.940 1139.900 ;
        RECT 1386.100 1139.900 1435.540 1141.500 ;
        RECT 1386.100 1134.700 1387.700 1139.900 ;
        RECT 1337.340 1133.100 1387.700 1134.700 ;
        RECT 1433.940 1134.700 1435.540 1139.900 ;
        RECT 1482.700 1139.900 1532.140 1141.500 ;
        RECT 1482.700 1134.700 1484.300 1139.900 ;
        RECT 1433.940 1133.100 1484.300 1134.700 ;
        RECT 1530.540 1134.700 1532.140 1139.900 ;
        RECT 1579.300 1139.900 1628.740 1141.500 ;
        RECT 1579.300 1134.700 1580.900 1139.900 ;
        RECT 1530.540 1133.100 1580.900 1134.700 ;
        RECT 1627.140 1134.700 1628.740 1139.900 ;
        RECT 1675.900 1139.900 1725.340 1141.500 ;
        RECT 1675.900 1134.700 1677.500 1139.900 ;
        RECT 1627.140 1133.100 1677.500 1134.700 ;
        RECT 1723.740 1134.700 1725.340 1139.900 ;
        RECT 1772.500 1139.900 1821.940 1141.500 ;
        RECT 1772.500 1134.700 1774.100 1139.900 ;
        RECT 1723.740 1133.100 1774.100 1134.700 ;
        RECT 1820.340 1134.700 1821.940 1139.900 ;
        RECT 1869.100 1139.900 1918.540 1141.500 ;
        RECT 1869.100 1134.700 1870.700 1139.900 ;
        RECT 1820.340 1133.100 1870.700 1134.700 ;
        RECT 1916.940 1134.700 1918.540 1139.900 ;
        RECT 1965.700 1139.900 2015.140 1141.500 ;
        RECT 1965.700 1134.700 1967.300 1139.900 ;
        RECT 1916.940 1133.100 1967.300 1134.700 ;
        RECT 2013.540 1134.700 2015.140 1139.900 ;
        RECT 2062.300 1139.900 2111.740 1141.500 ;
        RECT 2062.300 1134.700 2063.900 1139.900 ;
        RECT 2013.540 1133.100 2063.900 1134.700 ;
        RECT 2110.140 1134.700 2111.740 1139.900 ;
        RECT 2158.900 1139.900 2208.340 1141.500 ;
        RECT 2158.900 1134.700 2160.500 1139.900 ;
        RECT 2110.140 1133.100 2160.500 1134.700 ;
        RECT 2206.740 1134.700 2208.340 1139.900 ;
        RECT 2255.500 1139.900 2304.940 1141.500 ;
        RECT 2255.500 1134.700 2257.100 1139.900 ;
        RECT 2206.740 1133.100 2257.100 1134.700 ;
        RECT 2303.340 1134.700 2304.940 1139.900 ;
        RECT 2352.100 1139.900 2361.060 1141.500 ;
        RECT 2352.100 1134.700 2353.700 1139.900 ;
        RECT 2359.460 1138.100 2361.060 1139.900 ;
        RECT 2407.300 1139.900 2510.100 1141.500 ;
        RECT 2407.300 1138.100 2408.900 1139.900 ;
        RECT 2359.460 1136.500 2408.900 1138.100 ;
        RECT 2303.340 1133.100 2353.700 1134.700 ;
        RECT 2406.380 1133.100 2408.900 1136.500 ;
        RECT 2535.180 1133.100 2558.860 1134.700 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2408.170 3017.060 2408.490 3017.120 ;
        RECT 2659.790 3017.060 2660.110 3017.120 ;
        RECT 2408.170 3016.920 2660.110 3017.060 ;
        RECT 2408.170 3016.860 2408.490 3016.920 ;
        RECT 2659.790 3016.860 2660.110 3016.920 ;
        RECT 2659.790 1145.360 2660.110 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2659.790 1145.220 2901.150 1145.360 ;
        RECT 2659.790 1145.160 2660.110 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2408.200 3016.860 2408.460 3017.120 ;
        RECT 2659.820 3016.860 2660.080 3017.120 ;
        RECT 2659.820 1145.160 2660.080 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2408.200 3016.830 2408.460 3017.150 ;
        RECT 2659.820 3016.830 2660.080 3017.150 ;
        RECT 2408.260 3010.000 2408.400 3016.830 ;
        RECT 2408.260 3009.340 2408.610 3010.000 ;
        RECT 2408.330 3006.000 2408.610 3009.340 ;
        RECT 2659.880 1145.450 2660.020 3016.830 ;
        RECT 2659.820 1145.130 2660.080 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 3031.000 1049.650 3031.060 ;
        RECT 2770.190 3031.000 2770.510 3031.060 ;
        RECT 1049.330 3030.860 2770.510 3031.000 ;
        RECT 1049.330 3030.800 1049.650 3030.860 ;
        RECT 2770.190 3030.800 2770.510 3030.860 ;
        RECT 2770.190 1379.960 2770.510 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2770.190 1379.820 2901.150 1379.960 ;
        RECT 2770.190 1379.760 2770.510 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 1049.360 3030.800 1049.620 3031.060 ;
        RECT 2770.220 3030.800 2770.480 3031.060 ;
        RECT 2770.220 1379.760 2770.480 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 1049.360 3030.770 1049.620 3031.090 ;
        RECT 2770.220 3030.770 2770.480 3031.090 ;
        RECT 1049.420 3010.000 1049.560 3030.770 ;
        RECT 1049.420 3009.340 1049.770 3010.000 ;
        RECT 1049.490 3006.000 1049.770 3009.340 ;
        RECT 2770.280 1380.050 2770.420 3030.770 ;
        RECT 2770.220 1379.730 2770.480 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2508.450 2998.360 2508.770 2998.420 ;
        RECT 2570.090 2998.360 2570.410 2998.420 ;
        RECT 2508.450 2998.220 2570.410 2998.360 ;
        RECT 2508.450 2998.160 2508.770 2998.220 ;
        RECT 2570.090 2998.160 2570.410 2998.220 ;
        RECT 2570.090 1614.560 2570.410 1614.620 ;
        RECT 2900.830 1614.560 2901.150 1614.620 ;
        RECT 2570.090 1614.420 2901.150 1614.560 ;
        RECT 2570.090 1614.360 2570.410 1614.420 ;
        RECT 2900.830 1614.360 2901.150 1614.420 ;
      LAYER via ;
        RECT 2508.480 2998.160 2508.740 2998.420 ;
        RECT 2570.120 2998.160 2570.380 2998.420 ;
        RECT 2570.120 1614.360 2570.380 1614.620 ;
        RECT 2900.860 1614.360 2901.120 1614.620 ;
      LAYER met2 ;
        RECT 2506.770 3006.690 2507.050 3010.000 ;
        RECT 2506.770 3006.550 2508.680 3006.690 ;
        RECT 2506.770 3006.000 2507.050 3006.550 ;
        RECT 2508.540 2998.450 2508.680 3006.550 ;
        RECT 2508.480 2998.130 2508.740 2998.450 ;
        RECT 2570.120 2998.130 2570.380 2998.450 ;
        RECT 2570.180 1614.650 2570.320 2998.130 ;
        RECT 2570.120 1614.330 2570.380 1614.650 ;
        RECT 2900.860 1614.330 2901.120 1614.650 ;
        RECT 2900.920 1613.485 2901.060 1614.330 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2570.550 1842.700 2570.870 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2570.550 1842.560 2901.150 1842.700 ;
        RECT 2570.550 1842.500 2570.870 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
        RECT 1462.410 503.440 1462.730 503.500 ;
        RECT 2570.550 503.440 2570.870 503.500 ;
        RECT 1462.410 503.300 2570.870 503.440 ;
        RECT 1462.410 503.240 1462.730 503.300 ;
        RECT 2570.550 503.240 2570.870 503.300 ;
      LAYER via ;
        RECT 2570.580 1842.500 2570.840 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
        RECT 1462.440 503.240 1462.700 503.500 ;
        RECT 2570.580 503.240 2570.840 503.500 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2570.580 1842.470 2570.840 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 1462.570 510.340 1462.850 514.000 ;
        RECT 1462.500 510.000 1462.850 510.340 ;
        RECT 1462.500 503.530 1462.640 510.000 ;
        RECT 2570.640 503.530 2570.780 1842.470 ;
        RECT 1462.440 503.210 1462.700 503.530 ;
        RECT 2570.580 503.210 2570.840 503.530 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2507.605 2997.865 2507.775 3018.095 ;
      LAYER mcon ;
        RECT 2507.605 3017.925 2507.775 3018.095 ;
      LAYER met1 ;
        RECT 2111.930 3018.080 2112.250 3018.140 ;
        RECT 2507.545 3018.080 2507.835 3018.125 ;
        RECT 2111.930 3017.940 2507.835 3018.080 ;
        RECT 2111.930 3017.880 2112.250 3017.940 ;
        RECT 2507.545 3017.895 2507.835 3017.940 ;
        RECT 2507.545 2998.020 2507.835 2998.065 ;
        RECT 2901.750 2998.020 2902.070 2998.080 ;
        RECT 2507.545 2997.880 2902.070 2998.020 ;
        RECT 2507.545 2997.835 2507.835 2997.880 ;
        RECT 2901.750 2997.820 2902.070 2997.880 ;
      LAYER via ;
        RECT 2111.960 3017.880 2112.220 3018.140 ;
        RECT 2901.780 2997.820 2902.040 2998.080 ;
      LAYER met2 ;
        RECT 2111.960 3017.850 2112.220 3018.170 ;
        RECT 2112.020 3010.000 2112.160 3017.850 ;
        RECT 2112.020 3009.340 2112.370 3010.000 ;
        RECT 2112.090 3006.000 2112.370 3009.340 ;
        RECT 2901.780 2997.790 2902.040 2998.110 ;
        RECT 2901.840 2082.685 2901.980 2997.790 ;
        RECT 2901.770 2082.315 2902.050 2082.685 ;
      LAYER via2 ;
        RECT 2901.770 2082.360 2902.050 2082.640 ;
      LAYER met3 ;
        RECT 2901.745 2082.650 2902.075 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2901.745 2082.350 2924.800 2082.650 ;
        RECT 2901.745 2082.335 2902.075 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 883.345 482.885 884.435 483.055 ;
        RECT 1060.905 482.885 1062.455 483.055 ;
        RECT 1782.185 482.885 1783.275 483.055 ;
        RECT 2563.725 482.885 2564.815 483.055 ;
      LAYER mcon ;
        RECT 884.265 482.885 884.435 483.055 ;
        RECT 1062.285 482.885 1062.455 483.055 ;
        RECT 1783.105 482.885 1783.275 483.055 ;
        RECT 2564.645 482.885 2564.815 483.055 ;
      LAYER met1 ;
        RECT 2825.390 2311.900 2825.710 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2825.390 2311.760 2901.150 2311.900 ;
        RECT 2825.390 2311.700 2825.710 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 844.170 483.040 844.490 483.100 ;
        RECT 883.285 483.040 883.575 483.085 ;
        RECT 844.170 482.900 883.575 483.040 ;
        RECT 844.170 482.840 844.490 482.900 ;
        RECT 883.285 482.855 883.575 482.900 ;
        RECT 884.205 483.040 884.495 483.085 ;
        RECT 1060.845 483.040 1061.135 483.085 ;
        RECT 884.205 482.900 1061.135 483.040 ;
        RECT 884.205 482.855 884.495 482.900 ;
        RECT 1060.845 482.855 1061.135 482.900 ;
        RECT 1062.225 483.040 1062.515 483.085 ;
        RECT 1782.125 483.040 1782.415 483.085 ;
        RECT 1062.225 482.900 1782.415 483.040 ;
        RECT 1062.225 482.855 1062.515 482.900 ;
        RECT 1782.125 482.855 1782.415 482.900 ;
        RECT 1783.045 483.040 1783.335 483.085 ;
        RECT 2563.665 483.040 2563.955 483.085 ;
        RECT 1783.045 482.900 2563.955 483.040 ;
        RECT 1783.045 482.855 1783.335 482.900 ;
        RECT 2563.665 482.855 2563.955 482.900 ;
        RECT 2564.585 483.040 2564.875 483.085 ;
        RECT 2825.390 483.040 2825.710 483.100 ;
        RECT 2564.585 482.900 2825.710 483.040 ;
        RECT 2564.585 482.855 2564.875 482.900 ;
        RECT 2825.390 482.840 2825.710 482.900 ;
      LAYER via ;
        RECT 2825.420 2311.700 2825.680 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 844.200 482.840 844.460 483.100 ;
        RECT 2825.420 482.840 2825.680 483.100 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2825.420 2311.670 2825.680 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 844.330 510.340 844.610 514.000 ;
        RECT 844.260 510.000 844.610 510.340 ;
        RECT 844.260 483.130 844.400 510.000 ;
        RECT 2825.480 483.130 2825.620 2311.670 ;
        RECT 844.200 482.810 844.460 483.130 ;
        RECT 2825.420 482.810 2825.680 483.130 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2765.590 146.100 2765.910 146.160 ;
        RECT 2801.010 146.100 2801.330 146.160 ;
        RECT 2765.590 145.960 2801.330 146.100 ;
        RECT 2765.590 145.900 2765.910 145.960 ;
        RECT 2801.010 145.900 2801.330 145.960 ;
      LAYER via ;
        RECT 2765.620 145.900 2765.880 146.160 ;
        RECT 2801.040 145.900 2801.300 146.160 ;
      LAYER met2 ;
        RECT 926.070 3029.555 926.350 3029.925 ;
        RECT 926.140 3010.000 926.280 3029.555 ;
        RECT 926.140 3009.340 926.490 3010.000 ;
        RECT 926.210 3006.000 926.490 3009.340 ;
        RECT 2801.030 146.355 2801.310 146.725 ;
        RECT 2801.100 146.190 2801.240 146.355 ;
        RECT 2765.620 146.045 2765.880 146.190 ;
        RECT 2765.610 145.675 2765.890 146.045 ;
        RECT 2801.040 145.870 2801.300 146.190 ;
      LAYER via2 ;
        RECT 926.070 3029.600 926.350 3029.880 ;
        RECT 2801.030 146.400 2801.310 146.680 ;
        RECT 2765.610 145.720 2765.890 146.000 ;
      LAYER met3 ;
        RECT 926.045 3029.890 926.375 3029.905 ;
        RECT 2583.630 3029.890 2584.010 3029.900 ;
        RECT 926.045 3029.590 2584.010 3029.890 ;
        RECT 926.045 3029.575 926.375 3029.590 ;
        RECT 2583.630 3029.580 2584.010 3029.590 ;
        RECT 2801.005 146.690 2801.335 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2670.150 146.390 2719.210 146.690 ;
        RECT 2583.630 145.330 2584.010 145.340 ;
        RECT 2670.150 145.330 2670.450 146.390 ;
        RECT 2718.910 146.010 2719.210 146.390 ;
        RECT 2801.005 146.390 2863.650 146.690 ;
        RECT 2801.005 146.375 2801.335 146.390 ;
        RECT 2765.585 146.010 2765.915 146.025 ;
        RECT 2718.910 145.710 2765.915 146.010 ;
        RECT 2765.585 145.695 2765.915 145.710 ;
        RECT 2583.630 145.030 2670.450 145.330 ;
        RECT 2863.350 145.330 2863.650 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 145.330 2917.010 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2863.350 145.030 2917.010 145.330 ;
        RECT 2583.630 145.020 2584.010 145.030 ;
      LAYER via3 ;
        RECT 2583.660 3029.580 2583.980 3029.900 ;
        RECT 2583.660 145.020 2583.980 145.340 ;
      LAYER met4 ;
        RECT 2583.655 3029.575 2583.985 3029.905 ;
        RECT 2583.670 145.345 2583.970 3029.575 ;
        RECT 2583.655 145.015 2583.985 145.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 826.690 3030.660 827.010 3030.720 ;
        RECT 2542.490 3030.660 2542.810 3030.720 ;
        RECT 826.690 3030.520 2542.810 3030.660 ;
        RECT 826.690 3030.460 827.010 3030.520 ;
        RECT 2542.490 3030.460 2542.810 3030.520 ;
        RECT 2542.490 2497.540 2542.810 2497.600 ;
        RECT 2900.830 2497.540 2901.150 2497.600 ;
        RECT 2542.490 2497.400 2901.150 2497.540 ;
        RECT 2542.490 2497.340 2542.810 2497.400 ;
        RECT 2900.830 2497.340 2901.150 2497.400 ;
      LAYER via ;
        RECT 826.720 3030.460 826.980 3030.720 ;
        RECT 2542.520 3030.460 2542.780 3030.720 ;
        RECT 2542.520 2497.340 2542.780 2497.600 ;
        RECT 2900.860 2497.340 2901.120 2497.600 ;
      LAYER met2 ;
        RECT 826.720 3030.430 826.980 3030.750 ;
        RECT 2542.520 3030.430 2542.780 3030.750 ;
        RECT 826.780 3010.000 826.920 3030.430 ;
        RECT 826.780 3009.340 827.130 3010.000 ;
        RECT 826.850 3006.000 827.130 3009.340 ;
        RECT 2542.580 2497.630 2542.720 3030.430 ;
        RECT 2542.520 2497.310 2542.780 2497.630 ;
        RECT 2900.860 2497.310 2901.120 2497.630 ;
        RECT 2900.920 2493.405 2901.060 2497.310 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1061.825 482.205 1062.455 482.375 ;
      LAYER mcon ;
        RECT 1062.285 482.205 1062.455 482.375 ;
      LAYER met1 ;
        RECT 2563.190 2725.680 2563.510 2725.740 ;
        RECT 2899.450 2725.680 2899.770 2725.740 ;
        RECT 2563.190 2725.540 2899.770 2725.680 ;
        RECT 2563.190 2725.480 2563.510 2725.540 ;
        RECT 2899.450 2725.480 2899.770 2725.540 ;
        RECT 955.490 482.360 955.810 482.420 ;
        RECT 1061.765 482.360 1062.055 482.405 ;
        RECT 955.490 482.220 1062.055 482.360 ;
        RECT 955.490 482.160 955.810 482.220 ;
        RECT 1061.765 482.175 1062.055 482.220 ;
        RECT 1062.225 482.360 1062.515 482.405 ;
        RECT 2563.190 482.360 2563.510 482.420 ;
        RECT 1062.225 482.220 1739.100 482.360 ;
        RECT 1062.225 482.175 1062.515 482.220 ;
        RECT 1738.960 482.020 1739.100 482.220 ;
        RECT 1783.120 482.220 2563.510 482.360 ;
        RECT 1783.120 482.020 1783.260 482.220 ;
        RECT 2563.190 482.160 2563.510 482.220 ;
        RECT 1738.960 481.880 1783.260 482.020 ;
      LAYER via ;
        RECT 2563.220 2725.480 2563.480 2725.740 ;
        RECT 2899.480 2725.480 2899.740 2725.740 ;
        RECT 955.520 482.160 955.780 482.420 ;
        RECT 2563.220 482.160 2563.480 482.420 ;
      LAYER met2 ;
        RECT 2899.470 2727.635 2899.750 2728.005 ;
        RECT 2899.540 2725.770 2899.680 2727.635 ;
        RECT 2563.220 2725.450 2563.480 2725.770 ;
        RECT 2899.480 2725.450 2899.740 2725.770 ;
        RECT 955.650 510.340 955.930 514.000 ;
        RECT 955.580 510.000 955.930 510.340 ;
        RECT 955.580 482.450 955.720 510.000 ;
        RECT 2563.280 482.450 2563.420 2725.450 ;
        RECT 955.520 482.130 955.780 482.450 ;
        RECT 2563.220 482.130 2563.480 482.450 ;
      LAYER via2 ;
        RECT 2899.470 2727.680 2899.750 2727.960 ;
      LAYER met3 ;
        RECT 2899.445 2727.970 2899.775 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2899.445 2727.670 2924.800 2727.970 ;
        RECT 2899.445 2727.655 2899.775 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2556.290 2960.280 2556.610 2960.340 ;
        RECT 2899.450 2960.280 2899.770 2960.340 ;
        RECT 2556.290 2960.140 2899.770 2960.280 ;
        RECT 2556.290 2960.080 2556.610 2960.140 ;
        RECT 2899.450 2960.080 2899.770 2960.140 ;
        RECT 1944.490 502.420 1944.810 502.480 ;
        RECT 2556.290 502.420 2556.610 502.480 ;
        RECT 1944.490 502.280 2556.610 502.420 ;
        RECT 1944.490 502.220 1944.810 502.280 ;
        RECT 2556.290 502.220 2556.610 502.280 ;
      LAYER via ;
        RECT 2556.320 2960.080 2556.580 2960.340 ;
        RECT 2899.480 2960.080 2899.740 2960.340 ;
        RECT 1944.520 502.220 1944.780 502.480 ;
        RECT 2556.320 502.220 2556.580 502.480 ;
      LAYER met2 ;
        RECT 2899.470 2962.235 2899.750 2962.605 ;
        RECT 2899.540 2960.370 2899.680 2962.235 ;
        RECT 2556.320 2960.050 2556.580 2960.370 ;
        RECT 2899.480 2960.050 2899.740 2960.370 ;
        RECT 1944.650 510.340 1944.930 514.000 ;
        RECT 1944.580 510.000 1944.930 510.340 ;
        RECT 1944.580 502.510 1944.720 510.000 ;
        RECT 2556.380 502.510 2556.520 2960.050 ;
        RECT 1944.520 502.190 1944.780 502.510 ;
        RECT 2556.320 502.190 2556.580 502.510 ;
      LAYER via2 ;
        RECT 2899.470 2962.280 2899.750 2962.560 ;
      LAYER met3 ;
        RECT 2899.445 2962.570 2899.775 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2899.445 2962.270 2924.800 2962.570 ;
        RECT 2899.445 2962.255 2899.775 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2576.990 3194.880 2577.310 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2576.990 3194.740 2901.150 3194.880 ;
        RECT 2576.990 3194.680 2577.310 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
        RECT 2018.090 501.740 2018.410 501.800 ;
        RECT 2576.990 501.740 2577.310 501.800 ;
        RECT 2018.090 501.600 2577.310 501.740 ;
        RECT 2018.090 501.540 2018.410 501.600 ;
        RECT 2576.990 501.540 2577.310 501.600 ;
      LAYER via ;
        RECT 2577.020 3194.680 2577.280 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
        RECT 2018.120 501.540 2018.380 501.800 ;
        RECT 2577.020 501.540 2577.280 501.800 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2577.020 3194.650 2577.280 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2018.250 510.340 2018.530 514.000 ;
        RECT 2018.180 510.000 2018.530 510.340 ;
        RECT 2018.180 501.830 2018.320 510.000 ;
        RECT 2577.080 501.830 2577.220 3194.650 ;
        RECT 2018.120 501.510 2018.380 501.830 ;
        RECT 2577.020 501.510 2577.280 501.830 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2611.490 3429.480 2611.810 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2611.490 3429.340 2901.150 3429.480 ;
        RECT 2611.490 3429.280 2611.810 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 2519.490 1876.700 2519.810 1876.760 ;
        RECT 2611.490 1876.700 2611.810 1876.760 ;
        RECT 2519.490 1876.560 2611.810 1876.700 ;
        RECT 2519.490 1876.500 2519.810 1876.560 ;
        RECT 2611.490 1876.500 2611.810 1876.560 ;
      LAYER via ;
        RECT 2611.520 3429.280 2611.780 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 2519.520 1876.500 2519.780 1876.760 ;
        RECT 2611.520 1876.500 2611.780 1876.760 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2611.520 3429.250 2611.780 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2611.580 1876.790 2611.720 3429.250 ;
        RECT 2519.520 1876.470 2519.780 1876.790 ;
        RECT 2611.520 1876.470 2611.780 1876.790 ;
        RECT 2519.580 1873.245 2519.720 1876.470 ;
        RECT 2519.510 1872.875 2519.790 1873.245 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2519.510 1872.920 2519.790 1873.200 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2506.000 1873.210 2510.000 1873.360 ;
        RECT 2519.485 1873.210 2519.815 1873.225 ;
        RECT 2506.000 1872.910 2519.815 1873.210 ;
        RECT 2506.000 1872.760 2510.000 1872.910 ;
        RECT 2519.485 1872.895 2519.815 1872.910 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2645.990 3501.560 2646.310 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 2645.990 3501.420 2717.610 3501.560 ;
        RECT 2645.990 3501.360 2646.310 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
        RECT 2519.490 2773.620 2519.810 2773.680 ;
        RECT 2645.990 2773.620 2646.310 2773.680 ;
        RECT 2519.490 2773.480 2646.310 2773.620 ;
        RECT 2519.490 2773.420 2519.810 2773.480 ;
        RECT 2645.990 2773.420 2646.310 2773.480 ;
      LAYER via ;
        RECT 2646.020 3501.360 2646.280 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
        RECT 2519.520 2773.420 2519.780 2773.680 ;
        RECT 2646.020 2773.420 2646.280 2773.680 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 2646.020 3501.330 2646.280 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 2646.080 2773.710 2646.220 3501.330 ;
        RECT 2519.520 2773.390 2519.780 2773.710 ;
        RECT 2646.020 2773.390 2646.280 2773.710 ;
        RECT 2519.580 2768.125 2519.720 2773.390 ;
        RECT 2519.510 2767.755 2519.790 2768.125 ;
      LAYER via2 ;
        RECT 2519.510 2767.800 2519.790 2768.080 ;
      LAYER met3 ;
        RECT 2506.000 2768.090 2510.000 2768.240 ;
        RECT 2519.485 2768.090 2519.815 2768.105 ;
        RECT 2506.000 2767.790 2519.815 2768.090 ;
        RECT 2506.000 2767.640 2510.000 2767.790 ;
        RECT 2519.485 2767.775 2519.815 2767.790 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.470 3464.160 2387.790 3464.220 ;
        RECT 2392.990 3464.160 2393.310 3464.220 ;
        RECT 2387.470 3464.020 2393.310 3464.160 ;
        RECT 2387.470 3463.960 2387.790 3464.020 ;
        RECT 2392.990 3463.960 2393.310 3464.020 ;
        RECT 2387.470 3367.600 2387.790 3367.660 ;
        RECT 2388.390 3367.600 2388.710 3367.660 ;
        RECT 2387.470 3367.460 2388.710 3367.600 ;
        RECT 2387.470 3367.400 2387.790 3367.460 ;
        RECT 2388.390 3367.400 2388.710 3367.460 ;
        RECT 2387.470 3270.700 2387.790 3270.760 ;
        RECT 2388.390 3270.700 2388.710 3270.760 ;
        RECT 2387.470 3270.560 2388.710 3270.700 ;
        RECT 2387.470 3270.500 2387.790 3270.560 ;
        RECT 2388.390 3270.500 2388.710 3270.560 ;
        RECT 2387.470 3174.140 2387.790 3174.200 ;
        RECT 2388.390 3174.140 2388.710 3174.200 ;
        RECT 2387.470 3174.000 2388.710 3174.140 ;
        RECT 2387.470 3173.940 2387.790 3174.000 ;
        RECT 2388.390 3173.940 2388.710 3174.000 ;
        RECT 399.350 3087.780 399.670 3087.840 ;
        RECT 2388.390 3087.780 2388.710 3087.840 ;
        RECT 399.350 3087.640 2388.710 3087.780 ;
        RECT 399.350 3087.580 399.670 3087.640 ;
        RECT 2388.390 3087.580 2388.710 3087.640 ;
      LAYER via ;
        RECT 2387.500 3463.960 2387.760 3464.220 ;
        RECT 2393.020 3463.960 2393.280 3464.220 ;
        RECT 2387.500 3367.400 2387.760 3367.660 ;
        RECT 2388.420 3367.400 2388.680 3367.660 ;
        RECT 2387.500 3270.500 2387.760 3270.760 ;
        RECT 2388.420 3270.500 2388.680 3270.760 ;
        RECT 2387.500 3173.940 2387.760 3174.200 ;
        RECT 2388.420 3173.940 2388.680 3174.200 ;
        RECT 399.380 3087.580 399.640 3087.840 ;
        RECT 2388.420 3087.580 2388.680 3087.840 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.620 3517.230 2393.220 3517.370 ;
        RECT 2393.080 3464.250 2393.220 3517.230 ;
        RECT 2387.500 3463.930 2387.760 3464.250 ;
        RECT 2393.020 3463.930 2393.280 3464.250 ;
        RECT 2387.560 3415.370 2387.700 3463.930 ;
        RECT 2387.560 3415.230 2388.620 3415.370 ;
        RECT 2388.480 3367.690 2388.620 3415.230 ;
        RECT 2387.500 3367.370 2387.760 3367.690 ;
        RECT 2388.420 3367.370 2388.680 3367.690 ;
        RECT 2387.560 3318.810 2387.700 3367.370 ;
        RECT 2387.560 3318.670 2388.620 3318.810 ;
        RECT 2388.480 3270.790 2388.620 3318.670 ;
        RECT 2387.500 3270.470 2387.760 3270.790 ;
        RECT 2388.420 3270.470 2388.680 3270.790 ;
        RECT 2387.560 3222.250 2387.700 3270.470 ;
        RECT 2387.560 3222.110 2388.620 3222.250 ;
        RECT 2388.480 3174.230 2388.620 3222.110 ;
        RECT 2387.500 3173.910 2387.760 3174.230 ;
        RECT 2388.420 3173.910 2388.680 3174.230 ;
        RECT 2387.560 3125.690 2387.700 3173.910 ;
        RECT 2387.560 3125.550 2388.620 3125.690 ;
        RECT 2388.480 3087.870 2388.620 3125.550 ;
        RECT 399.380 3087.550 399.640 3087.870 ;
        RECT 2388.420 3087.550 2388.680 3087.870 ;
        RECT 399.440 2651.165 399.580 3087.550 ;
        RECT 399.370 2650.795 399.650 2651.165 ;
      LAYER via2 ;
        RECT 399.370 2650.840 399.650 2651.120 ;
      LAYER met3 ;
        RECT 399.345 2651.130 399.675 2651.145 ;
        RECT 410.000 2651.130 414.000 2651.280 ;
        RECT 399.345 2650.830 414.000 2651.130 ;
        RECT 399.345 2650.815 399.675 2650.830 ;
        RECT 410.000 2650.680 414.000 2650.830 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 337.250 3501.900 337.570 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 337.250 3501.760 2068.550 3501.900 ;
        RECT 337.250 3501.700 337.570 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 337.280 3501.700 337.540 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 337.280 3501.670 337.540 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 337.340 502.365 337.480 3501.670 ;
        RECT 436.770 510.340 437.050 514.000 ;
        RECT 436.700 510.000 437.050 510.340 ;
        RECT 436.700 502.365 436.840 510.000 ;
        RECT 337.270 501.995 337.550 502.365 ;
        RECT 436.630 501.995 436.910 502.365 ;
      LAYER via2 ;
        RECT 337.270 502.040 337.550 502.320 ;
        RECT 436.630 502.040 436.910 502.320 ;
      LAYER met3 ;
        RECT 337.245 502.330 337.575 502.345 ;
        RECT 436.605 502.330 436.935 502.345 ;
        RECT 337.245 502.030 436.935 502.330 ;
        RECT 337.245 502.015 337.575 502.030 ;
        RECT 436.605 502.015 436.935 502.030 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 386.010 3502.240 386.330 3502.300 ;
        RECT 1743.930 3502.240 1744.250 3502.300 ;
        RECT 386.010 3502.100 1744.250 3502.240 ;
        RECT 386.010 3502.040 386.330 3502.100 ;
        RECT 1743.930 3502.040 1744.250 3502.100 ;
      LAYER via ;
        RECT 386.040 3502.040 386.300 3502.300 ;
        RECT 1743.960 3502.040 1744.220 3502.300 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.330 1744.160 3517.600 ;
        RECT 386.040 3502.010 386.300 3502.330 ;
        RECT 1743.960 3502.010 1744.220 3502.330 ;
        RECT 386.100 503.045 386.240 3502.010 ;
        RECT 622.610 510.340 622.890 514.000 ;
        RECT 622.540 510.000 622.890 510.340 ;
        RECT 622.540 503.045 622.680 510.000 ;
        RECT 386.030 502.675 386.310 503.045 ;
        RECT 622.470 502.675 622.750 503.045 ;
      LAYER via2 ;
        RECT 386.030 502.720 386.310 503.000 ;
        RECT 622.470 502.720 622.750 503.000 ;
      LAYER met3 ;
        RECT 386.005 503.010 386.335 503.025 ;
        RECT 622.445 503.010 622.775 503.025 ;
        RECT 386.005 502.710 622.775 503.010 ;
        RECT 386.005 502.695 386.335 502.710 ;
        RECT 622.445 502.695 622.775 502.710 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3502.580 1419.490 3502.640 ;
        RECT 1493.690 3502.580 1494.010 3502.640 ;
        RECT 1419.170 3502.440 1494.010 3502.580 ;
        RECT 1419.170 3502.380 1419.490 3502.440 ;
        RECT 1493.690 3502.380 1494.010 3502.440 ;
        RECT 1493.690 3039.500 1494.010 3039.560 ;
        RECT 1691.490 3039.500 1691.810 3039.560 ;
        RECT 1493.690 3039.360 1691.810 3039.500 ;
        RECT 1493.690 3039.300 1494.010 3039.360 ;
        RECT 1691.490 3039.300 1691.810 3039.360 ;
      LAYER via ;
        RECT 1419.200 3502.380 1419.460 3502.640 ;
        RECT 1493.720 3502.380 1493.980 3502.640 ;
        RECT 1493.720 3039.300 1493.980 3039.560 ;
        RECT 1691.520 3039.300 1691.780 3039.560 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3502.670 1419.400 3517.600 ;
        RECT 1419.200 3502.350 1419.460 3502.670 ;
        RECT 1493.720 3502.350 1493.980 3502.670 ;
        RECT 1493.780 3039.590 1493.920 3502.350 ;
        RECT 1493.720 3039.270 1493.980 3039.590 ;
        RECT 1691.520 3039.270 1691.780 3039.590 ;
        RECT 1691.580 3010.000 1691.720 3039.270 ;
        RECT 1691.580 3009.340 1691.930 3010.000 ;
        RECT 1691.650 3006.000 1691.930 3009.340 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1061.825 385.985 1062.455 386.155 ;
      LAYER mcon ;
        RECT 1062.285 385.985 1062.455 386.155 ;
      LAYER met1 ;
        RECT 362.550 1055.940 362.870 1056.000 ;
        RECT 393.370 1055.940 393.690 1056.000 ;
        RECT 362.550 1055.800 393.690 1055.940 ;
        RECT 362.550 1055.740 362.870 1055.800 ;
        RECT 393.370 1055.740 393.690 1055.800 ;
        RECT 362.550 386.140 362.870 386.200 ;
        RECT 1061.765 386.140 1062.055 386.185 ;
        RECT 362.550 386.000 1062.055 386.140 ;
        RECT 362.550 385.940 362.870 386.000 ;
        RECT 1061.765 385.955 1062.055 386.000 ;
        RECT 1062.225 386.140 1062.515 386.185 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 1062.225 386.000 2901.150 386.140 ;
        RECT 1062.225 385.955 1062.515 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 362.580 1055.740 362.840 1056.000 ;
        RECT 393.400 1055.740 393.660 1056.000 ;
        RECT 362.580 385.940 362.840 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 393.390 1060.955 393.670 1061.325 ;
        RECT 393.460 1056.030 393.600 1060.955 ;
        RECT 362.580 1055.710 362.840 1056.030 ;
        RECT 393.400 1055.710 393.660 1056.030 ;
        RECT 362.640 386.230 362.780 1055.710 ;
        RECT 362.580 385.910 362.840 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 393.390 1061.000 393.670 1061.280 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 393.365 1061.290 393.695 1061.305 ;
        RECT 410.000 1061.290 414.000 1061.440 ;
        RECT 393.365 1060.990 414.000 1061.290 ;
        RECT 393.365 1060.975 393.695 1060.990 ;
        RECT 410.000 1060.840 414.000 1060.990 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 425.185 500.565 425.355 502.775 ;
      LAYER mcon ;
        RECT 425.185 502.605 425.355 502.775 ;
      LAYER met1 ;
        RECT 406.710 3502.920 407.030 3502.980 ;
        RECT 1094.870 3502.920 1095.190 3502.980 ;
        RECT 406.710 3502.780 1095.190 3502.920 ;
        RECT 406.710 3502.720 407.030 3502.780 ;
        RECT 1094.870 3502.720 1095.190 3502.780 ;
        RECT 425.125 502.760 425.415 502.805 ;
        RECT 1647.330 502.760 1647.650 502.820 ;
        RECT 425.125 502.620 1647.650 502.760 ;
        RECT 425.125 502.575 425.415 502.620 ;
        RECT 1647.330 502.560 1647.650 502.620 ;
        RECT 406.710 500.720 407.030 500.780 ;
        RECT 425.125 500.720 425.415 500.765 ;
        RECT 406.710 500.580 425.415 500.720 ;
        RECT 406.710 500.520 407.030 500.580 ;
        RECT 425.125 500.535 425.415 500.580 ;
      LAYER via ;
        RECT 406.740 3502.720 407.000 3502.980 ;
        RECT 1094.900 3502.720 1095.160 3502.980 ;
        RECT 1647.360 502.560 1647.620 502.820 ;
        RECT 406.740 500.520 407.000 500.780 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3503.010 1095.100 3517.600 ;
        RECT 406.740 3502.690 407.000 3503.010 ;
        RECT 1094.900 3502.690 1095.160 3503.010 ;
        RECT 406.800 500.810 406.940 3502.690 ;
        RECT 1647.490 510.340 1647.770 514.000 ;
        RECT 1647.420 510.000 1647.770 510.340 ;
        RECT 1647.420 502.850 1647.560 510.000 ;
        RECT 1647.360 502.530 1647.620 502.850 ;
        RECT 406.740 500.490 407.000 500.810 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 351.510 3503.260 351.830 3503.320 ;
        RECT 770.570 3503.260 770.890 3503.320 ;
        RECT 351.510 3503.120 770.890 3503.260 ;
        RECT 351.510 3503.060 351.830 3503.120 ;
        RECT 770.570 3503.060 770.890 3503.120 ;
        RECT 351.510 501.400 351.830 501.460 ;
        RECT 659.250 501.400 659.570 501.460 ;
        RECT 351.510 501.260 659.570 501.400 ;
        RECT 351.510 501.200 351.830 501.260 ;
        RECT 659.250 501.200 659.570 501.260 ;
      LAYER via ;
        RECT 351.540 3503.060 351.800 3503.320 ;
        RECT 770.600 3503.060 770.860 3503.320 ;
        RECT 351.540 501.200 351.800 501.460 ;
        RECT 659.280 501.200 659.540 501.460 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.350 770.800 3517.600 ;
        RECT 351.540 3503.030 351.800 3503.350 ;
        RECT 770.600 3503.030 770.860 3503.350 ;
        RECT 351.600 501.490 351.740 3503.030 ;
        RECT 659.410 510.340 659.690 514.000 ;
        RECT 659.340 510.000 659.690 510.340 ;
        RECT 659.340 501.490 659.480 510.000 ;
        RECT 351.540 501.170 351.800 501.490 ;
        RECT 659.280 501.170 659.540 501.490 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 441.670 3498.500 441.990 3498.560 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 441.670 3498.360 446.130 3498.500 ;
        RECT 441.670 3498.300 441.990 3498.360 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 344.150 3012.300 344.470 3012.360 ;
        RECT 441.210 3012.300 441.530 3012.360 ;
        RECT 344.150 3012.160 441.530 3012.300 ;
        RECT 344.150 3012.100 344.470 3012.160 ;
        RECT 441.210 3012.100 441.530 3012.160 ;
        RECT 344.150 502.420 344.470 502.480 ;
        RECT 930.650 502.420 930.970 502.480 ;
        RECT 344.150 502.280 930.970 502.420 ;
        RECT 344.150 502.220 344.470 502.280 ;
        RECT 930.650 502.220 930.970 502.280 ;
      LAYER via ;
        RECT 441.700 3498.300 441.960 3498.560 ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 344.180 3012.100 344.440 3012.360 ;
        RECT 441.240 3012.100 441.500 3012.360 ;
        RECT 344.180 502.220 344.440 502.480 ;
        RECT 930.680 502.220 930.940 502.480 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 441.700 3498.270 441.960 3498.590 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 441.760 3016.210 441.900 3498.270 ;
        RECT 441.300 3016.070 441.900 3016.210 ;
        RECT 441.300 3012.390 441.440 3016.070 ;
        RECT 344.180 3012.070 344.440 3012.390 ;
        RECT 441.240 3012.070 441.500 3012.390 ;
        RECT 344.240 502.510 344.380 3012.070 ;
        RECT 930.810 510.340 931.090 514.000 ;
        RECT 930.740 510.000 931.090 510.340 ;
        RECT 930.740 502.510 930.880 510.000 ;
        RECT 344.180 502.190 344.440 502.510 ;
        RECT 930.680 502.190 930.940 502.510 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 441.670 504.460 441.990 504.520 ;
        RECT 2097.210 504.460 2097.530 504.520 ;
        RECT 441.670 504.320 2097.530 504.460 ;
        RECT 441.670 504.260 441.990 504.320 ;
        RECT 2097.210 504.260 2097.530 504.320 ;
        RECT 2097.210 501.400 2097.530 501.460 ;
        RECT 2203.930 501.400 2204.250 501.460 ;
        RECT 2097.210 501.260 2204.250 501.400 ;
        RECT 2097.210 501.200 2097.530 501.260 ;
        RECT 2203.930 501.200 2204.250 501.260 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 441.700 504.260 441.960 504.520 ;
        RECT 2097.240 504.260 2097.500 504.520 ;
        RECT 2097.240 501.200 2097.500 501.460 ;
        RECT 2203.960 501.200 2204.220 501.460 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 510.525 124.040 3498.270 ;
        RECT 123.830 510.155 124.110 510.525 ;
        RECT 441.690 510.155 441.970 510.525 ;
        RECT 2204.090 510.340 2204.370 514.000 ;
        RECT 441.760 504.550 441.900 510.155 ;
        RECT 2204.020 510.000 2204.370 510.340 ;
        RECT 441.700 504.230 441.960 504.550 ;
        RECT 2097.240 504.230 2097.500 504.550 ;
        RECT 2097.300 501.490 2097.440 504.230 ;
        RECT 2204.020 501.490 2204.160 510.000 ;
        RECT 2097.240 501.170 2097.500 501.490 ;
        RECT 2203.960 501.170 2204.220 501.490 ;
      LAYER via2 ;
        RECT 123.830 510.200 124.110 510.480 ;
        RECT 441.690 510.200 441.970 510.480 ;
      LAYER met3 ;
        RECT 123.805 510.490 124.135 510.505 ;
        RECT 441.665 510.490 441.995 510.505 ;
        RECT 123.805 510.190 441.995 510.490 ;
        RECT 123.805 510.175 124.135 510.190 ;
        RECT 441.665 510.175 441.995 510.190 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 2512.130 3339.720 2512.450 3339.780 ;
        RECT 17.090 3339.580 2512.450 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 2512.130 3339.520 2512.450 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 2512.160 3339.520 2512.420 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 2512.160 3339.490 2512.420 3339.810 ;
        RECT 2512.220 2074.525 2512.360 3339.490 ;
        RECT 2512.150 2074.155 2512.430 2074.525 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 2512.150 2074.200 2512.430 2074.480 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 2506.000 2074.490 2510.000 2074.640 ;
        RECT 2512.125 2074.490 2512.455 2074.505 ;
        RECT 2506.000 2074.190 2512.455 2074.490 ;
        RECT 2506.000 2074.040 2510.000 2074.190 ;
        RECT 2512.125 2074.175 2512.455 2074.190 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 244.790 3050.040 245.110 3050.100 ;
        RECT 17.090 3049.900 245.110 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 244.790 3049.840 245.110 3049.900 ;
        RECT 244.790 2359.840 245.110 2359.900 ;
        RECT 393.370 2359.840 393.690 2359.900 ;
        RECT 244.790 2359.700 393.690 2359.840 ;
        RECT 244.790 2359.640 245.110 2359.700 ;
        RECT 393.370 2359.640 393.690 2359.700 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 244.820 3049.840 245.080 3050.100 ;
        RECT 244.820 2359.640 245.080 2359.900 ;
        RECT 393.400 2359.640 393.660 2359.900 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 244.820 3049.810 245.080 3050.130 ;
        RECT 244.880 2359.930 245.020 3049.810 ;
        RECT 244.820 2359.610 245.080 2359.930 ;
        RECT 393.400 2359.610 393.660 2359.930 ;
        RECT 393.460 2358.765 393.600 2359.610 ;
        RECT 393.390 2358.395 393.670 2358.765 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 393.390 2358.440 393.670 2358.720 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 393.365 2358.730 393.695 2358.745 ;
        RECT 410.000 2358.730 414.000 2358.880 ;
        RECT 393.365 2358.430 414.000 2358.730 ;
        RECT 393.365 2358.415 393.695 2358.430 ;
        RECT 410.000 2358.280 414.000 2358.430 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 196.490 2760.360 196.810 2760.420 ;
        RECT 15.710 2760.220 196.810 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 196.490 2760.160 196.810 2760.220 ;
        RECT 196.490 504.120 196.810 504.180 ;
        RECT 832.210 504.120 832.530 504.180 ;
        RECT 196.490 503.980 832.530 504.120 ;
        RECT 196.490 503.920 196.810 503.980 ;
        RECT 832.210 503.920 832.530 503.980 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 196.520 2760.160 196.780 2760.420 ;
        RECT 196.520 503.920 196.780 504.180 ;
        RECT 832.240 503.920 832.500 504.180 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 196.520 2760.130 196.780 2760.450 ;
        RECT 196.580 504.210 196.720 2760.130 ;
        RECT 832.370 510.340 832.650 514.000 ;
        RECT 832.300 510.000 832.650 510.340 ;
        RECT 832.300 504.210 832.440 510.000 ;
        RECT 196.520 503.890 196.780 504.210 ;
        RECT 832.240 503.890 832.500 504.210 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 936.705 3002.285 936.875 3006.535 ;
        RECT 396.205 2483.785 396.375 2508.775 ;
      LAYER mcon ;
        RECT 936.705 3006.365 936.875 3006.535 ;
        RECT 396.205 2508.605 396.375 2508.775 ;
      LAYER met1 ;
        RECT 936.630 3006.520 936.950 3006.580 ;
        RECT 936.435 3006.380 936.950 3006.520 ;
        RECT 936.630 3006.320 936.950 3006.380 ;
        RECT 418.210 3002.440 418.530 3002.500 ;
        RECT 936.645 3002.440 936.935 3002.485 ;
        RECT 418.210 3002.300 936.935 3002.440 ;
        RECT 418.210 3002.240 418.530 3002.300 ;
        RECT 936.645 3002.255 936.935 3002.300 ;
        RECT 396.145 2508.760 396.435 2508.805 ;
        RECT 414.530 2508.760 414.850 2508.820 ;
        RECT 396.145 2508.620 414.850 2508.760 ;
        RECT 396.145 2508.575 396.435 2508.620 ;
        RECT 414.530 2508.560 414.850 2508.620 ;
        RECT 17.090 2483.940 17.410 2484.000 ;
        RECT 396.145 2483.940 396.435 2483.985 ;
        RECT 17.090 2483.800 396.435 2483.940 ;
        RECT 17.090 2483.740 17.410 2483.800 ;
        RECT 396.145 2483.755 396.435 2483.800 ;
      LAYER via ;
        RECT 936.660 3006.320 936.920 3006.580 ;
        RECT 418.240 3002.240 418.500 3002.500 ;
        RECT 414.560 2508.560 414.820 2508.820 ;
        RECT 17.120 2483.740 17.380 2484.000 ;
      LAYER met2 ;
        RECT 938.170 3006.690 938.450 3010.000 ;
        RECT 936.720 3006.610 938.450 3006.690 ;
        RECT 936.660 3006.550 938.450 3006.610 ;
        RECT 936.660 3006.290 936.920 3006.550 ;
        RECT 938.170 3006.000 938.450 3006.550 ;
        RECT 418.240 3002.210 418.500 3002.530 ;
        RECT 418.300 2509.610 418.440 3002.210 ;
        RECT 414.620 2509.470 418.440 2509.610 ;
        RECT 414.620 2508.850 414.760 2509.470 ;
        RECT 414.560 2508.530 414.820 2508.850 ;
        RECT 17.120 2483.710 17.380 2484.030 ;
        RECT 17.180 2477.765 17.320 2483.710 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
      LAYER via2 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2087.160 17.410 2087.220 ;
        RECT 348.750 2087.160 349.070 2087.220 ;
        RECT 17.090 2087.020 349.070 2087.160 ;
        RECT 17.090 2086.960 17.410 2087.020 ;
        RECT 348.750 2086.960 349.070 2087.020 ;
        RECT 348.750 502.080 349.070 502.140 ;
        RECT 881.890 502.080 882.210 502.140 ;
        RECT 348.750 501.940 882.210 502.080 ;
        RECT 348.750 501.880 349.070 501.940 ;
        RECT 881.890 501.880 882.210 501.940 ;
      LAYER via ;
        RECT 17.120 2086.960 17.380 2087.220 ;
        RECT 348.780 2086.960 349.040 2087.220 ;
        RECT 348.780 501.880 349.040 502.140 ;
        RECT 881.920 501.880 882.180 502.140 ;
      LAYER met2 ;
        RECT 17.110 2189.755 17.390 2190.125 ;
        RECT 17.180 2087.250 17.320 2189.755 ;
        RECT 17.120 2086.930 17.380 2087.250 ;
        RECT 348.780 2086.930 349.040 2087.250 ;
        RECT 348.840 502.170 348.980 2086.930 ;
        RECT 882.050 510.340 882.330 514.000 ;
        RECT 881.980 510.000 882.330 510.340 ;
        RECT 881.980 502.170 882.120 510.000 ;
        RECT 348.780 501.850 349.040 502.170 ;
        RECT 881.920 501.850 882.180 502.170 ;
      LAYER via2 ;
        RECT 17.110 2189.800 17.390 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.085 2190.090 17.415 2190.105 ;
        RECT -4.800 2189.790 17.415 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.085 2189.775 17.415 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1897.780 17.410 1897.840 ;
        RECT 65.850 1897.780 66.170 1897.840 ;
        RECT 17.090 1897.640 66.170 1897.780 ;
        RECT 17.090 1897.580 17.410 1897.640 ;
        RECT 65.850 1897.580 66.170 1897.640 ;
        RECT 65.850 1759.400 66.170 1759.460 ;
        RECT 393.370 1759.400 393.690 1759.460 ;
        RECT 65.850 1759.260 393.690 1759.400 ;
        RECT 65.850 1759.200 66.170 1759.260 ;
        RECT 393.370 1759.200 393.690 1759.260 ;
      LAYER via ;
        RECT 17.120 1897.580 17.380 1897.840 ;
        RECT 65.880 1897.580 66.140 1897.840 ;
        RECT 65.880 1759.200 66.140 1759.460 ;
        RECT 393.400 1759.200 393.660 1759.460 ;
      LAYER met2 ;
        RECT 17.110 1902.795 17.390 1903.165 ;
        RECT 17.180 1897.870 17.320 1902.795 ;
        RECT 17.120 1897.550 17.380 1897.870 ;
        RECT 65.880 1897.550 66.140 1897.870 ;
        RECT 65.940 1759.490 66.080 1897.550 ;
        RECT 65.880 1759.170 66.140 1759.490 ;
        RECT 393.400 1759.170 393.660 1759.490 ;
        RECT 393.460 1756.285 393.600 1759.170 ;
        RECT 393.390 1755.915 393.670 1756.285 ;
      LAYER via2 ;
        RECT 17.110 1902.840 17.390 1903.120 ;
        RECT 393.390 1755.960 393.670 1756.240 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.085 1903.130 17.415 1903.145 ;
        RECT -4.800 1902.830 17.415 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.085 1902.815 17.415 1902.830 ;
        RECT 393.365 1756.250 393.695 1756.265 ;
        RECT 410.000 1756.250 414.000 1756.400 ;
        RECT 393.365 1755.950 414.000 1756.250 ;
        RECT 393.365 1755.935 393.695 1755.950 ;
        RECT 410.000 1755.800 414.000 1755.950 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2856.920 2519.810 2856.980 ;
        RECT 2694.290 2856.920 2694.610 2856.980 ;
        RECT 2519.490 2856.780 2694.610 2856.920 ;
        RECT 2519.490 2856.720 2519.810 2856.780 ;
        RECT 2694.290 2856.720 2694.610 2856.780 ;
        RECT 2694.290 620.740 2694.610 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2694.290 620.600 2901.150 620.740 ;
        RECT 2694.290 620.540 2694.610 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2519.520 2856.720 2519.780 2856.980 ;
        RECT 2694.320 2856.720 2694.580 2856.980 ;
        RECT 2694.320 620.540 2694.580 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2519.510 2858.875 2519.790 2859.245 ;
        RECT 2519.580 2857.010 2519.720 2858.875 ;
        RECT 2519.520 2856.690 2519.780 2857.010 ;
        RECT 2694.320 2856.690 2694.580 2857.010 ;
        RECT 2694.380 620.830 2694.520 2856.690 ;
        RECT 2694.320 620.510 2694.580 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2519.510 2858.920 2519.790 2859.200 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2506.000 2859.210 2510.000 2859.360 ;
        RECT 2519.485 2859.210 2519.815 2859.225 ;
        RECT 2506.000 2858.910 2519.815 2859.210 ;
        RECT 2506.000 2858.760 2510.000 2858.910 ;
        RECT 2519.485 2858.895 2519.815 2858.910 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1357.145 3003.305 1357.315 3006.535 ;
      LAYER mcon ;
        RECT 1357.145 3006.365 1357.315 3006.535 ;
      LAYER met1 ;
        RECT 1357.070 3006.520 1357.390 3006.580 ;
        RECT 1356.875 3006.380 1357.390 3006.520 ;
        RECT 1357.070 3006.320 1357.390 3006.380 ;
        RECT 382.790 3003.460 383.110 3003.520 ;
        RECT 1357.085 3003.460 1357.375 3003.505 ;
        RECT 382.790 3003.320 1357.375 3003.460 ;
        RECT 382.790 3003.260 383.110 3003.320 ;
        RECT 1357.085 3003.275 1357.375 3003.320 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 382.790 1621.360 383.110 1621.420 ;
        RECT 16.170 1621.220 383.110 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 382.790 1621.160 383.110 1621.220 ;
      LAYER via ;
        RECT 1357.100 3006.320 1357.360 3006.580 ;
        RECT 382.820 3003.260 383.080 3003.520 ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 382.820 1621.160 383.080 1621.420 ;
      LAYER met2 ;
        RECT 1358.610 3006.690 1358.890 3010.000 ;
        RECT 1357.160 3006.610 1358.890 3006.690 ;
        RECT 1357.100 3006.550 1358.890 3006.610 ;
        RECT 1357.100 3006.290 1357.360 3006.550 ;
        RECT 1358.610 3006.000 1358.890 3006.550 ;
        RECT 382.820 3003.230 383.080 3003.550 ;
        RECT 382.880 1621.450 383.020 3003.230 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 382.820 1621.130 383.080 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 17.180 1394.525 17.320 1400.275 ;
        RECT 17.110 1394.155 17.390 1394.525 ;
      LAYER via2 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
        RECT 17.110 1394.200 17.390 1394.480 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
        RECT 17.085 1394.490 17.415 1394.505 ;
        RECT 106.070 1394.490 106.450 1394.500 ;
        RECT 17.085 1394.190 106.450 1394.490 ;
        RECT 17.085 1394.175 17.415 1394.190 ;
        RECT 106.070 1394.180 106.450 1394.190 ;
        RECT 2506.000 1032.280 2510.000 1032.880 ;
        RECT 2507.310 1028.660 2507.610 1032.280 ;
        RECT 306.630 1028.650 307.010 1028.660 ;
        RECT 379.310 1028.650 379.690 1028.660 ;
        RECT 306.630 1028.350 379.690 1028.650 ;
        RECT 306.630 1028.340 307.010 1028.350 ;
        RECT 379.310 1028.340 379.690 1028.350 ;
        RECT 2507.270 1028.340 2507.650 1028.660 ;
        RECT 379.310 1025.250 379.690 1025.260 ;
        RECT 394.950 1025.250 395.330 1025.260 ;
        RECT 379.310 1024.950 395.330 1025.250 ;
        RECT 379.310 1024.940 379.690 1024.950 ;
        RECT 394.950 1024.940 395.330 1024.950 ;
      LAYER via3 ;
        RECT 106.100 1394.180 106.420 1394.500 ;
        RECT 306.660 1028.340 306.980 1028.660 ;
        RECT 379.340 1028.340 379.660 1028.660 ;
        RECT 2507.300 1028.340 2507.620 1028.660 ;
        RECT 379.340 1024.940 379.660 1025.260 ;
        RECT 394.980 1024.940 395.300 1025.260 ;
      LAYER met4 ;
        RECT 106.095 1394.175 106.425 1394.505 ;
        RECT 106.110 1032.490 106.410 1394.175 ;
        RECT 2433.270 1041.510 2434.450 1042.690 ;
        RECT 2460.870 1041.510 2462.050 1042.690 ;
        RECT 2433.710 1032.490 2434.010 1041.510 ;
        RECT 105.670 1031.310 106.850 1032.490 ;
        RECT 306.230 1031.310 307.410 1032.490 ;
        RECT 2433.270 1031.310 2434.450 1032.490 ;
        RECT 306.670 1028.665 306.970 1031.310 ;
        RECT 2461.310 1029.090 2461.610 1041.510 ;
        RECT 306.655 1028.335 306.985 1028.665 ;
        RECT 379.335 1028.335 379.665 1028.665 ;
        RECT 379.350 1025.265 379.650 1028.335 ;
        RECT 2460.870 1027.910 2462.050 1029.090 ;
        RECT 2505.030 1028.650 2506.210 1029.090 ;
        RECT 2507.295 1028.650 2507.625 1028.665 ;
        RECT 2505.030 1028.350 2507.625 1028.650 ;
        RECT 2505.030 1027.910 2506.210 1028.350 ;
        RECT 2507.295 1028.335 2507.625 1028.350 ;
        RECT 379.335 1024.935 379.665 1025.265 ;
        RECT 394.550 1024.510 395.730 1025.690 ;
      LAYER met5 ;
        RECT 2433.060 1041.300 2462.260 1042.900 ;
        RECT -179.395 1031.100 131.900 1032.700 ;
        RECT 130.300 1025.900 131.900 1031.100 ;
        RECT 253.580 1031.100 307.620 1032.700 ;
        RECT 457.820 1031.100 470.460 1032.700 ;
        RECT 253.580 1025.900 255.180 1031.100 ;
        RECT 457.820 1025.900 459.420 1031.100 ;
        RECT 130.300 1024.300 255.180 1025.900 ;
        RECT 394.340 1024.300 459.420 1025.900 ;
        RECT 468.860 1025.900 470.460 1031.100 ;
        RECT 473.460 1031.100 518.300 1032.700 ;
        RECT 473.460 1025.900 475.060 1031.100 ;
        RECT 468.860 1024.300 475.060 1025.900 ;
        RECT 516.700 1025.900 518.300 1031.100 ;
        RECT 564.540 1031.100 614.900 1032.700 ;
        RECT 564.540 1025.900 566.140 1031.100 ;
        RECT 516.700 1024.300 566.140 1025.900 ;
        RECT 613.300 1025.900 614.900 1031.100 ;
        RECT 661.140 1031.100 711.500 1032.700 ;
        RECT 661.140 1025.900 662.740 1031.100 ;
        RECT 613.300 1024.300 662.740 1025.900 ;
        RECT 709.900 1025.900 711.500 1031.100 ;
        RECT 757.740 1031.100 808.100 1032.700 ;
        RECT 757.740 1025.900 759.340 1031.100 ;
        RECT 709.900 1024.300 759.340 1025.900 ;
        RECT 806.500 1025.900 808.100 1031.100 ;
        RECT 854.340 1031.100 904.700 1032.700 ;
        RECT 854.340 1025.900 855.940 1031.100 ;
        RECT 806.500 1024.300 855.940 1025.900 ;
        RECT 903.100 1025.900 904.700 1031.100 ;
        RECT 950.940 1031.100 1001.300 1032.700 ;
        RECT 950.940 1025.900 952.540 1031.100 ;
        RECT 903.100 1024.300 952.540 1025.900 ;
        RECT 999.700 1025.900 1001.300 1031.100 ;
        RECT 1047.540 1031.100 1097.900 1032.700 ;
        RECT 1047.540 1025.900 1049.140 1031.100 ;
        RECT 999.700 1024.300 1049.140 1025.900 ;
        RECT 1096.300 1025.900 1097.900 1031.100 ;
        RECT 1144.140 1031.100 1194.500 1032.700 ;
        RECT 1144.140 1025.900 1145.740 1031.100 ;
        RECT 1096.300 1024.300 1145.740 1025.900 ;
        RECT 1192.900 1025.900 1194.500 1031.100 ;
        RECT 1240.740 1031.100 1291.100 1032.700 ;
        RECT 1240.740 1025.900 1242.340 1031.100 ;
        RECT 1192.900 1024.300 1242.340 1025.900 ;
        RECT 1289.500 1025.900 1291.100 1031.100 ;
        RECT 1337.340 1031.100 1387.700 1032.700 ;
        RECT 1337.340 1025.900 1338.940 1031.100 ;
        RECT 1289.500 1024.300 1338.940 1025.900 ;
        RECT 1386.100 1025.900 1387.700 1031.100 ;
        RECT 1433.940 1031.100 1484.300 1032.700 ;
        RECT 1433.940 1025.900 1435.540 1031.100 ;
        RECT 1386.100 1024.300 1435.540 1025.900 ;
        RECT 1482.700 1025.900 1484.300 1031.100 ;
        RECT 1530.540 1031.100 1580.900 1032.700 ;
        RECT 1530.540 1025.900 1532.140 1031.100 ;
        RECT 1482.700 1024.300 1532.140 1025.900 ;
        RECT 1579.300 1025.900 1580.900 1031.100 ;
        RECT 1627.140 1031.100 1677.500 1032.700 ;
        RECT 1627.140 1025.900 1628.740 1031.100 ;
        RECT 1579.300 1024.300 1628.740 1025.900 ;
        RECT 1675.900 1025.900 1677.500 1031.100 ;
        RECT 1723.740 1031.100 1774.100 1032.700 ;
        RECT 1723.740 1025.900 1725.340 1031.100 ;
        RECT 1675.900 1024.300 1725.340 1025.900 ;
        RECT 1772.500 1025.900 1774.100 1031.100 ;
        RECT 1820.340 1031.100 1870.700 1032.700 ;
        RECT 1820.340 1025.900 1821.940 1031.100 ;
        RECT 1772.500 1024.300 1821.940 1025.900 ;
        RECT 1869.100 1025.900 1870.700 1031.100 ;
        RECT 1916.940 1031.100 1967.300 1032.700 ;
        RECT 1916.940 1025.900 1918.540 1031.100 ;
        RECT 1869.100 1024.300 1918.540 1025.900 ;
        RECT 1965.700 1025.900 1967.300 1031.100 ;
        RECT 2013.540 1031.100 2063.900 1032.700 ;
        RECT 2013.540 1025.900 2015.140 1031.100 ;
        RECT 1965.700 1024.300 2015.140 1025.900 ;
        RECT 2062.300 1025.900 2063.900 1031.100 ;
        RECT 2110.140 1031.100 2160.500 1032.700 ;
        RECT 2110.140 1025.900 2111.740 1031.100 ;
        RECT 2062.300 1024.300 2111.740 1025.900 ;
        RECT 2158.900 1025.900 2160.500 1031.100 ;
        RECT 2206.740 1031.100 2257.100 1032.700 ;
        RECT 2206.740 1025.900 2208.340 1031.100 ;
        RECT 2158.900 1024.300 2208.340 1025.900 ;
        RECT 2255.500 1025.900 2257.100 1031.100 ;
        RECT 2303.340 1031.100 2353.700 1032.700 ;
        RECT 2303.340 1025.900 2304.940 1031.100 ;
        RECT 2255.500 1024.300 2304.940 1025.900 ;
        RECT 2352.100 1025.900 2353.700 1031.100 ;
        RECT 2415.580 1031.100 2434.660 1032.700 ;
        RECT 2415.580 1025.900 2417.180 1031.100 ;
        RECT 2460.660 1027.700 2506.420 1029.300 ;
        RECT 2352.100 1024.300 2417.180 1025.900 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1739.865 3002.965 1740.035 3006.535 ;
      LAYER mcon ;
        RECT 1739.865 3006.365 1740.035 3006.535 ;
      LAYER met1 ;
        RECT 1739.790 3006.520 1740.110 3006.580 ;
        RECT 1739.595 3006.380 1740.110 3006.520 ;
        RECT 1739.790 3006.320 1740.110 3006.380 ;
        RECT 348.290 3003.120 348.610 3003.180 ;
        RECT 1739.805 3003.120 1740.095 3003.165 ;
        RECT 348.290 3002.980 1740.095 3003.120 ;
        RECT 348.290 3002.920 348.610 3002.980 ;
        RECT 1739.805 3002.935 1740.095 3002.980 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 348.290 1186.840 348.610 1186.900 ;
        RECT 17.090 1186.700 348.610 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 348.290 1186.640 348.610 1186.700 ;
      LAYER via ;
        RECT 1739.820 3006.320 1740.080 3006.580 ;
        RECT 348.320 3002.920 348.580 3003.180 ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 348.320 1186.640 348.580 1186.900 ;
      LAYER met2 ;
        RECT 1741.330 3006.690 1741.610 3010.000 ;
        RECT 1739.880 3006.610 1741.610 3006.690 ;
        RECT 1739.820 3006.550 1741.610 3006.610 ;
        RECT 1739.820 3006.290 1740.080 3006.550 ;
        RECT 1741.330 3006.000 1741.610 3006.550 ;
        RECT 348.320 3002.890 348.580 3003.210 ;
        RECT 348.380 1186.930 348.520 3002.890 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 348.320 1186.610 348.580 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1271.050 3006.320 1271.370 3006.580 ;
        RECT 355.650 3004.140 355.970 3004.200 ;
        RECT 1271.140 3004.140 1271.280 3006.320 ;
        RECT 355.650 3004.000 1271.280 3004.140 ;
        RECT 355.650 3003.940 355.970 3004.000 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 355.650 972.640 355.970 972.700 ;
        RECT 15.710 972.500 355.970 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 355.650 972.440 355.970 972.500 ;
      LAYER via ;
        RECT 1271.080 3006.320 1271.340 3006.580 ;
        RECT 355.680 3003.940 355.940 3004.200 ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 355.680 972.440 355.940 972.700 ;
      LAYER met2 ;
        RECT 1272.130 3006.690 1272.410 3010.000 ;
        RECT 1271.140 3006.610 1272.410 3006.690 ;
        RECT 1271.080 3006.550 1272.410 3006.610 ;
        RECT 1271.080 3006.290 1271.340 3006.550 ;
        RECT 1272.130 3006.000 1272.410 3006.550 ;
        RECT 355.680 3003.910 355.940 3004.230 ;
        RECT 355.740 972.730 355.880 3003.910 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 355.680 972.410 355.940 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 3022.840 341.710 3022.900 ;
        RECT 765.050 3022.840 765.370 3022.900 ;
        RECT 341.390 3022.700 765.370 3022.840 ;
        RECT 341.390 3022.640 341.710 3022.700 ;
        RECT 765.050 3022.640 765.370 3022.700 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 341.390 758.780 341.710 758.840 ;
        RECT 15.710 758.640 341.710 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 341.390 758.580 341.710 758.640 ;
      LAYER via ;
        RECT 341.420 3022.640 341.680 3022.900 ;
        RECT 765.080 3022.640 765.340 3022.900 ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 341.420 758.580 341.680 758.840 ;
      LAYER met2 ;
        RECT 341.420 3022.610 341.680 3022.930 ;
        RECT 765.080 3022.610 765.340 3022.930 ;
        RECT 341.480 758.870 341.620 3022.610 ;
        RECT 765.140 3010.000 765.280 3022.610 ;
        RECT 765.140 3009.340 765.490 3010.000 ;
        RECT 765.210 3006.000 765.490 3009.340 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 341.420 758.550 341.680 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1138.900 2520.730 1138.960 ;
        RECT 2554.450 1138.900 2554.770 1138.960 ;
        RECT 2520.410 1138.760 2554.770 1138.900 ;
        RECT 2520.410 1138.700 2520.730 1138.760 ;
        RECT 2554.450 1138.700 2554.770 1138.760 ;
        RECT 20.310 538.460 20.630 538.520 ;
        RECT 371.290 538.460 371.610 538.520 ;
        RECT 20.310 538.320 371.610 538.460 ;
        RECT 20.310 538.260 20.630 538.320 ;
        RECT 371.290 538.260 371.610 538.320 ;
        RECT 371.290 510.580 371.610 510.640 ;
        RECT 2554.450 510.580 2554.770 510.640 ;
        RECT 371.290 510.440 2554.770 510.580 ;
        RECT 371.290 510.380 371.610 510.440 ;
        RECT 2554.450 510.380 2554.770 510.440 ;
      LAYER via ;
        RECT 2520.440 1138.700 2520.700 1138.960 ;
        RECT 2554.480 1138.700 2554.740 1138.960 ;
        RECT 20.340 538.260 20.600 538.520 ;
        RECT 371.320 538.260 371.580 538.520 ;
        RECT 371.320 510.380 371.580 510.640 ;
        RECT 2554.480 510.380 2554.740 510.640 ;
      LAYER met2 ;
        RECT 2520.430 1142.555 2520.710 1142.925 ;
        RECT 2520.500 1138.990 2520.640 1142.555 ;
        RECT 2520.440 1138.670 2520.700 1138.990 ;
        RECT 2554.480 1138.670 2554.740 1138.990 ;
        RECT 20.340 538.405 20.600 538.550 ;
        RECT 20.330 538.035 20.610 538.405 ;
        RECT 371.320 538.230 371.580 538.550 ;
        RECT 371.380 510.670 371.520 538.230 ;
        RECT 2554.540 510.670 2554.680 1138.670 ;
        RECT 371.320 510.350 371.580 510.670 ;
        RECT 2554.480 510.350 2554.740 510.670 ;
      LAYER via2 ;
        RECT 2520.430 1142.600 2520.710 1142.880 ;
        RECT 20.330 538.080 20.610 538.360 ;
      LAYER met3 ;
        RECT 2506.000 1142.890 2510.000 1143.040 ;
        RECT 2520.405 1142.890 2520.735 1142.905 ;
        RECT 2506.000 1142.590 2520.735 1142.890 ;
        RECT 2506.000 1142.440 2510.000 1142.590 ;
        RECT 2520.405 1142.575 2520.735 1142.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 20.305 538.370 20.635 538.385 ;
        RECT -4.800 538.070 20.635 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 20.305 538.055 20.635 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 168.890 1987.540 169.210 1987.600 ;
        RECT 393.370 1987.540 393.690 1987.600 ;
        RECT 168.890 1987.400 393.690 1987.540 ;
        RECT 168.890 1987.340 169.210 1987.400 ;
        RECT 393.370 1987.340 393.690 1987.400 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 168.890 324.260 169.210 324.320 ;
        RECT 16.630 324.120 169.210 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 168.890 324.060 169.210 324.120 ;
      LAYER via ;
        RECT 168.920 1987.340 169.180 1987.600 ;
        RECT 393.400 1987.340 393.660 1987.600 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 168.920 324.060 169.180 324.320 ;
      LAYER met2 ;
        RECT 393.390 1992.555 393.670 1992.925 ;
        RECT 393.460 1987.630 393.600 1992.555 ;
        RECT 168.920 1987.310 169.180 1987.630 ;
        RECT 393.400 1987.310 393.660 1987.630 ;
        RECT 168.980 324.350 169.120 1987.310 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 168.920 324.030 169.180 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 393.390 1992.600 393.670 1992.880 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 393.365 1992.890 393.695 1992.905 ;
        RECT 410.000 1992.890 414.000 1993.040 ;
        RECT 393.365 1992.590 414.000 1992.890 ;
        RECT 393.365 1992.575 393.695 1992.590 ;
        RECT 410.000 1992.440 414.000 1992.590 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2822.240 2519.810 2822.300 ;
        RECT 2574.230 2822.240 2574.550 2822.300 ;
        RECT 2519.490 2822.100 2574.550 2822.240 ;
        RECT 2519.490 2822.040 2519.810 2822.100 ;
        RECT 2574.230 2822.040 2574.550 2822.100 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 2574.230 110.400 2574.550 110.460 ;
        RECT 15.710 110.260 2574.550 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 2574.230 110.200 2574.550 110.260 ;
      LAYER via ;
        RECT 2519.520 2822.040 2519.780 2822.300 ;
        RECT 2574.260 2822.040 2574.520 2822.300 ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 2574.260 110.200 2574.520 110.460 ;
      LAYER met2 ;
        RECT 2519.510 2822.155 2519.790 2822.525 ;
        RECT 2519.520 2822.010 2519.780 2822.155 ;
        RECT 2574.260 2822.010 2574.520 2822.330 ;
        RECT 2574.320 110.490 2574.460 2822.010 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 2574.260 110.170 2574.520 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 2519.510 2822.200 2519.790 2822.480 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 2506.000 2822.490 2510.000 2822.640 ;
        RECT 2519.485 2822.490 2519.815 2822.505 ;
        RECT 2506.000 2822.190 2519.815 2822.490 ;
        RECT 2506.000 2822.040 2510.000 2822.190 ;
        RECT 2519.485 2822.175 2519.815 2822.190 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.350 3006.320 1779.670 3006.580 ;
        RECT 1779.440 3003.800 1779.580 3006.320 ;
        RECT 2556.750 3003.800 2557.070 3003.860 ;
        RECT 1779.440 3003.660 2557.070 3003.800 ;
        RECT 2556.750 3003.600 2557.070 3003.660 ;
        RECT 2556.750 855.340 2557.070 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2556.750 855.200 2901.150 855.340 ;
        RECT 2556.750 855.140 2557.070 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 1779.380 3006.320 1779.640 3006.580 ;
        RECT 2556.780 3003.600 2557.040 3003.860 ;
        RECT 2556.780 855.140 2557.040 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 1778.130 3006.690 1778.410 3010.000 ;
        RECT 1778.130 3006.610 1779.580 3006.690 ;
        RECT 1778.130 3006.550 1779.640 3006.610 ;
        RECT 1778.130 3006.000 1778.410 3006.550 ;
        RECT 1779.380 3006.290 1779.640 3006.550 ;
        RECT 2556.780 3003.570 2557.040 3003.890 ;
        RECT 2556.840 855.430 2556.980 3003.570 ;
        RECT 2556.780 855.110 2557.040 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1428.580 2520.730 1428.640 ;
        RECT 2701.190 1428.580 2701.510 1428.640 ;
        RECT 2520.410 1428.440 2701.510 1428.580 ;
        RECT 2520.410 1428.380 2520.730 1428.440 ;
        RECT 2701.190 1428.380 2701.510 1428.440 ;
        RECT 2701.190 1089.940 2701.510 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2701.190 1089.800 2901.150 1089.940 ;
        RECT 2701.190 1089.740 2701.510 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2520.440 1428.380 2520.700 1428.640 ;
        RECT 2701.220 1428.380 2701.480 1428.640 ;
        RECT 2701.220 1089.740 2701.480 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2520.430 1434.955 2520.710 1435.325 ;
        RECT 2520.500 1428.670 2520.640 1434.955 ;
        RECT 2520.440 1428.350 2520.700 1428.670 ;
        RECT 2701.220 1428.350 2701.480 1428.670 ;
        RECT 2701.280 1090.030 2701.420 1428.350 ;
        RECT 2701.220 1089.710 2701.480 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2520.430 1435.000 2520.710 1435.280 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2506.000 1435.290 2510.000 1435.440 ;
        RECT 2520.405 1435.290 2520.735 1435.305 ;
        RECT 2506.000 1434.990 2520.735 1435.290 ;
        RECT 2506.000 1434.840 2510.000 1434.990 ;
        RECT 2520.405 1434.975 2520.735 1434.990 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 412.430 1885.140 412.810 1885.460 ;
        RECT 412.470 1884.240 412.770 1885.140 ;
        RECT 410.000 1883.640 414.000 1884.240 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2691.310 1319.390 2739.450 1319.690 ;
        RECT 2645.270 1318.330 2645.650 1318.340 ;
        RECT 2691.310 1318.330 2691.610 1319.390 ;
        RECT 2739.150 1319.010 2739.450 1319.390 ;
        RECT 2787.910 1319.390 2836.050 1319.690 ;
        RECT 2739.150 1318.710 2787.290 1319.010 ;
        RECT 2645.270 1318.030 2691.610 1318.330 ;
        RECT 2786.990 1318.330 2787.290 1318.710 ;
        RECT 2787.910 1318.330 2788.210 1319.390 ;
        RECT 2835.750 1319.010 2836.050 1319.390 ;
        RECT 2916.710 1319.390 2924.800 1319.690 ;
        RECT 2835.750 1318.710 2883.890 1319.010 ;
        RECT 2786.990 1318.030 2788.210 1318.330 ;
        RECT 2883.590 1318.330 2883.890 1318.710 ;
        RECT 2916.710 1318.330 2917.010 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 2883.590 1318.030 2917.010 1318.330 ;
        RECT 2645.270 1318.020 2645.650 1318.030 ;
      LAYER via3 ;
        RECT 412.460 1885.140 412.780 1885.460 ;
        RECT 2645.300 1318.020 2645.620 1318.340 ;
      LAYER met4 ;
        RECT 2644.870 1888.110 2646.050 1889.290 ;
        RECT 412.030 1884.710 413.210 1885.890 ;
        RECT 2645.310 1318.345 2645.610 1888.110 ;
        RECT 2645.295 1318.015 2645.625 1318.345 ;
      LAYER met5 ;
        RECT 2552.660 1891.300 2601.180 1892.900 ;
        RECT 882.860 1887.900 931.380 1889.500 ;
        RECT 411.820 1884.500 448.380 1886.100 ;
        RECT 446.780 1882.700 448.380 1884.500 ;
        RECT 446.780 1881.100 484.260 1882.700 ;
        RECT 482.660 1875.900 484.260 1881.100 ;
        RECT 529.580 1881.100 580.860 1882.700 ;
        RECT 529.580 1875.900 531.180 1881.100 ;
        RECT 482.660 1874.300 531.180 1875.900 ;
        RECT 579.260 1875.900 580.860 1881.100 ;
        RECT 626.180 1881.100 677.460 1882.700 ;
        RECT 626.180 1875.900 627.780 1881.100 ;
        RECT 579.260 1874.300 627.780 1875.900 ;
        RECT 675.860 1875.900 677.460 1881.100 ;
        RECT 722.780 1881.100 774.060 1882.700 ;
        RECT 722.780 1875.900 724.380 1881.100 ;
        RECT 675.860 1874.300 724.380 1875.900 ;
        RECT 772.460 1875.900 774.060 1881.100 ;
        RECT 819.380 1881.100 870.660 1882.700 ;
        RECT 819.380 1875.900 820.980 1881.100 ;
        RECT 772.460 1874.300 820.980 1875.900 ;
        RECT 869.060 1872.500 870.660 1881.100 ;
        RECT 882.860 1872.500 884.460 1887.900 ;
        RECT 929.780 1882.700 931.380 1887.900 ;
        RECT 979.460 1887.900 1027.980 1889.500 ;
        RECT 929.780 1881.100 967.260 1882.700 ;
        RECT 869.060 1870.900 884.460 1872.500 ;
        RECT 965.660 1872.500 967.260 1881.100 ;
        RECT 979.460 1872.500 981.060 1887.900 ;
        RECT 1026.380 1882.700 1027.980 1887.900 ;
        RECT 1076.060 1887.900 1124.580 1889.500 ;
        RECT 1026.380 1881.100 1063.860 1882.700 ;
        RECT 965.660 1870.900 981.060 1872.500 ;
        RECT 1062.260 1872.500 1063.860 1881.100 ;
        RECT 1076.060 1872.500 1077.660 1887.900 ;
        RECT 1122.980 1882.700 1124.580 1887.900 ;
        RECT 1172.660 1887.900 1221.180 1889.500 ;
        RECT 1122.980 1881.100 1160.460 1882.700 ;
        RECT 1062.260 1870.900 1077.660 1872.500 ;
        RECT 1158.860 1872.500 1160.460 1881.100 ;
        RECT 1172.660 1872.500 1174.260 1887.900 ;
        RECT 1219.580 1882.700 1221.180 1887.900 ;
        RECT 1269.260 1887.900 1317.780 1889.500 ;
        RECT 1219.580 1881.100 1257.060 1882.700 ;
        RECT 1158.860 1870.900 1174.260 1872.500 ;
        RECT 1255.460 1872.500 1257.060 1881.100 ;
        RECT 1269.260 1872.500 1270.860 1887.900 ;
        RECT 1316.180 1882.700 1317.780 1887.900 ;
        RECT 1365.860 1887.900 1414.380 1889.500 ;
        RECT 1316.180 1881.100 1353.660 1882.700 ;
        RECT 1255.460 1870.900 1270.860 1872.500 ;
        RECT 1352.060 1872.500 1353.660 1881.100 ;
        RECT 1365.860 1872.500 1367.460 1887.900 ;
        RECT 1412.780 1882.700 1414.380 1887.900 ;
        RECT 1462.460 1887.900 1510.980 1889.500 ;
        RECT 1412.780 1881.100 1450.260 1882.700 ;
        RECT 1352.060 1870.900 1367.460 1872.500 ;
        RECT 1448.660 1872.500 1450.260 1881.100 ;
        RECT 1462.460 1872.500 1464.060 1887.900 ;
        RECT 1509.380 1882.700 1510.980 1887.900 ;
        RECT 1559.060 1887.900 1607.580 1889.500 ;
        RECT 1509.380 1881.100 1546.860 1882.700 ;
        RECT 1448.660 1870.900 1464.060 1872.500 ;
        RECT 1545.260 1872.500 1546.860 1881.100 ;
        RECT 1559.060 1872.500 1560.660 1887.900 ;
        RECT 1605.980 1882.700 1607.580 1887.900 ;
        RECT 1655.660 1887.900 1704.180 1889.500 ;
        RECT 1605.980 1881.100 1643.460 1882.700 ;
        RECT 1545.260 1870.900 1560.660 1872.500 ;
        RECT 1641.860 1872.500 1643.460 1881.100 ;
        RECT 1655.660 1872.500 1657.260 1887.900 ;
        RECT 1702.580 1882.700 1704.180 1887.900 ;
        RECT 1752.260 1887.900 1800.780 1889.500 ;
        RECT 1702.580 1881.100 1740.060 1882.700 ;
        RECT 1641.860 1870.900 1657.260 1872.500 ;
        RECT 1738.460 1872.500 1740.060 1881.100 ;
        RECT 1752.260 1872.500 1753.860 1887.900 ;
        RECT 1799.180 1882.700 1800.780 1887.900 ;
        RECT 1848.860 1887.900 1897.380 1889.500 ;
        RECT 1799.180 1881.100 1836.660 1882.700 ;
        RECT 1738.460 1870.900 1753.860 1872.500 ;
        RECT 1835.060 1872.500 1836.660 1881.100 ;
        RECT 1848.860 1872.500 1850.460 1887.900 ;
        RECT 1895.780 1882.700 1897.380 1887.900 ;
        RECT 1945.460 1887.900 1993.980 1889.500 ;
        RECT 1895.780 1881.100 1933.260 1882.700 ;
        RECT 1835.060 1870.900 1850.460 1872.500 ;
        RECT 1931.660 1872.500 1933.260 1881.100 ;
        RECT 1945.460 1872.500 1947.060 1887.900 ;
        RECT 1992.380 1882.700 1993.980 1887.900 ;
        RECT 2042.060 1887.900 2090.580 1889.500 ;
        RECT 1992.380 1881.100 2029.860 1882.700 ;
        RECT 1931.660 1870.900 1947.060 1872.500 ;
        RECT 2028.260 1872.500 2029.860 1881.100 ;
        RECT 2042.060 1872.500 2043.660 1887.900 ;
        RECT 2088.980 1882.700 2090.580 1887.900 ;
        RECT 2138.660 1887.900 2187.180 1889.500 ;
        RECT 2088.980 1881.100 2126.460 1882.700 ;
        RECT 2028.260 1870.900 2043.660 1872.500 ;
        RECT 2124.860 1872.500 2126.460 1881.100 ;
        RECT 2138.660 1872.500 2140.260 1887.900 ;
        RECT 2185.580 1882.700 2187.180 1887.900 ;
        RECT 2235.260 1887.900 2283.780 1889.500 ;
        RECT 2185.580 1881.100 2223.060 1882.700 ;
        RECT 2124.860 1870.900 2140.260 1872.500 ;
        RECT 2221.460 1872.500 2223.060 1881.100 ;
        RECT 2235.260 1872.500 2236.860 1887.900 ;
        RECT 2282.180 1882.700 2283.780 1887.900 ;
        RECT 2331.860 1887.900 2374.860 1889.500 ;
        RECT 2282.180 1881.100 2319.660 1882.700 ;
        RECT 2221.460 1870.900 2236.860 1872.500 ;
        RECT 2318.060 1872.500 2319.660 1881.100 ;
        RECT 2331.860 1872.500 2333.460 1887.900 ;
        RECT 2373.260 1886.100 2374.860 1887.900 ;
        RECT 2552.660 1886.100 2554.260 1891.300 ;
        RECT 2373.260 1884.500 2381.300 1886.100 ;
        RECT 2379.700 1882.700 2381.300 1884.500 ;
        RECT 2407.300 1884.500 2430.060 1886.100 ;
        RECT 2407.300 1882.700 2408.900 1884.500 ;
        RECT 2379.700 1881.100 2408.900 1882.700 ;
        RECT 2428.460 1882.700 2430.060 1884.500 ;
        RECT 2455.140 1884.500 2554.260 1886.100 ;
        RECT 2455.140 1882.700 2456.740 1884.500 ;
        RECT 2428.460 1881.100 2456.740 1882.700 ;
        RECT 2599.580 1882.700 2601.180 1891.300 ;
        RECT 2621.660 1887.900 2646.260 1889.500 ;
        RECT 2621.660 1882.700 2623.260 1887.900 ;
        RECT 2599.580 1881.100 2623.260 1882.700 ;
        RECT 2318.060 1870.900 2333.460 1872.500 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2161.610 3017.740 2161.930 3017.800 ;
        RECT 2577.450 3017.740 2577.770 3017.800 ;
        RECT 2161.610 3017.600 2577.770 3017.740 ;
        RECT 2161.610 3017.540 2161.930 3017.600 ;
        RECT 2577.450 3017.540 2577.770 3017.600 ;
        RECT 2577.450 1559.140 2577.770 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 2577.450 1559.000 2901.150 1559.140 ;
        RECT 2577.450 1558.940 2577.770 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 2161.640 3017.540 2161.900 3017.800 ;
        RECT 2577.480 3017.540 2577.740 3017.800 ;
        RECT 2577.480 1558.940 2577.740 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 2161.640 3017.510 2161.900 3017.830 ;
        RECT 2577.480 3017.510 2577.740 3017.830 ;
        RECT 2161.700 3010.000 2161.840 3017.510 ;
        RECT 2161.700 3009.340 2162.050 3010.000 ;
        RECT 2161.770 3006.000 2162.050 3009.340 ;
        RECT 2577.540 1559.230 2577.680 3017.510 ;
        RECT 2577.480 1558.910 2577.740 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2846.090 1787.280 2846.410 1787.340 ;
        RECT 2900.830 1787.280 2901.150 1787.340 ;
        RECT 2846.090 1787.140 2901.150 1787.280 ;
        RECT 2846.090 1787.080 2846.410 1787.140 ;
        RECT 2900.830 1787.080 2901.150 1787.140 ;
      LAYER via ;
        RECT 2846.120 1787.080 2846.380 1787.340 ;
        RECT 2900.860 1787.080 2901.120 1787.340 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1787.370 2901.060 1789.235 ;
        RECT 2846.120 1787.050 2846.380 1787.370 ;
        RECT 2900.860 1787.050 2901.120 1787.370 ;
        RECT 968.530 510.340 968.810 514.000 ;
        RECT 968.460 510.000 968.810 510.340 ;
        RECT 968.460 504.405 968.600 510.000 ;
        RECT 2846.180 504.405 2846.320 1787.050 ;
        RECT 968.390 504.035 968.670 504.405 ;
        RECT 2846.110 504.035 2846.390 504.405 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 968.390 504.080 968.670 504.360 ;
        RECT 2846.110 504.080 2846.390 504.360 ;
      LAYER met3 ;
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 968.365 504.370 968.695 504.385 ;
        RECT 2846.085 504.370 2846.415 504.385 ;
        RECT 968.365 504.070 2846.415 504.370 ;
        RECT 968.365 504.055 968.695 504.070 ;
        RECT 2846.085 504.055 2846.415 504.070 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2583.890 2021.880 2584.210 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 2583.890 2021.740 2901.150 2021.880 ;
        RECT 2583.890 2021.680 2584.210 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
        RECT 1635.370 503.100 1635.690 503.160 ;
        RECT 2583.890 503.100 2584.210 503.160 ;
        RECT 1635.370 502.960 2584.210 503.100 ;
        RECT 1635.370 502.900 1635.690 502.960 ;
        RECT 2583.890 502.900 2584.210 502.960 ;
      LAYER via ;
        RECT 2583.920 2021.680 2584.180 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
        RECT 1635.400 502.900 1635.660 503.160 ;
        RECT 2583.920 502.900 2584.180 503.160 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 2583.920 2021.650 2584.180 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 1635.530 510.340 1635.810 514.000 ;
        RECT 1635.460 510.000 1635.810 510.340 ;
        RECT 1635.460 503.190 1635.600 510.000 ;
        RECT 2583.980 503.190 2584.120 2021.650 ;
        RECT 1635.400 502.870 1635.660 503.190 ;
        RECT 2583.920 502.870 2584.180 503.190 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 655.185 3001.605 655.355 3006.535 ;
      LAYER mcon ;
        RECT 655.185 3006.365 655.355 3006.535 ;
      LAYER met1 ;
        RECT 655.110 3006.520 655.430 3006.580 ;
        RECT 654.915 3006.380 655.430 3006.520 ;
        RECT 655.110 3006.320 655.430 3006.380 ;
        RECT 655.125 3001.760 655.415 3001.805 ;
        RECT 2549.390 3001.760 2549.710 3001.820 ;
        RECT 655.125 3001.620 2549.710 3001.760 ;
        RECT 655.125 3001.575 655.415 3001.620 ;
        RECT 2549.390 3001.560 2549.710 3001.620 ;
        RECT 2549.390 2262.940 2549.710 2263.000 ;
        RECT 2900.830 2262.940 2901.150 2263.000 ;
        RECT 2549.390 2262.800 2901.150 2262.940 ;
        RECT 2549.390 2262.740 2549.710 2262.800 ;
        RECT 2900.830 2262.740 2901.150 2262.800 ;
      LAYER via ;
        RECT 655.140 3006.320 655.400 3006.580 ;
        RECT 2549.420 3001.560 2549.680 3001.820 ;
        RECT 2549.420 2262.740 2549.680 2263.000 ;
        RECT 2900.860 2262.740 2901.120 2263.000 ;
      LAYER met2 ;
        RECT 653.890 3006.690 654.170 3010.000 ;
        RECT 653.890 3006.610 655.340 3006.690 ;
        RECT 653.890 3006.550 655.400 3006.610 ;
        RECT 653.890 3006.000 654.170 3006.550 ;
        RECT 655.140 3006.290 655.400 3006.550 ;
        RECT 2549.420 3001.530 2549.680 3001.850 ;
        RECT 2549.480 2263.030 2549.620 3001.530 ;
        RECT 2549.420 2262.710 2549.680 2263.030 ;
        RECT 2900.860 2262.710 2901.120 2263.030 ;
        RECT 2900.920 2258.805 2901.060 2262.710 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.410 65.520 634.730 65.580 ;
        RECT 1469.770 65.520 1470.090 65.580 ;
        RECT 634.410 65.380 1470.090 65.520 ;
        RECT 634.410 65.320 634.730 65.380 ;
        RECT 1469.770 65.320 1470.090 65.380 ;
      LAYER via ;
        RECT 634.440 65.320 634.700 65.580 ;
        RECT 1469.800 65.320 1470.060 65.580 ;
      LAYER met2 ;
        RECT 1474.530 510.410 1474.810 514.000 ;
        RECT 1469.860 510.270 1474.810 510.410 ;
        RECT 1469.860 65.610 1470.000 510.270 ;
        RECT 1474.530 510.000 1474.810 510.270 ;
        RECT 634.440 65.290 634.700 65.610 ;
        RECT 1469.800 65.290 1470.060 65.610 ;
        RECT 634.500 17.410 634.640 65.290 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.870 972.980 2521.190 973.040 ;
        RECT 2569.630 972.980 2569.950 973.040 ;
        RECT 2520.870 972.840 2569.950 972.980 ;
        RECT 2520.870 972.780 2521.190 972.840 ;
        RECT 2569.630 972.780 2569.950 972.840 ;
        RECT 2421.510 508.540 2421.830 508.600 ;
        RECT 2569.630 508.540 2569.950 508.600 ;
        RECT 2421.510 508.400 2569.950 508.540 ;
        RECT 2421.510 508.340 2421.830 508.400 ;
        RECT 2569.630 508.340 2569.950 508.400 ;
        RECT 2417.370 16.900 2417.690 16.960 ;
        RECT 2421.510 16.900 2421.830 16.960 ;
        RECT 2417.370 16.760 2421.830 16.900 ;
        RECT 2417.370 16.700 2417.690 16.760 ;
        RECT 2421.510 16.700 2421.830 16.760 ;
      LAYER via ;
        RECT 2520.900 972.780 2521.160 973.040 ;
        RECT 2569.660 972.780 2569.920 973.040 ;
        RECT 2421.540 508.340 2421.800 508.600 ;
        RECT 2569.660 508.340 2569.920 508.600 ;
        RECT 2417.400 16.700 2417.660 16.960 ;
        RECT 2421.540 16.700 2421.800 16.960 ;
      LAYER met2 ;
        RECT 2520.890 977.995 2521.170 978.365 ;
        RECT 2520.960 973.070 2521.100 977.995 ;
        RECT 2520.900 972.750 2521.160 973.070 ;
        RECT 2569.660 972.750 2569.920 973.070 ;
        RECT 2569.720 508.630 2569.860 972.750 ;
        RECT 2421.540 508.310 2421.800 508.630 ;
        RECT 2569.660 508.310 2569.920 508.630 ;
        RECT 2421.600 16.990 2421.740 508.310 ;
        RECT 2417.400 16.670 2417.660 16.990 ;
        RECT 2421.540 16.670 2421.800 16.990 ;
        RECT 2417.460 2.400 2417.600 16.670 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 2520.890 978.040 2521.170 978.320 ;
      LAYER met3 ;
        RECT 2506.000 978.330 2510.000 978.480 ;
        RECT 2520.865 978.330 2521.195 978.345 ;
        RECT 2506.000 978.030 2521.195 978.330 ;
        RECT 2506.000 977.880 2510.000 978.030 ;
        RECT 2520.865 978.015 2521.195 978.030 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.710 628.220 2523.030 628.280 ;
        RECT 2548.930 628.220 2549.250 628.280 ;
        RECT 2522.710 628.080 2549.250 628.220 ;
        RECT 2522.710 628.020 2523.030 628.080 ;
        RECT 2548.930 628.020 2549.250 628.080 ;
        RECT 2435.310 508.880 2435.630 508.940 ;
        RECT 2548.930 508.880 2549.250 508.940 ;
        RECT 2435.310 508.740 2549.250 508.880 ;
        RECT 2435.310 508.680 2435.630 508.740 ;
        RECT 2548.930 508.680 2549.250 508.740 ;
        RECT 2434.390 62.120 2434.710 62.180 ;
        RECT 2435.310 62.120 2435.630 62.180 ;
        RECT 2434.390 61.980 2435.630 62.120 ;
        RECT 2434.390 61.920 2434.710 61.980 ;
        RECT 2435.310 61.920 2435.630 61.980 ;
      LAYER via ;
        RECT 2522.740 628.020 2523.000 628.280 ;
        RECT 2548.960 628.020 2549.220 628.280 ;
        RECT 2435.340 508.680 2435.600 508.940 ;
        RECT 2548.960 508.680 2549.220 508.940 ;
        RECT 2434.420 61.920 2434.680 62.180 ;
        RECT 2435.340 61.920 2435.600 62.180 ;
      LAYER met2 ;
        RECT 2522.730 631.195 2523.010 631.565 ;
        RECT 2522.800 628.310 2522.940 631.195 ;
        RECT 2522.740 627.990 2523.000 628.310 ;
        RECT 2548.960 627.990 2549.220 628.310 ;
        RECT 2549.020 508.970 2549.160 627.990 ;
        RECT 2435.340 508.650 2435.600 508.970 ;
        RECT 2548.960 508.650 2549.220 508.970 ;
        RECT 2435.400 62.210 2435.540 508.650 ;
        RECT 2434.420 61.890 2434.680 62.210 ;
        RECT 2435.340 61.890 2435.600 62.210 ;
        RECT 2434.480 19.450 2434.620 61.890 ;
        RECT 2434.480 19.310 2435.080 19.450 ;
        RECT 2434.940 2.400 2435.080 19.310 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 2522.730 631.240 2523.010 631.520 ;
      LAYER met3 ;
        RECT 2506.000 631.530 2510.000 631.680 ;
        RECT 2522.705 631.530 2523.035 631.545 ;
        RECT 2506.000 631.230 2523.035 631.530 ;
        RECT 2506.000 631.080 2510.000 631.230 ;
        RECT 2522.705 631.215 2523.035 631.230 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.310 3017.315 1061.590 3017.685 ;
        RECT 2580.690 3017.315 2580.970 3017.685 ;
        RECT 1061.380 3010.000 1061.520 3017.315 ;
        RECT 1061.380 3009.340 1061.730 3010.000 ;
        RECT 1061.450 3006.000 1061.730 3009.340 ;
        RECT 2580.760 18.885 2580.900 3017.315 ;
        RECT 2452.810 18.515 2453.090 18.885 ;
        RECT 2580.690 18.515 2580.970 18.885 ;
        RECT 2452.880 2.400 2453.020 18.515 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 1061.310 3017.360 1061.590 3017.640 ;
        RECT 2580.690 3017.360 2580.970 3017.640 ;
        RECT 2452.810 18.560 2453.090 18.840 ;
        RECT 2580.690 18.560 2580.970 18.840 ;
      LAYER met3 ;
        RECT 1061.285 3017.650 1061.615 3017.665 ;
        RECT 2580.665 3017.650 2580.995 3017.665 ;
        RECT 1061.285 3017.350 2580.995 3017.650 ;
        RECT 1061.285 3017.335 1061.615 3017.350 ;
        RECT 2580.665 3017.335 2580.995 3017.350 ;
        RECT 2452.785 18.850 2453.115 18.865 ;
        RECT 2580.665 18.850 2580.995 18.865 ;
        RECT 2452.785 18.550 2580.995 18.850 ;
        RECT 2452.785 18.535 2453.115 18.550 ;
        RECT 2580.665 18.535 2580.995 18.550 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2518.645 16.405 2518.815 20.315 ;
        RECT 2542.565 19.465 2542.735 20.315 ;
      LAYER mcon ;
        RECT 2518.645 20.145 2518.815 20.315 ;
        RECT 2542.565 20.145 2542.735 20.315 ;
      LAYER met1 ;
        RECT 2272.010 3018.760 2272.330 3018.820 ;
        RECT 2567.330 3018.760 2567.650 3018.820 ;
        RECT 2272.010 3018.620 2567.650 3018.760 ;
        RECT 2272.010 3018.560 2272.330 3018.620 ;
        RECT 2567.330 3018.560 2567.650 3018.620 ;
        RECT 2518.585 20.300 2518.875 20.345 ;
        RECT 2542.505 20.300 2542.795 20.345 ;
        RECT 2518.585 20.160 2542.795 20.300 ;
        RECT 2518.585 20.115 2518.875 20.160 ;
        RECT 2542.505 20.115 2542.795 20.160 ;
        RECT 2542.505 19.620 2542.795 19.665 ;
        RECT 2567.330 19.620 2567.650 19.680 ;
        RECT 2542.505 19.480 2567.650 19.620 ;
        RECT 2542.505 19.435 2542.795 19.480 ;
        RECT 2567.330 19.420 2567.650 19.480 ;
        RECT 2470.730 16.560 2471.050 16.620 ;
        RECT 2518.585 16.560 2518.875 16.605 ;
        RECT 2470.730 16.420 2518.875 16.560 ;
        RECT 2470.730 16.360 2471.050 16.420 ;
        RECT 2518.585 16.375 2518.875 16.420 ;
      LAYER via ;
        RECT 2272.040 3018.560 2272.300 3018.820 ;
        RECT 2567.360 3018.560 2567.620 3018.820 ;
        RECT 2567.360 19.420 2567.620 19.680 ;
        RECT 2470.760 16.360 2471.020 16.620 ;
      LAYER met2 ;
        RECT 2272.040 3018.530 2272.300 3018.850 ;
        RECT 2567.360 3018.530 2567.620 3018.850 ;
        RECT 2272.100 3010.000 2272.240 3018.530 ;
        RECT 2272.100 3009.340 2272.450 3010.000 ;
        RECT 2272.170 3006.000 2272.450 3009.340 ;
        RECT 2567.420 19.710 2567.560 3018.530 ;
        RECT 2567.360 19.390 2567.620 19.710 ;
        RECT 2470.760 16.330 2471.020 16.650 ;
        RECT 2470.820 2.400 2470.960 16.330 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1815.690 3019.440 1816.010 3019.500 ;
        RECT 2408.630 3019.440 2408.950 3019.500 ;
        RECT 1815.690 3019.300 2408.950 3019.440 ;
        RECT 1815.690 3019.240 1816.010 3019.300 ;
        RECT 2408.630 3019.240 2408.950 3019.300 ;
        RECT 2408.630 3012.300 2408.950 3012.360 ;
        RECT 2588.490 3012.300 2588.810 3012.360 ;
        RECT 2408.630 3012.160 2588.810 3012.300 ;
        RECT 2408.630 3012.100 2408.950 3012.160 ;
        RECT 2588.490 3012.100 2588.810 3012.160 ;
        RECT 2488.670 19.960 2488.990 20.020 ;
        RECT 2588.490 19.960 2588.810 20.020 ;
        RECT 2488.670 19.820 2588.810 19.960 ;
        RECT 2488.670 19.760 2488.990 19.820 ;
        RECT 2588.490 19.760 2588.810 19.820 ;
      LAYER via ;
        RECT 1815.720 3019.240 1815.980 3019.500 ;
        RECT 2408.660 3019.240 2408.920 3019.500 ;
        RECT 2408.660 3012.100 2408.920 3012.360 ;
        RECT 2588.520 3012.100 2588.780 3012.360 ;
        RECT 2488.700 19.760 2488.960 20.020 ;
        RECT 2588.520 19.760 2588.780 20.020 ;
      LAYER met2 ;
        RECT 1815.720 3019.210 1815.980 3019.530 ;
        RECT 2408.660 3019.210 2408.920 3019.530 ;
        RECT 1815.780 3010.000 1815.920 3019.210 ;
        RECT 2408.720 3012.390 2408.860 3019.210 ;
        RECT 2408.660 3012.070 2408.920 3012.390 ;
        RECT 2588.520 3012.070 2588.780 3012.390 ;
        RECT 1815.780 3009.340 1816.130 3010.000 ;
        RECT 1815.850 3006.000 1816.130 3009.340 ;
        RECT 2588.580 20.050 2588.720 3012.070 ;
        RECT 2488.700 19.730 2488.960 20.050 ;
        RECT 2588.520 19.730 2588.780 20.050 ;
        RECT 2488.760 2.400 2488.900 19.730 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 65.520 2132.030 65.580 ;
        RECT 2504.770 65.520 2505.090 65.580 ;
        RECT 2131.710 65.380 2505.090 65.520 ;
        RECT 2131.710 65.320 2132.030 65.380 ;
        RECT 2504.770 65.320 2505.090 65.380 ;
        RECT 2504.770 2.960 2505.090 3.020 ;
        RECT 2506.150 2.960 2506.470 3.020 ;
        RECT 2504.770 2.820 2506.470 2.960 ;
        RECT 2504.770 2.760 2505.090 2.820 ;
        RECT 2506.150 2.760 2506.470 2.820 ;
      LAYER via ;
        RECT 2131.740 65.320 2132.000 65.580 ;
        RECT 2504.800 65.320 2505.060 65.580 ;
        RECT 2504.800 2.760 2505.060 3.020 ;
        RECT 2506.180 2.760 2506.440 3.020 ;
      LAYER met2 ;
        RECT 2129.570 510.410 2129.850 514.000 ;
        RECT 2129.570 510.270 2131.940 510.410 ;
        RECT 2129.570 510.000 2129.850 510.270 ;
        RECT 2131.800 65.610 2131.940 510.270 ;
        RECT 2131.740 65.290 2132.000 65.610 ;
        RECT 2504.800 65.290 2505.060 65.610 ;
        RECT 2504.860 3.050 2505.000 65.290 ;
        RECT 2504.800 2.730 2505.060 3.050 ;
        RECT 2506.180 2.730 2506.440 3.050 ;
        RECT 2506.240 2.400 2506.380 2.730 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 356.570 1552.680 356.890 1552.740 ;
        RECT 393.370 1552.680 393.690 1552.740 ;
        RECT 356.570 1552.540 393.690 1552.680 ;
        RECT 356.570 1552.480 356.890 1552.540 ;
        RECT 393.370 1552.480 393.690 1552.540 ;
      LAYER via ;
        RECT 356.600 1552.480 356.860 1552.740 ;
        RECT 393.400 1552.480 393.660 1552.740 ;
      LAYER met2 ;
        RECT 393.390 1554.635 393.670 1555.005 ;
        RECT 393.460 1552.770 393.600 1554.635 ;
        RECT 356.600 1552.450 356.860 1552.770 ;
        RECT 393.400 1552.450 393.660 1552.770 ;
        RECT 356.660 16.845 356.800 1552.450 ;
        RECT 356.590 16.475 356.870 16.845 ;
        RECT 2524.110 16.475 2524.390 16.845 ;
        RECT 2524.180 2.400 2524.320 16.475 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
      LAYER via2 ;
        RECT 393.390 1554.680 393.670 1554.960 ;
        RECT 356.590 16.520 356.870 16.800 ;
        RECT 2524.110 16.520 2524.390 16.800 ;
      LAYER met3 ;
        RECT 393.365 1554.970 393.695 1554.985 ;
        RECT 410.000 1554.970 414.000 1555.120 ;
        RECT 393.365 1554.670 414.000 1554.970 ;
        RECT 393.365 1554.655 393.695 1554.670 ;
        RECT 410.000 1554.520 414.000 1554.670 ;
        RECT 356.565 16.810 356.895 16.825 ;
        RECT 2524.085 16.810 2524.415 16.825 ;
        RECT 356.565 16.510 2524.415 16.810 ;
        RECT 356.565 16.495 356.895 16.510 ;
        RECT 2524.085 16.495 2524.415 16.510 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1283.740 2520.730 1283.800 ;
        RECT 2540.650 1283.740 2540.970 1283.800 ;
        RECT 2520.410 1283.600 2540.970 1283.740 ;
        RECT 2520.410 1283.540 2520.730 1283.600 ;
        RECT 2540.650 1283.540 2540.970 1283.600 ;
        RECT 2540.650 2.960 2540.970 3.020 ;
        RECT 2542.030 2.960 2542.350 3.020 ;
        RECT 2540.650 2.820 2542.350 2.960 ;
        RECT 2540.650 2.760 2540.970 2.820 ;
        RECT 2542.030 2.760 2542.350 2.820 ;
      LAYER via ;
        RECT 2520.440 1283.540 2520.700 1283.800 ;
        RECT 2540.680 1283.540 2540.940 1283.800 ;
        RECT 2540.680 2.760 2540.940 3.020 ;
        RECT 2542.060 2.760 2542.320 3.020 ;
      LAYER met2 ;
        RECT 2520.430 1288.075 2520.710 1288.445 ;
        RECT 2520.500 1283.830 2520.640 1288.075 ;
        RECT 2520.440 1283.510 2520.700 1283.830 ;
        RECT 2540.680 1283.510 2540.940 1283.830 ;
        RECT 2540.740 3.050 2540.880 1283.510 ;
        RECT 2540.680 2.730 2540.940 3.050 ;
        RECT 2542.060 2.730 2542.320 3.050 ;
        RECT 2542.120 2.400 2542.260 2.730 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1288.120 2520.710 1288.400 ;
      LAYER met3 ;
        RECT 2506.000 1288.410 2510.000 1288.560 ;
        RECT 2520.405 1288.410 2520.735 1288.425 ;
        RECT 2506.000 1288.110 2520.735 1288.410 ;
        RECT 2506.000 1287.960 2510.000 1288.110 ;
        RECT 2520.405 1288.095 2520.735 1288.110 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2564.185 2408.305 2564.355 2456.415 ;
        RECT 2564.185 2311.745 2564.355 2359.855 ;
        RECT 2564.185 2214.845 2564.355 2262.615 ;
        RECT 2564.185 2118.285 2564.355 2166.395 ;
        RECT 2564.185 2021.725 2564.355 2069.835 ;
        RECT 2564.185 1925.505 2564.355 1973.275 ;
        RECT 2564.185 1828.605 2564.355 1876.375 ;
        RECT 2564.185 1732.045 2564.355 1780.155 ;
        RECT 2564.185 1635.485 2564.355 1683.595 ;
        RECT 2564.185 766.105 2564.355 814.215 ;
        RECT 2564.185 669.545 2564.355 717.655 ;
        RECT 2564.185 572.645 2564.355 620.755 ;
        RECT 2563.265 476.085 2563.435 524.195 ;
        RECT 2564.185 379.525 2564.355 427.635 ;
        RECT 2564.185 282.965 2564.355 331.075 ;
        RECT 2564.185 186.405 2564.355 234.515 ;
        RECT 2562.345 48.365 2562.515 137.955 ;
      LAYER mcon ;
        RECT 2564.185 2456.245 2564.355 2456.415 ;
        RECT 2564.185 2359.685 2564.355 2359.855 ;
        RECT 2564.185 2262.445 2564.355 2262.615 ;
        RECT 2564.185 2166.225 2564.355 2166.395 ;
        RECT 2564.185 2069.665 2564.355 2069.835 ;
        RECT 2564.185 1973.105 2564.355 1973.275 ;
        RECT 2564.185 1876.205 2564.355 1876.375 ;
        RECT 2564.185 1779.985 2564.355 1780.155 ;
        RECT 2564.185 1683.425 2564.355 1683.595 ;
        RECT 2564.185 814.045 2564.355 814.215 ;
        RECT 2564.185 717.485 2564.355 717.655 ;
        RECT 2564.185 620.585 2564.355 620.755 ;
        RECT 2563.265 524.025 2563.435 524.195 ;
        RECT 2564.185 427.465 2564.355 427.635 ;
        RECT 2564.185 330.905 2564.355 331.075 ;
        RECT 2564.185 234.345 2564.355 234.515 ;
        RECT 2562.345 137.785 2562.515 137.955 ;
      LAYER met1 ;
        RECT 2396.210 3018.420 2396.530 3018.480 ;
        RECT 2511.210 3018.420 2511.530 3018.480 ;
        RECT 2396.210 3018.280 2511.530 3018.420 ;
        RECT 2396.210 3018.220 2396.530 3018.280 ;
        RECT 2511.210 3018.220 2511.530 3018.280 ;
        RECT 2511.210 2984.080 2511.530 2984.140 ;
        RECT 2564.110 2984.080 2564.430 2984.140 ;
        RECT 2511.210 2983.940 2564.430 2984.080 ;
        RECT 2511.210 2983.880 2511.530 2983.940 ;
        RECT 2564.110 2983.880 2564.430 2983.940 ;
        RECT 2564.110 2794.700 2564.430 2794.760 ;
        RECT 2565.030 2794.700 2565.350 2794.760 ;
        RECT 2564.110 2794.560 2565.350 2794.700 ;
        RECT 2564.110 2794.500 2564.430 2794.560 ;
        RECT 2565.030 2794.500 2565.350 2794.560 ;
        RECT 2564.110 2656.660 2564.430 2656.720 ;
        RECT 2565.030 2656.660 2565.350 2656.720 ;
        RECT 2564.110 2656.520 2565.350 2656.660 ;
        RECT 2564.110 2656.460 2564.430 2656.520 ;
        RECT 2565.030 2656.460 2565.350 2656.520 ;
        RECT 2564.110 2649.520 2564.430 2649.580 ;
        RECT 2565.030 2649.520 2565.350 2649.580 ;
        RECT 2564.110 2649.380 2565.350 2649.520 ;
        RECT 2564.110 2649.320 2564.430 2649.380 ;
        RECT 2565.030 2649.320 2565.350 2649.380 ;
        RECT 2564.110 2560.100 2564.430 2560.160 ;
        RECT 2565.030 2560.100 2565.350 2560.160 ;
        RECT 2564.110 2559.960 2565.350 2560.100 ;
        RECT 2564.110 2559.900 2564.430 2559.960 ;
        RECT 2565.030 2559.900 2565.350 2559.960 ;
        RECT 2564.110 2552.960 2564.430 2553.020 ;
        RECT 2565.030 2552.960 2565.350 2553.020 ;
        RECT 2564.110 2552.820 2565.350 2552.960 ;
        RECT 2564.110 2552.760 2564.430 2552.820 ;
        RECT 2565.030 2552.760 2565.350 2552.820 ;
        RECT 2564.110 2456.400 2564.430 2456.460 ;
        RECT 2563.915 2456.260 2564.430 2456.400 ;
        RECT 2564.110 2456.200 2564.430 2456.260 ;
        RECT 2564.110 2408.460 2564.430 2408.520 ;
        RECT 2563.915 2408.320 2564.430 2408.460 ;
        RECT 2564.110 2408.260 2564.430 2408.320 ;
        RECT 2564.110 2359.840 2564.430 2359.900 ;
        RECT 2563.915 2359.700 2564.430 2359.840 ;
        RECT 2564.110 2359.640 2564.430 2359.700 ;
        RECT 2564.110 2311.900 2564.430 2311.960 ;
        RECT 2563.915 2311.760 2564.430 2311.900 ;
        RECT 2564.110 2311.700 2564.430 2311.760 ;
        RECT 2564.110 2262.600 2564.430 2262.660 ;
        RECT 2563.915 2262.460 2564.430 2262.600 ;
        RECT 2564.110 2262.400 2564.430 2262.460 ;
        RECT 2564.110 2215.000 2564.430 2215.060 ;
        RECT 2563.915 2214.860 2564.430 2215.000 ;
        RECT 2564.110 2214.800 2564.430 2214.860 ;
        RECT 2564.110 2166.380 2564.430 2166.440 ;
        RECT 2563.915 2166.240 2564.430 2166.380 ;
        RECT 2564.110 2166.180 2564.430 2166.240 ;
        RECT 2564.110 2118.440 2564.430 2118.500 ;
        RECT 2563.915 2118.300 2564.430 2118.440 ;
        RECT 2564.110 2118.240 2564.430 2118.300 ;
        RECT 2564.110 2069.820 2564.430 2069.880 ;
        RECT 2563.915 2069.680 2564.430 2069.820 ;
        RECT 2564.110 2069.620 2564.430 2069.680 ;
        RECT 2564.110 2021.880 2564.430 2021.940 ;
        RECT 2563.915 2021.740 2564.430 2021.880 ;
        RECT 2564.110 2021.680 2564.430 2021.740 ;
        RECT 2564.110 1973.260 2564.430 1973.320 ;
        RECT 2563.915 1973.120 2564.430 1973.260 ;
        RECT 2564.110 1973.060 2564.430 1973.120 ;
        RECT 2564.110 1925.660 2564.430 1925.720 ;
        RECT 2563.915 1925.520 2564.430 1925.660 ;
        RECT 2564.110 1925.460 2564.430 1925.520 ;
        RECT 2564.110 1876.360 2564.430 1876.420 ;
        RECT 2563.915 1876.220 2564.430 1876.360 ;
        RECT 2564.110 1876.160 2564.430 1876.220 ;
        RECT 2564.110 1828.760 2564.430 1828.820 ;
        RECT 2563.915 1828.620 2564.430 1828.760 ;
        RECT 2564.110 1828.560 2564.430 1828.620 ;
        RECT 2564.110 1787.760 2564.430 1788.020 ;
        RECT 2564.200 1787.340 2564.340 1787.760 ;
        RECT 2564.110 1787.080 2564.430 1787.340 ;
        RECT 2564.110 1780.140 2564.430 1780.200 ;
        RECT 2563.915 1780.000 2564.430 1780.140 ;
        RECT 2564.110 1779.940 2564.430 1780.000 ;
        RECT 2564.110 1732.200 2564.430 1732.260 ;
        RECT 2563.915 1732.060 2564.430 1732.200 ;
        RECT 2564.110 1732.000 2564.430 1732.060 ;
        RECT 2564.110 1683.580 2564.430 1683.640 ;
        RECT 2563.915 1683.440 2564.430 1683.580 ;
        RECT 2564.110 1683.380 2564.430 1683.440 ;
        RECT 2564.110 1635.640 2564.430 1635.700 ;
        RECT 2563.915 1635.500 2564.430 1635.640 ;
        RECT 2564.110 1635.440 2564.430 1635.500 ;
        RECT 2564.110 1587.020 2564.430 1587.080 ;
        RECT 2564.570 1587.020 2564.890 1587.080 ;
        RECT 2564.110 1586.880 2564.890 1587.020 ;
        RECT 2564.110 1586.820 2564.430 1586.880 ;
        RECT 2564.570 1586.820 2564.890 1586.880 ;
        RECT 2564.110 1490.460 2564.430 1490.520 ;
        RECT 2564.570 1490.460 2564.890 1490.520 ;
        RECT 2564.110 1490.320 2564.890 1490.460 ;
        RECT 2564.110 1490.260 2564.430 1490.320 ;
        RECT 2564.570 1490.260 2564.890 1490.320 ;
        RECT 2564.110 1345.620 2564.430 1345.680 ;
        RECT 2565.030 1345.620 2565.350 1345.680 ;
        RECT 2564.110 1345.480 2565.350 1345.620 ;
        RECT 2564.110 1345.420 2564.430 1345.480 ;
        RECT 2565.030 1345.420 2565.350 1345.480 ;
        RECT 2564.110 1249.400 2564.430 1249.460 ;
        RECT 2565.030 1249.400 2565.350 1249.460 ;
        RECT 2564.110 1249.260 2565.350 1249.400 ;
        RECT 2564.110 1249.200 2564.430 1249.260 ;
        RECT 2565.030 1249.200 2565.350 1249.260 ;
        RECT 2564.110 1152.500 2564.430 1152.560 ;
        RECT 2565.030 1152.500 2565.350 1152.560 ;
        RECT 2564.110 1152.360 2565.350 1152.500 ;
        RECT 2564.110 1152.300 2564.430 1152.360 ;
        RECT 2565.030 1152.300 2565.350 1152.360 ;
        RECT 2564.110 1007.320 2564.430 1007.380 ;
        RECT 2565.030 1007.320 2565.350 1007.380 ;
        RECT 2564.110 1007.180 2565.350 1007.320 ;
        RECT 2564.110 1007.120 2564.430 1007.180 ;
        RECT 2565.030 1007.120 2565.350 1007.180 ;
        RECT 2564.110 910.760 2564.430 910.820 ;
        RECT 2565.030 910.760 2565.350 910.820 ;
        RECT 2564.110 910.620 2565.350 910.760 ;
        RECT 2564.110 910.560 2564.430 910.620 ;
        RECT 2565.030 910.560 2565.350 910.620 ;
        RECT 2564.110 814.200 2564.430 814.260 ;
        RECT 2563.915 814.060 2564.430 814.200 ;
        RECT 2564.110 814.000 2564.430 814.060 ;
        RECT 2564.110 766.260 2564.430 766.320 ;
        RECT 2563.915 766.120 2564.430 766.260 ;
        RECT 2564.110 766.060 2564.430 766.120 ;
        RECT 2564.110 717.640 2564.430 717.700 ;
        RECT 2563.915 717.500 2564.430 717.640 ;
        RECT 2564.110 717.440 2564.430 717.500 ;
        RECT 2564.110 669.700 2564.430 669.760 ;
        RECT 2563.915 669.560 2564.430 669.700 ;
        RECT 2564.110 669.500 2564.430 669.560 ;
        RECT 2564.110 620.740 2564.430 620.800 ;
        RECT 2563.915 620.600 2564.430 620.740 ;
        RECT 2564.110 620.540 2564.430 620.600 ;
        RECT 2564.110 572.800 2564.430 572.860 ;
        RECT 2563.915 572.660 2564.430 572.800 ;
        RECT 2564.110 572.600 2564.430 572.660 ;
        RECT 2563.205 524.180 2563.495 524.225 ;
        RECT 2564.110 524.180 2564.430 524.240 ;
        RECT 2563.205 524.040 2564.430 524.180 ;
        RECT 2563.205 523.995 2563.495 524.040 ;
        RECT 2564.110 523.980 2564.430 524.040 ;
        RECT 2563.205 476.240 2563.495 476.285 ;
        RECT 2563.650 476.240 2563.970 476.300 ;
        RECT 2563.205 476.100 2563.970 476.240 ;
        RECT 2563.205 476.055 2563.495 476.100 ;
        RECT 2563.650 476.040 2563.970 476.100 ;
        RECT 2563.650 435.100 2563.970 435.160 ;
        RECT 2564.110 435.100 2564.430 435.160 ;
        RECT 2563.650 434.960 2564.430 435.100 ;
        RECT 2563.650 434.900 2563.970 434.960 ;
        RECT 2564.110 434.900 2564.430 434.960 ;
        RECT 2564.110 427.620 2564.430 427.680 ;
        RECT 2563.915 427.480 2564.430 427.620 ;
        RECT 2564.110 427.420 2564.430 427.480 ;
        RECT 2564.110 379.680 2564.430 379.740 ;
        RECT 2563.915 379.540 2564.430 379.680 ;
        RECT 2564.110 379.480 2564.430 379.540 ;
        RECT 2564.110 331.060 2564.430 331.120 ;
        RECT 2563.915 330.920 2564.430 331.060 ;
        RECT 2564.110 330.860 2564.430 330.920 ;
        RECT 2564.110 283.120 2564.430 283.180 ;
        RECT 2563.915 282.980 2564.430 283.120 ;
        RECT 2564.110 282.920 2564.430 282.980 ;
        RECT 2564.110 234.500 2564.430 234.560 ;
        RECT 2563.915 234.360 2564.430 234.500 ;
        RECT 2564.110 234.300 2564.430 234.360 ;
        RECT 2564.110 186.560 2564.430 186.620 ;
        RECT 2563.915 186.420 2564.430 186.560 ;
        RECT 2564.110 186.360 2564.430 186.420 ;
        RECT 2562.285 137.940 2562.575 137.985 ;
        RECT 2564.110 137.940 2564.430 138.000 ;
        RECT 2562.285 137.800 2564.430 137.940 ;
        RECT 2562.285 137.755 2562.575 137.800 ;
        RECT 2564.110 137.740 2564.430 137.800 ;
        RECT 2562.270 48.520 2562.590 48.580 ;
        RECT 2562.075 48.380 2562.590 48.520 ;
        RECT 2562.270 48.320 2562.590 48.380 ;
        RECT 2559.970 13.840 2560.290 13.900 ;
        RECT 2562.730 13.840 2563.050 13.900 ;
        RECT 2559.970 13.700 2563.050 13.840 ;
        RECT 2559.970 13.640 2560.290 13.700 ;
        RECT 2562.730 13.640 2563.050 13.700 ;
      LAYER via ;
        RECT 2396.240 3018.220 2396.500 3018.480 ;
        RECT 2511.240 3018.220 2511.500 3018.480 ;
        RECT 2511.240 2983.880 2511.500 2984.140 ;
        RECT 2564.140 2983.880 2564.400 2984.140 ;
        RECT 2564.140 2794.500 2564.400 2794.760 ;
        RECT 2565.060 2794.500 2565.320 2794.760 ;
        RECT 2564.140 2656.460 2564.400 2656.720 ;
        RECT 2565.060 2656.460 2565.320 2656.720 ;
        RECT 2564.140 2649.320 2564.400 2649.580 ;
        RECT 2565.060 2649.320 2565.320 2649.580 ;
        RECT 2564.140 2559.900 2564.400 2560.160 ;
        RECT 2565.060 2559.900 2565.320 2560.160 ;
        RECT 2564.140 2552.760 2564.400 2553.020 ;
        RECT 2565.060 2552.760 2565.320 2553.020 ;
        RECT 2564.140 2456.200 2564.400 2456.460 ;
        RECT 2564.140 2408.260 2564.400 2408.520 ;
        RECT 2564.140 2359.640 2564.400 2359.900 ;
        RECT 2564.140 2311.700 2564.400 2311.960 ;
        RECT 2564.140 2262.400 2564.400 2262.660 ;
        RECT 2564.140 2214.800 2564.400 2215.060 ;
        RECT 2564.140 2166.180 2564.400 2166.440 ;
        RECT 2564.140 2118.240 2564.400 2118.500 ;
        RECT 2564.140 2069.620 2564.400 2069.880 ;
        RECT 2564.140 2021.680 2564.400 2021.940 ;
        RECT 2564.140 1973.060 2564.400 1973.320 ;
        RECT 2564.140 1925.460 2564.400 1925.720 ;
        RECT 2564.140 1876.160 2564.400 1876.420 ;
        RECT 2564.140 1828.560 2564.400 1828.820 ;
        RECT 2564.140 1787.760 2564.400 1788.020 ;
        RECT 2564.140 1787.080 2564.400 1787.340 ;
        RECT 2564.140 1779.940 2564.400 1780.200 ;
        RECT 2564.140 1732.000 2564.400 1732.260 ;
        RECT 2564.140 1683.380 2564.400 1683.640 ;
        RECT 2564.140 1635.440 2564.400 1635.700 ;
        RECT 2564.140 1586.820 2564.400 1587.080 ;
        RECT 2564.600 1586.820 2564.860 1587.080 ;
        RECT 2564.140 1490.260 2564.400 1490.520 ;
        RECT 2564.600 1490.260 2564.860 1490.520 ;
        RECT 2564.140 1345.420 2564.400 1345.680 ;
        RECT 2565.060 1345.420 2565.320 1345.680 ;
        RECT 2564.140 1249.200 2564.400 1249.460 ;
        RECT 2565.060 1249.200 2565.320 1249.460 ;
        RECT 2564.140 1152.300 2564.400 1152.560 ;
        RECT 2565.060 1152.300 2565.320 1152.560 ;
        RECT 2564.140 1007.120 2564.400 1007.380 ;
        RECT 2565.060 1007.120 2565.320 1007.380 ;
        RECT 2564.140 910.560 2564.400 910.820 ;
        RECT 2565.060 910.560 2565.320 910.820 ;
        RECT 2564.140 814.000 2564.400 814.260 ;
        RECT 2564.140 766.060 2564.400 766.320 ;
        RECT 2564.140 717.440 2564.400 717.700 ;
        RECT 2564.140 669.500 2564.400 669.760 ;
        RECT 2564.140 620.540 2564.400 620.800 ;
        RECT 2564.140 572.600 2564.400 572.860 ;
        RECT 2564.140 523.980 2564.400 524.240 ;
        RECT 2563.680 476.040 2563.940 476.300 ;
        RECT 2563.680 434.900 2563.940 435.160 ;
        RECT 2564.140 434.900 2564.400 435.160 ;
        RECT 2564.140 427.420 2564.400 427.680 ;
        RECT 2564.140 379.480 2564.400 379.740 ;
        RECT 2564.140 330.860 2564.400 331.120 ;
        RECT 2564.140 282.920 2564.400 283.180 ;
        RECT 2564.140 234.300 2564.400 234.560 ;
        RECT 2564.140 186.360 2564.400 186.620 ;
        RECT 2564.140 137.740 2564.400 138.000 ;
        RECT 2562.300 48.320 2562.560 48.580 ;
        RECT 2560.000 13.640 2560.260 13.900 ;
        RECT 2562.760 13.640 2563.020 13.900 ;
      LAYER met2 ;
        RECT 2396.240 3018.190 2396.500 3018.510 ;
        RECT 2511.240 3018.190 2511.500 3018.510 ;
        RECT 2396.300 3010.000 2396.440 3018.190 ;
        RECT 2396.300 3009.340 2396.650 3010.000 ;
        RECT 2396.370 3006.000 2396.650 3009.340 ;
        RECT 2511.300 2984.170 2511.440 3018.190 ;
        RECT 2511.240 2983.850 2511.500 2984.170 ;
        RECT 2564.140 2983.850 2564.400 2984.170 ;
        RECT 2564.200 2851.085 2564.340 2983.850 ;
        RECT 2564.130 2850.715 2564.410 2851.085 ;
        RECT 2564.130 2850.035 2564.410 2850.405 ;
        RECT 2564.200 2842.925 2564.340 2850.035 ;
        RECT 2564.130 2842.555 2564.410 2842.925 ;
        RECT 2565.050 2842.555 2565.330 2842.925 ;
        RECT 2565.120 2794.790 2565.260 2842.555 ;
        RECT 2564.140 2794.470 2564.400 2794.790 ;
        RECT 2565.060 2794.470 2565.320 2794.790 ;
        RECT 2564.200 2746.365 2564.340 2794.470 ;
        RECT 2564.130 2745.995 2564.410 2746.365 ;
        RECT 2565.050 2745.995 2565.330 2746.365 ;
        RECT 2565.120 2656.750 2565.260 2745.995 ;
        RECT 2564.140 2656.430 2564.400 2656.750 ;
        RECT 2565.060 2656.430 2565.320 2656.750 ;
        RECT 2564.200 2649.610 2564.340 2656.430 ;
        RECT 2564.140 2649.290 2564.400 2649.610 ;
        RECT 2565.060 2649.290 2565.320 2649.610 ;
        RECT 2565.120 2560.190 2565.260 2649.290 ;
        RECT 2564.140 2559.870 2564.400 2560.190 ;
        RECT 2565.060 2559.870 2565.320 2560.190 ;
        RECT 2564.200 2553.050 2564.340 2559.870 ;
        RECT 2564.140 2552.730 2564.400 2553.050 ;
        RECT 2565.060 2552.730 2565.320 2553.050 ;
        RECT 2565.120 2504.965 2565.260 2552.730 ;
        RECT 2564.130 2504.595 2564.410 2504.965 ;
        RECT 2565.050 2504.595 2565.330 2504.965 ;
        RECT 2564.200 2456.490 2564.340 2504.595 ;
        RECT 2564.140 2456.170 2564.400 2456.490 ;
        RECT 2564.140 2408.230 2564.400 2408.550 ;
        RECT 2564.200 2359.930 2564.340 2408.230 ;
        RECT 2564.140 2359.610 2564.400 2359.930 ;
        RECT 2564.140 2311.670 2564.400 2311.990 ;
        RECT 2564.200 2262.690 2564.340 2311.670 ;
        RECT 2564.140 2262.370 2564.400 2262.690 ;
        RECT 2564.140 2214.770 2564.400 2215.090 ;
        RECT 2564.200 2166.470 2564.340 2214.770 ;
        RECT 2564.140 2166.150 2564.400 2166.470 ;
        RECT 2564.140 2118.210 2564.400 2118.530 ;
        RECT 2564.200 2069.910 2564.340 2118.210 ;
        RECT 2564.140 2069.590 2564.400 2069.910 ;
        RECT 2564.140 2021.650 2564.400 2021.970 ;
        RECT 2564.200 1973.350 2564.340 2021.650 ;
        RECT 2564.140 1973.030 2564.400 1973.350 ;
        RECT 2564.140 1925.430 2564.400 1925.750 ;
        RECT 2564.200 1885.370 2564.340 1925.430 ;
        RECT 2564.200 1885.230 2564.800 1885.370 ;
        RECT 2564.660 1884.010 2564.800 1885.230 ;
        RECT 2564.200 1883.870 2564.800 1884.010 ;
        RECT 2564.200 1876.450 2564.340 1883.870 ;
        RECT 2564.140 1876.130 2564.400 1876.450 ;
        RECT 2564.140 1828.530 2564.400 1828.850 ;
        RECT 2564.200 1788.050 2564.340 1828.530 ;
        RECT 2564.140 1787.730 2564.400 1788.050 ;
        RECT 2564.140 1787.050 2564.400 1787.370 ;
        RECT 2564.200 1780.230 2564.340 1787.050 ;
        RECT 2564.140 1779.910 2564.400 1780.230 ;
        RECT 2564.140 1731.970 2564.400 1732.290 ;
        RECT 2564.200 1683.670 2564.340 1731.970 ;
        RECT 2564.140 1683.350 2564.400 1683.670 ;
        RECT 2564.140 1635.410 2564.400 1635.730 ;
        RECT 2564.200 1587.110 2564.340 1635.410 ;
        RECT 2564.140 1586.790 2564.400 1587.110 ;
        RECT 2564.600 1586.790 2564.860 1587.110 ;
        RECT 2564.660 1497.770 2564.800 1586.790 ;
        RECT 2564.200 1497.630 2564.800 1497.770 ;
        RECT 2564.200 1490.550 2564.340 1497.630 ;
        RECT 2564.140 1490.230 2564.400 1490.550 ;
        RECT 2564.600 1490.230 2564.860 1490.550 ;
        RECT 2564.660 1401.210 2564.800 1490.230 ;
        RECT 2564.200 1401.070 2564.800 1401.210 ;
        RECT 2564.200 1393.845 2564.340 1401.070 ;
        RECT 2564.130 1393.475 2564.410 1393.845 ;
        RECT 2565.050 1393.475 2565.330 1393.845 ;
        RECT 2565.120 1345.710 2565.260 1393.475 ;
        RECT 2564.140 1345.390 2564.400 1345.710 ;
        RECT 2565.060 1345.390 2565.320 1345.710 ;
        RECT 2564.200 1305.330 2564.340 1345.390 ;
        RECT 2564.200 1305.190 2564.800 1305.330 ;
        RECT 2564.660 1304.650 2564.800 1305.190 ;
        RECT 2564.200 1304.510 2564.800 1304.650 ;
        RECT 2564.200 1297.285 2564.340 1304.510 ;
        RECT 2564.130 1296.915 2564.410 1297.285 ;
        RECT 2565.050 1296.915 2565.330 1297.285 ;
        RECT 2565.120 1249.490 2565.260 1296.915 ;
        RECT 2564.140 1249.170 2564.400 1249.490 ;
        RECT 2565.060 1249.170 2565.320 1249.490 ;
        RECT 2564.200 1200.725 2564.340 1249.170 ;
        RECT 2564.130 1200.355 2564.410 1200.725 ;
        RECT 2565.050 1200.355 2565.330 1200.725 ;
        RECT 2565.120 1152.590 2565.260 1200.355 ;
        RECT 2564.140 1152.270 2564.400 1152.590 ;
        RECT 2565.060 1152.270 2565.320 1152.590 ;
        RECT 2564.200 1104.165 2564.340 1152.270 ;
        RECT 2564.130 1103.795 2564.410 1104.165 ;
        RECT 2565.050 1103.795 2565.330 1104.165 ;
        RECT 2565.120 1055.885 2565.260 1103.795 ;
        RECT 2564.130 1055.515 2564.410 1055.885 ;
        RECT 2565.050 1055.515 2565.330 1055.885 ;
        RECT 2564.200 1007.410 2564.340 1055.515 ;
        RECT 2564.140 1007.090 2564.400 1007.410 ;
        RECT 2565.060 1007.090 2565.320 1007.410 ;
        RECT 2565.120 959.325 2565.260 1007.090 ;
        RECT 2564.130 958.955 2564.410 959.325 ;
        RECT 2565.050 958.955 2565.330 959.325 ;
        RECT 2564.200 910.850 2564.340 958.955 ;
        RECT 2564.140 910.530 2564.400 910.850 ;
        RECT 2565.060 910.530 2565.320 910.850 ;
        RECT 2565.120 862.765 2565.260 910.530 ;
        RECT 2564.130 862.395 2564.410 862.765 ;
        RECT 2565.050 862.395 2565.330 862.765 ;
        RECT 2564.200 814.290 2564.340 862.395 ;
        RECT 2564.140 813.970 2564.400 814.290 ;
        RECT 2564.140 766.030 2564.400 766.350 ;
        RECT 2564.200 717.730 2564.340 766.030 ;
        RECT 2564.140 717.410 2564.400 717.730 ;
        RECT 2564.140 669.470 2564.400 669.790 ;
        RECT 2564.200 620.830 2564.340 669.470 ;
        RECT 2564.140 620.510 2564.400 620.830 ;
        RECT 2564.140 572.570 2564.400 572.890 ;
        RECT 2564.200 524.270 2564.340 572.570 ;
        RECT 2564.140 523.950 2564.400 524.270 ;
        RECT 2563.680 476.010 2563.940 476.330 ;
        RECT 2563.740 435.190 2563.880 476.010 ;
        RECT 2563.680 434.870 2563.940 435.190 ;
        RECT 2564.140 434.870 2564.400 435.190 ;
        RECT 2564.200 427.710 2564.340 434.870 ;
        RECT 2564.140 427.390 2564.400 427.710 ;
        RECT 2564.140 379.450 2564.400 379.770 ;
        RECT 2564.200 331.150 2564.340 379.450 ;
        RECT 2564.140 330.830 2564.400 331.150 ;
        RECT 2564.140 282.890 2564.400 283.210 ;
        RECT 2564.200 234.590 2564.340 282.890 ;
        RECT 2564.140 234.270 2564.400 234.590 ;
        RECT 2564.140 186.330 2564.400 186.650 ;
        RECT 2564.200 138.030 2564.340 186.330 ;
        RECT 2564.140 137.710 2564.400 138.030 ;
        RECT 2562.300 48.290 2562.560 48.610 ;
        RECT 2562.360 48.010 2562.500 48.290 ;
        RECT 2562.360 47.870 2562.960 48.010 ;
        RECT 2562.820 13.930 2562.960 47.870 ;
        RECT 2560.000 13.610 2560.260 13.930 ;
        RECT 2562.760 13.610 2563.020 13.930 ;
        RECT 2560.060 2.400 2560.200 13.610 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
      LAYER via2 ;
        RECT 2564.130 2850.760 2564.410 2851.040 ;
        RECT 2564.130 2850.080 2564.410 2850.360 ;
        RECT 2564.130 2842.600 2564.410 2842.880 ;
        RECT 2565.050 2842.600 2565.330 2842.880 ;
        RECT 2564.130 2746.040 2564.410 2746.320 ;
        RECT 2565.050 2746.040 2565.330 2746.320 ;
        RECT 2564.130 2504.640 2564.410 2504.920 ;
        RECT 2565.050 2504.640 2565.330 2504.920 ;
        RECT 2564.130 1393.520 2564.410 1393.800 ;
        RECT 2565.050 1393.520 2565.330 1393.800 ;
        RECT 2564.130 1296.960 2564.410 1297.240 ;
        RECT 2565.050 1296.960 2565.330 1297.240 ;
        RECT 2564.130 1200.400 2564.410 1200.680 ;
        RECT 2565.050 1200.400 2565.330 1200.680 ;
        RECT 2564.130 1103.840 2564.410 1104.120 ;
        RECT 2565.050 1103.840 2565.330 1104.120 ;
        RECT 2564.130 1055.560 2564.410 1055.840 ;
        RECT 2565.050 1055.560 2565.330 1055.840 ;
        RECT 2564.130 959.000 2564.410 959.280 ;
        RECT 2565.050 959.000 2565.330 959.280 ;
        RECT 2564.130 862.440 2564.410 862.720 ;
        RECT 2565.050 862.440 2565.330 862.720 ;
      LAYER met3 ;
        RECT 2564.105 2851.050 2564.435 2851.065 ;
        RECT 2563.430 2850.750 2564.435 2851.050 ;
        RECT 2563.430 2850.370 2563.730 2850.750 ;
        RECT 2564.105 2850.735 2564.435 2850.750 ;
        RECT 2564.105 2850.370 2564.435 2850.385 ;
        RECT 2563.430 2850.070 2564.435 2850.370 ;
        RECT 2564.105 2850.055 2564.435 2850.070 ;
        RECT 2564.105 2842.890 2564.435 2842.905 ;
        RECT 2565.025 2842.890 2565.355 2842.905 ;
        RECT 2564.105 2842.590 2565.355 2842.890 ;
        RECT 2564.105 2842.575 2564.435 2842.590 ;
        RECT 2565.025 2842.575 2565.355 2842.590 ;
        RECT 2564.105 2746.330 2564.435 2746.345 ;
        RECT 2565.025 2746.330 2565.355 2746.345 ;
        RECT 2564.105 2746.030 2565.355 2746.330 ;
        RECT 2564.105 2746.015 2564.435 2746.030 ;
        RECT 2565.025 2746.015 2565.355 2746.030 ;
        RECT 2564.105 2504.930 2564.435 2504.945 ;
        RECT 2565.025 2504.930 2565.355 2504.945 ;
        RECT 2564.105 2504.630 2565.355 2504.930 ;
        RECT 2564.105 2504.615 2564.435 2504.630 ;
        RECT 2565.025 2504.615 2565.355 2504.630 ;
        RECT 2564.105 1393.810 2564.435 1393.825 ;
        RECT 2565.025 1393.810 2565.355 1393.825 ;
        RECT 2564.105 1393.510 2565.355 1393.810 ;
        RECT 2564.105 1393.495 2564.435 1393.510 ;
        RECT 2565.025 1393.495 2565.355 1393.510 ;
        RECT 2564.105 1297.250 2564.435 1297.265 ;
        RECT 2565.025 1297.250 2565.355 1297.265 ;
        RECT 2564.105 1296.950 2565.355 1297.250 ;
        RECT 2564.105 1296.935 2564.435 1296.950 ;
        RECT 2565.025 1296.935 2565.355 1296.950 ;
        RECT 2564.105 1200.690 2564.435 1200.705 ;
        RECT 2565.025 1200.690 2565.355 1200.705 ;
        RECT 2564.105 1200.390 2565.355 1200.690 ;
        RECT 2564.105 1200.375 2564.435 1200.390 ;
        RECT 2565.025 1200.375 2565.355 1200.390 ;
        RECT 2564.105 1104.130 2564.435 1104.145 ;
        RECT 2565.025 1104.130 2565.355 1104.145 ;
        RECT 2564.105 1103.830 2565.355 1104.130 ;
        RECT 2564.105 1103.815 2564.435 1103.830 ;
        RECT 2565.025 1103.815 2565.355 1103.830 ;
        RECT 2564.105 1055.850 2564.435 1055.865 ;
        RECT 2565.025 1055.850 2565.355 1055.865 ;
        RECT 2564.105 1055.550 2565.355 1055.850 ;
        RECT 2564.105 1055.535 2564.435 1055.550 ;
        RECT 2565.025 1055.535 2565.355 1055.550 ;
        RECT 2564.105 959.290 2564.435 959.305 ;
        RECT 2565.025 959.290 2565.355 959.305 ;
        RECT 2564.105 958.990 2565.355 959.290 ;
        RECT 2564.105 958.975 2564.435 958.990 ;
        RECT 2565.025 958.975 2565.355 958.990 ;
        RECT 2564.105 862.730 2564.435 862.745 ;
        RECT 2565.025 862.730 2565.355 862.745 ;
        RECT 2564.105 862.430 2565.355 862.730 ;
        RECT 2564.105 862.415 2564.435 862.430 ;
        RECT 2565.025 862.415 2565.355 862.430 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 363.930 1407.840 364.250 1407.900 ;
        RECT 393.370 1407.840 393.690 1407.900 ;
        RECT 363.930 1407.700 393.690 1407.840 ;
        RECT 363.930 1407.640 364.250 1407.700 ;
        RECT 393.370 1407.640 393.690 1407.700 ;
        RECT 2577.910 17.580 2578.230 17.640 ;
        RECT 364.940 17.440 2578.230 17.580 ;
        RECT 363.930 17.240 364.250 17.300 ;
        RECT 364.940 17.240 365.080 17.440 ;
        RECT 2577.910 17.380 2578.230 17.440 ;
        RECT 363.930 17.100 365.080 17.240 ;
        RECT 363.930 17.040 364.250 17.100 ;
      LAYER via ;
        RECT 363.960 1407.640 364.220 1407.900 ;
        RECT 393.400 1407.640 393.660 1407.900 ;
        RECT 363.960 17.040 364.220 17.300 ;
        RECT 2577.940 17.380 2578.200 17.640 ;
      LAYER met2 ;
        RECT 363.960 1407.610 364.220 1407.930 ;
        RECT 393.390 1407.755 393.670 1408.125 ;
        RECT 393.400 1407.610 393.660 1407.755 ;
        RECT 364.020 17.330 364.160 1407.610 ;
        RECT 2577.940 17.350 2578.200 17.670 ;
        RECT 363.960 17.010 364.220 17.330 ;
        RECT 2578.000 2.400 2578.140 17.350 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
      LAYER via2 ;
        RECT 393.390 1407.800 393.670 1408.080 ;
      LAYER met3 ;
        RECT 393.365 1408.090 393.695 1408.105 ;
        RECT 410.000 1408.090 414.000 1408.240 ;
        RECT 393.365 1407.790 414.000 1408.090 ;
        RECT 393.365 1407.775 393.695 1407.790 ;
        RECT 410.000 1407.640 414.000 1407.790 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 343.230 2297.960 343.550 2298.020 ;
        RECT 393.370 2297.960 393.690 2298.020 ;
        RECT 343.230 2297.820 393.690 2297.960 ;
        RECT 343.230 2297.760 343.550 2297.820 ;
        RECT 393.370 2297.760 393.690 2297.820 ;
        RECT 343.230 19.620 343.550 19.680 ;
        RECT 811.510 19.620 811.830 19.680 ;
        RECT 343.230 19.480 811.830 19.620 ;
        RECT 343.230 19.420 343.550 19.480 ;
        RECT 811.510 19.420 811.830 19.480 ;
      LAYER via ;
        RECT 343.260 2297.760 343.520 2298.020 ;
        RECT 393.400 2297.760 393.660 2298.020 ;
        RECT 343.260 19.420 343.520 19.680 ;
        RECT 811.540 19.420 811.800 19.680 ;
      LAYER met2 ;
        RECT 393.390 2302.635 393.670 2303.005 ;
        RECT 393.460 2298.050 393.600 2302.635 ;
        RECT 343.260 2297.730 343.520 2298.050 ;
        RECT 393.400 2297.730 393.660 2298.050 ;
        RECT 343.320 19.710 343.460 2297.730 ;
        RECT 343.260 19.390 343.520 19.710 ;
        RECT 811.540 19.390 811.800 19.710 ;
        RECT 811.600 2.400 811.740 19.390 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 393.390 2302.680 393.670 2302.960 ;
      LAYER met3 ;
        RECT 393.365 2302.970 393.695 2302.985 ;
        RECT 410.000 2302.970 414.000 2303.120 ;
        RECT 393.365 2302.670 414.000 2302.970 ;
        RECT 393.365 2302.655 393.695 2302.670 ;
        RECT 410.000 2302.520 414.000 2302.670 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 449.490 500.720 449.810 500.780 ;
        RECT 455.010 500.720 455.330 500.780 ;
        RECT 449.490 500.580 455.330 500.720 ;
        RECT 449.490 500.520 449.810 500.580 ;
        RECT 455.010 500.520 455.330 500.580 ;
        RECT 455.010 86.260 455.330 86.320 ;
        RECT 2594.930 86.260 2595.250 86.320 ;
        RECT 455.010 86.120 2595.250 86.260 ;
        RECT 455.010 86.060 455.330 86.120 ;
        RECT 2594.930 86.060 2595.250 86.120 ;
      LAYER via ;
        RECT 449.520 500.520 449.780 500.780 ;
        RECT 455.040 500.520 455.300 500.780 ;
        RECT 455.040 86.060 455.300 86.320 ;
        RECT 2594.960 86.060 2595.220 86.320 ;
      LAYER met2 ;
        RECT 449.650 510.340 449.930 514.000 ;
        RECT 449.580 510.000 449.930 510.340 ;
        RECT 449.580 500.810 449.720 510.000 ;
        RECT 449.520 500.490 449.780 500.810 ;
        RECT 455.040 500.490 455.300 500.810 ;
        RECT 455.100 86.350 455.240 500.490 ;
        RECT 455.040 86.030 455.300 86.350 ;
        RECT 2594.960 86.030 2595.220 86.350 ;
        RECT 2595.020 7.890 2595.160 86.030 ;
        RECT 2595.020 7.750 2595.620 7.890 ;
        RECT 2595.480 2.400 2595.620 7.750 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 365.385 17.085 365.555 18.615 ;
      LAYER mcon ;
        RECT 365.385 18.445 365.555 18.615 ;
      LAYER met1 ;
        RECT 334.950 1387.100 335.270 1387.160 ;
        RECT 393.370 1387.100 393.690 1387.160 ;
        RECT 334.950 1386.960 393.690 1387.100 ;
        RECT 334.950 1386.900 335.270 1386.960 ;
        RECT 393.370 1386.900 393.690 1386.960 ;
        RECT 334.950 18.600 335.270 18.660 ;
        RECT 365.325 18.600 365.615 18.645 ;
        RECT 334.950 18.460 365.615 18.600 ;
        RECT 334.950 18.400 335.270 18.460 ;
        RECT 365.325 18.415 365.615 18.460 ;
        RECT 365.325 17.240 365.615 17.285 ;
        RECT 2613.330 17.240 2613.650 17.300 ;
        RECT 365.325 17.100 2613.650 17.240 ;
        RECT 365.325 17.055 365.615 17.100 ;
        RECT 2613.330 17.040 2613.650 17.100 ;
      LAYER via ;
        RECT 334.980 1386.900 335.240 1387.160 ;
        RECT 393.400 1386.900 393.660 1387.160 ;
        RECT 334.980 18.400 335.240 18.660 ;
        RECT 2613.360 17.040 2613.620 17.300 ;
      LAYER met2 ;
        RECT 393.390 1390.075 393.670 1390.445 ;
        RECT 393.460 1387.190 393.600 1390.075 ;
        RECT 334.980 1386.870 335.240 1387.190 ;
        RECT 393.400 1386.870 393.660 1387.190 ;
        RECT 335.040 18.690 335.180 1386.870 ;
        RECT 334.980 18.370 335.240 18.690 ;
        RECT 2613.360 17.010 2613.620 17.330 ;
        RECT 2613.420 2.400 2613.560 17.010 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
      LAYER via2 ;
        RECT 393.390 1390.120 393.670 1390.400 ;
      LAYER met3 ;
        RECT 393.365 1390.410 393.695 1390.425 ;
        RECT 410.000 1390.410 414.000 1390.560 ;
        RECT 393.365 1390.110 414.000 1390.410 ;
        RECT 393.365 1390.095 393.695 1390.110 ;
        RECT 410.000 1389.960 414.000 1390.110 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.110 79.460 2242.430 79.520 ;
        RECT 2628.970 79.460 2629.290 79.520 ;
        RECT 2242.110 79.320 2629.290 79.460 ;
        RECT 2242.110 79.260 2242.430 79.320 ;
        RECT 2628.970 79.260 2629.290 79.320 ;
      LAYER via ;
        RECT 2242.140 79.260 2242.400 79.520 ;
        RECT 2629.000 79.260 2629.260 79.520 ;
      LAYER met2 ;
        RECT 2240.890 510.410 2241.170 514.000 ;
        RECT 2240.890 510.270 2242.340 510.410 ;
        RECT 2240.890 510.000 2241.170 510.270 ;
        RECT 2242.200 79.550 2242.340 510.270 ;
        RECT 2242.140 79.230 2242.400 79.550 ;
        RECT 2629.000 79.230 2629.260 79.550 ;
        RECT 2629.060 16.730 2629.200 79.230 ;
        RECT 2629.060 16.590 2631.500 16.730 ;
        RECT 2631.360 2.400 2631.500 16.590 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2366.310 431.360 2366.630 431.420 ;
        RECT 2642.770 431.360 2643.090 431.420 ;
        RECT 2366.310 431.220 2643.090 431.360 ;
        RECT 2366.310 431.160 2366.630 431.220 ;
        RECT 2642.770 431.160 2643.090 431.220 ;
        RECT 2642.770 17.240 2643.090 17.300 ;
        RECT 2649.210 17.240 2649.530 17.300 ;
        RECT 2642.770 17.100 2649.530 17.240 ;
        RECT 2642.770 17.040 2643.090 17.100 ;
        RECT 2649.210 17.040 2649.530 17.100 ;
      LAYER via ;
        RECT 2366.340 431.160 2366.600 431.420 ;
        RECT 2642.800 431.160 2643.060 431.420 ;
        RECT 2642.800 17.040 2643.060 17.300 ;
        RECT 2649.240 17.040 2649.500 17.300 ;
      LAYER met2 ;
        RECT 2364.170 510.410 2364.450 514.000 ;
        RECT 2364.170 510.270 2366.540 510.410 ;
        RECT 2364.170 510.000 2364.450 510.270 ;
        RECT 2366.400 431.450 2366.540 510.270 ;
        RECT 2366.340 431.130 2366.600 431.450 ;
        RECT 2642.800 431.130 2643.060 431.450 ;
        RECT 2642.860 17.330 2643.000 431.130 ;
        RECT 2642.800 17.010 2643.060 17.330 ;
        RECT 2649.240 17.010 2649.500 17.330 ;
        RECT 2649.300 2.400 2649.440 17.010 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1088.045 3002.285 1088.215 3006.535 ;
      LAYER mcon ;
        RECT 1088.045 3006.365 1088.215 3006.535 ;
      LAYER met1 ;
        RECT 1087.970 3006.520 1088.290 3006.580 ;
        RECT 1087.775 3006.380 1088.290 3006.520 ;
        RECT 1087.970 3006.320 1088.290 3006.380 ;
        RECT 1087.985 3002.440 1088.275 3002.485 ;
        RECT 2663.470 3002.440 2663.790 3002.500 ;
        RECT 1087.985 3002.300 2663.790 3002.440 ;
        RECT 1087.985 3002.255 1088.275 3002.300 ;
        RECT 2663.470 3002.240 2663.790 3002.300 ;
      LAYER via ;
        RECT 1088.000 3006.320 1088.260 3006.580 ;
        RECT 2663.500 3002.240 2663.760 3002.500 ;
      LAYER met2 ;
        RECT 1086.290 3006.690 1086.570 3010.000 ;
        RECT 1086.290 3006.610 1088.200 3006.690 ;
        RECT 1086.290 3006.550 1088.260 3006.610 ;
        RECT 1086.290 3006.000 1086.570 3006.550 ;
        RECT 1088.000 3006.290 1088.260 3006.550 ;
        RECT 2663.500 3002.210 2663.760 3002.530 ;
        RECT 2663.560 17.410 2663.700 3002.210 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.650 30.755 2684.930 31.125 ;
        RECT 2684.720 2.400 2684.860 30.755 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
      LAYER via2 ;
        RECT 2684.650 30.800 2684.930 31.080 ;
      LAYER met3 ;
        RECT 410.000 1444.360 414.000 1444.960 ;
        RECT 349.870 1442.770 350.250 1442.780 ;
        RECT 410.630 1442.770 410.930 1444.360 ;
        RECT 349.870 1442.470 410.930 1442.770 ;
        RECT 349.870 1442.460 350.250 1442.470 ;
        RECT 349.870 31.090 350.250 31.100 ;
        RECT 2684.625 31.090 2684.955 31.105 ;
        RECT 349.870 30.790 2684.955 31.090 ;
        RECT 349.870 30.780 350.250 30.790 ;
        RECT 2684.625 30.775 2684.955 30.790 ;
      LAYER via3 ;
        RECT 349.900 1442.460 350.220 1442.780 ;
        RECT 349.900 30.780 350.220 31.100 ;
      LAYER met4 ;
        RECT 349.895 1442.455 350.225 1442.785 ;
        RECT 349.910 31.105 350.210 1442.455 ;
        RECT 349.895 30.775 350.225 31.105 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 757.765 386.665 757.935 405.535 ;
        RECT 757.305 338.045 757.475 385.815 ;
        RECT 757.765 193.205 757.935 241.315 ;
      LAYER mcon ;
        RECT 757.765 405.365 757.935 405.535 ;
        RECT 757.305 385.645 757.475 385.815 ;
        RECT 757.765 241.145 757.935 241.315 ;
      LAYER met1 ;
        RECT 757.690 435.100 758.010 435.160 ;
        RECT 758.150 435.100 758.470 435.160 ;
        RECT 757.690 434.960 758.470 435.100 ;
        RECT 757.690 434.900 758.010 434.960 ;
        RECT 758.150 434.900 758.470 434.960 ;
        RECT 757.690 405.520 758.010 405.580 ;
        RECT 757.495 405.380 758.010 405.520 ;
        RECT 757.690 405.320 758.010 405.380 ;
        RECT 757.690 386.820 758.010 386.880 ;
        RECT 757.495 386.680 758.010 386.820 ;
        RECT 757.690 386.620 758.010 386.680 ;
        RECT 757.230 385.800 757.550 385.860 ;
        RECT 757.035 385.660 757.550 385.800 ;
        RECT 757.230 385.600 757.550 385.660 ;
        RECT 757.245 338.200 757.535 338.245 ;
        RECT 757.690 338.200 758.010 338.260 ;
        RECT 757.245 338.060 758.010 338.200 ;
        RECT 757.245 338.015 757.535 338.060 ;
        RECT 757.690 338.000 758.010 338.060 ;
        RECT 757.690 304.200 758.010 304.260 ;
        RECT 757.320 304.060 758.010 304.200 ;
        RECT 757.320 303.580 757.460 304.060 ;
        RECT 757.690 304.000 758.010 304.060 ;
        RECT 757.230 303.320 757.550 303.580 ;
        RECT 757.230 255.240 757.550 255.300 ;
        RECT 758.150 255.240 758.470 255.300 ;
        RECT 757.230 255.100 758.470 255.240 ;
        RECT 757.230 255.040 757.550 255.100 ;
        RECT 758.150 255.040 758.470 255.100 ;
        RECT 757.705 241.300 757.995 241.345 ;
        RECT 758.150 241.300 758.470 241.360 ;
        RECT 757.705 241.160 758.470 241.300 ;
        RECT 757.705 241.115 757.995 241.160 ;
        RECT 758.150 241.100 758.470 241.160 ;
        RECT 757.690 193.360 758.010 193.420 ;
        RECT 757.495 193.220 758.010 193.360 ;
        RECT 757.690 193.160 758.010 193.220 ;
        RECT 757.230 134.540 757.550 134.600 ;
        RECT 2697.970 134.540 2698.290 134.600 ;
        RECT 757.230 134.400 2698.290 134.540 ;
        RECT 757.230 134.340 757.550 134.400 ;
        RECT 2697.970 134.340 2698.290 134.400 ;
      LAYER via ;
        RECT 757.720 434.900 757.980 435.160 ;
        RECT 758.180 434.900 758.440 435.160 ;
        RECT 757.720 405.320 757.980 405.580 ;
        RECT 757.720 386.620 757.980 386.880 ;
        RECT 757.260 385.600 757.520 385.860 ;
        RECT 757.720 338.000 757.980 338.260 ;
        RECT 757.720 304.000 757.980 304.260 ;
        RECT 757.260 303.320 757.520 303.580 ;
        RECT 757.260 255.040 757.520 255.300 ;
        RECT 758.180 255.040 758.440 255.300 ;
        RECT 758.180 241.100 758.440 241.360 ;
        RECT 757.720 193.160 757.980 193.420 ;
        RECT 757.260 134.340 757.520 134.600 ;
        RECT 2698.000 134.340 2698.260 134.600 ;
      LAYER met2 ;
        RECT 757.850 511.090 758.130 514.000 ;
        RECT 757.850 510.950 758.840 511.090 ;
        RECT 757.850 510.000 758.130 510.950 ;
        RECT 758.700 483.210 758.840 510.950 ;
        RECT 758.240 483.070 758.840 483.210 ;
        RECT 758.240 435.190 758.380 483.070 ;
        RECT 757.720 434.870 757.980 435.190 ;
        RECT 758.180 434.870 758.440 435.190 ;
        RECT 757.780 405.610 757.920 434.870 ;
        RECT 757.720 405.290 757.980 405.610 ;
        RECT 757.720 386.650 757.980 386.910 ;
        RECT 757.320 386.590 757.980 386.650 ;
        RECT 757.320 386.510 757.920 386.590 ;
        RECT 757.320 385.890 757.460 386.510 ;
        RECT 757.260 385.570 757.520 385.890 ;
        RECT 757.720 337.970 757.980 338.290 ;
        RECT 757.780 304.290 757.920 337.970 ;
        RECT 757.720 303.970 757.980 304.290 ;
        RECT 757.260 303.290 757.520 303.610 ;
        RECT 757.320 255.330 757.460 303.290 ;
        RECT 757.260 255.010 757.520 255.330 ;
        RECT 758.180 255.010 758.440 255.330 ;
        RECT 758.240 241.390 758.380 255.010 ;
        RECT 758.180 241.070 758.440 241.390 ;
        RECT 757.720 193.130 757.980 193.450 ;
        RECT 757.780 158.850 757.920 193.130 ;
        RECT 757.320 158.710 757.920 158.850 ;
        RECT 757.320 134.630 757.460 158.710 ;
        RECT 757.260 134.310 757.520 134.630 ;
        RECT 2698.000 134.310 2698.260 134.630 ;
        RECT 2698.060 17.410 2698.200 134.310 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2032.885 3004.665 2033.055 3015.715 ;
      LAYER mcon ;
        RECT 2032.885 3015.545 2033.055 3015.715 ;
      LAYER met1 ;
        RECT 1975.770 3015.700 1976.090 3015.760 ;
        RECT 2032.825 3015.700 2033.115 3015.745 ;
        RECT 1975.770 3015.560 2033.115 3015.700 ;
        RECT 1975.770 3015.500 1976.090 3015.560 ;
        RECT 2032.825 3015.515 2033.115 3015.560 ;
        RECT 2032.825 3004.820 2033.115 3004.865 ;
        RECT 2718.670 3004.820 2718.990 3004.880 ;
        RECT 2032.825 3004.680 2718.990 3004.820 ;
        RECT 2032.825 3004.635 2033.115 3004.680 ;
        RECT 2718.670 3004.620 2718.990 3004.680 ;
      LAYER via ;
        RECT 1975.800 3015.500 1976.060 3015.760 ;
        RECT 2718.700 3004.620 2718.960 3004.880 ;
      LAYER met2 ;
        RECT 1975.800 3015.470 1976.060 3015.790 ;
        RECT 1975.860 3010.000 1976.000 3015.470 ;
        RECT 1975.860 3009.340 1976.210 3010.000 ;
        RECT 1975.930 3006.000 1976.210 3009.340 ;
        RECT 2718.700 3004.590 2718.960 3004.910 ;
        RECT 2718.760 17.410 2718.900 3004.590 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 93.740 1821.530 93.800 ;
        RECT 2732.930 93.740 2733.250 93.800 ;
        RECT 1821.210 93.600 2733.250 93.740 ;
        RECT 1821.210 93.540 1821.530 93.600 ;
        RECT 2732.930 93.540 2733.250 93.600 ;
      LAYER via ;
        RECT 1821.240 93.540 1821.500 93.800 ;
        RECT 2732.960 93.540 2733.220 93.800 ;
      LAYER met2 ;
        RECT 1820.450 510.410 1820.730 514.000 ;
        RECT 1820.450 510.270 1821.440 510.410 ;
        RECT 1820.450 510.000 1820.730 510.270 ;
        RECT 1821.300 93.830 1821.440 510.270 ;
        RECT 1821.240 93.510 1821.500 93.830 ;
        RECT 2732.960 93.510 2733.220 93.830 ;
        RECT 2733.020 17.410 2733.160 93.510 ;
        RECT 2733.020 17.270 2738.680 17.410 ;
        RECT 2738.540 2.400 2738.680 17.270 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 127.740 551.930 127.800 ;
        RECT 2753.170 127.740 2753.490 127.800 ;
        RECT 551.610 127.600 2753.490 127.740 ;
        RECT 551.610 127.540 551.930 127.600 ;
        RECT 2753.170 127.540 2753.490 127.600 ;
      LAYER via ;
        RECT 551.640 127.540 551.900 127.800 ;
        RECT 2753.200 127.540 2753.460 127.800 ;
      LAYER met2 ;
        RECT 548.090 510.410 548.370 514.000 ;
        RECT 548.090 510.270 551.840 510.410 ;
        RECT 548.090 510.000 548.370 510.270 ;
        RECT 551.700 127.830 551.840 510.270 ;
        RECT 551.640 127.510 551.900 127.830 ;
        RECT 2753.200 127.510 2753.460 127.830 ;
        RECT 2753.260 17.410 2753.400 127.510 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.450 2994.960 323.770 2995.020 ;
        RECT 393.370 2994.960 393.690 2995.020 ;
        RECT 323.450 2994.820 393.690 2994.960 ;
        RECT 323.450 2994.760 323.770 2994.820 ;
        RECT 393.370 2994.760 393.690 2994.820 ;
        RECT 323.450 19.280 323.770 19.340 ;
        RECT 829.450 19.280 829.770 19.340 ;
        RECT 323.450 19.140 829.770 19.280 ;
        RECT 323.450 19.080 323.770 19.140 ;
        RECT 829.450 19.080 829.770 19.140 ;
      LAYER via ;
        RECT 323.480 2994.760 323.740 2995.020 ;
        RECT 393.400 2994.760 393.660 2995.020 ;
        RECT 323.480 19.080 323.740 19.340 ;
        RECT 829.480 19.080 829.740 19.340 ;
      LAYER met2 ;
        RECT 393.390 2997.595 393.670 2997.965 ;
        RECT 393.460 2995.050 393.600 2997.595 ;
        RECT 323.480 2994.730 323.740 2995.050 ;
        RECT 393.400 2994.730 393.660 2995.050 ;
        RECT 323.540 19.370 323.680 2994.730 ;
        RECT 323.480 19.050 323.740 19.370 ;
        RECT 829.480 19.050 829.740 19.370 ;
        RECT 829.540 2.400 829.680 19.050 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 393.390 2997.640 393.670 2997.920 ;
      LAYER met3 ;
        RECT 393.365 2997.930 393.695 2997.945 ;
        RECT 410.000 2997.930 414.000 2998.080 ;
        RECT 393.365 2997.630 414.000 2997.930 ;
        RECT 393.365 2997.615 393.695 2997.630 ;
        RECT 410.000 2997.480 414.000 2997.630 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 369.910 1207.580 370.230 1207.640 ;
        RECT 393.370 1207.580 393.690 1207.640 ;
        RECT 369.910 1207.440 393.690 1207.580 ;
        RECT 369.910 1207.380 370.230 1207.440 ;
        RECT 393.370 1207.380 393.690 1207.440 ;
        RECT 369.910 31.860 370.230 31.920 ;
        RECT 2774.330 31.860 2774.650 31.920 ;
        RECT 369.910 31.720 2774.650 31.860 ;
        RECT 369.910 31.660 370.230 31.720 ;
        RECT 2774.330 31.660 2774.650 31.720 ;
      LAYER via ;
        RECT 369.940 1207.380 370.200 1207.640 ;
        RECT 393.400 1207.380 393.660 1207.640 ;
        RECT 369.940 31.660 370.200 31.920 ;
        RECT 2774.360 31.660 2774.620 31.920 ;
      LAYER met2 ;
        RECT 393.390 1207.835 393.670 1208.205 ;
        RECT 393.460 1207.670 393.600 1207.835 ;
        RECT 369.940 1207.350 370.200 1207.670 ;
        RECT 393.400 1207.350 393.660 1207.670 ;
        RECT 370.000 31.950 370.140 1207.350 ;
        RECT 369.940 31.630 370.200 31.950 ;
        RECT 2774.360 31.630 2774.620 31.950 ;
        RECT 2774.420 16.730 2774.560 31.630 ;
        RECT 2773.960 16.590 2774.560 16.730 ;
        RECT 2773.960 2.400 2774.100 16.590 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
      LAYER via2 ;
        RECT 393.390 1207.880 393.670 1208.160 ;
      LAYER met3 ;
        RECT 393.365 1208.170 393.695 1208.185 ;
        RECT 410.000 1208.170 414.000 1208.320 ;
        RECT 393.365 1207.870 414.000 1208.170 ;
        RECT 393.365 1207.855 393.695 1207.870 ;
        RECT 410.000 1207.720 414.000 1207.870 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 330.350 2518.620 330.670 2518.680 ;
        RECT 393.370 2518.620 393.690 2518.680 ;
        RECT 330.350 2518.480 393.690 2518.620 ;
        RECT 330.350 2518.420 330.670 2518.480 ;
        RECT 393.370 2518.420 393.690 2518.480 ;
        RECT 330.350 31.520 330.670 31.580 ;
        RECT 2791.810 31.520 2792.130 31.580 ;
        RECT 330.350 31.380 2792.130 31.520 ;
        RECT 330.350 31.320 330.670 31.380 ;
        RECT 2791.810 31.320 2792.130 31.380 ;
      LAYER via ;
        RECT 330.380 2518.420 330.640 2518.680 ;
        RECT 393.400 2518.420 393.660 2518.680 ;
        RECT 330.380 31.320 330.640 31.580 ;
        RECT 2791.840 31.320 2792.100 31.580 ;
      LAYER met2 ;
        RECT 393.390 2522.955 393.670 2523.325 ;
        RECT 393.460 2518.710 393.600 2522.955 ;
        RECT 330.380 2518.390 330.640 2518.710 ;
        RECT 393.400 2518.390 393.660 2518.710 ;
        RECT 330.440 31.610 330.580 2518.390 ;
        RECT 330.380 31.290 330.640 31.610 ;
        RECT 2791.840 31.290 2792.100 31.610 ;
        RECT 2791.900 2.400 2792.040 31.290 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 393.390 2523.000 393.670 2523.280 ;
      LAYER met3 ;
        RECT 393.365 2523.290 393.695 2523.305 ;
        RECT 410.000 2523.290 414.000 2523.440 ;
        RECT 393.365 2522.990 414.000 2523.290 ;
        RECT 393.365 2522.975 393.695 2522.990 ;
        RECT 410.000 2522.840 414.000 2522.990 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 2429.200 330.210 2429.260 ;
        RECT 393.370 2429.200 393.690 2429.260 ;
        RECT 329.890 2429.060 393.690 2429.200 ;
        RECT 329.890 2429.000 330.210 2429.060 ;
        RECT 393.370 2429.000 393.690 2429.060 ;
        RECT 329.890 31.180 330.210 31.240 ;
        RECT 2809.750 31.180 2810.070 31.240 ;
        RECT 329.890 31.040 2810.070 31.180 ;
        RECT 329.890 30.980 330.210 31.040 ;
        RECT 2809.750 30.980 2810.070 31.040 ;
      LAYER via ;
        RECT 329.920 2429.000 330.180 2429.260 ;
        RECT 393.400 2429.000 393.660 2429.260 ;
        RECT 329.920 30.980 330.180 31.240 ;
        RECT 2809.780 30.980 2810.040 31.240 ;
      LAYER met2 ;
        RECT 393.390 2430.475 393.670 2430.845 ;
        RECT 393.460 2429.290 393.600 2430.475 ;
        RECT 329.920 2428.970 330.180 2429.290 ;
        RECT 393.400 2428.970 393.660 2429.290 ;
        RECT 329.980 31.270 330.120 2428.970 ;
        RECT 329.920 30.950 330.180 31.270 ;
        RECT 2809.780 30.950 2810.040 31.270 ;
        RECT 2809.840 2.400 2809.980 30.950 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
      LAYER via2 ;
        RECT 393.390 2430.520 393.670 2430.800 ;
      LAYER met3 ;
        RECT 393.365 2430.810 393.695 2430.825 ;
        RECT 410.000 2430.810 414.000 2430.960 ;
        RECT 393.365 2430.510 414.000 2430.810 ;
        RECT 393.365 2430.495 393.695 2430.510 ;
        RECT 410.000 2430.360 414.000 2430.510 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1580.220 2520.730 1580.280 ;
        RECT 2790.890 1580.220 2791.210 1580.280 ;
        RECT 2520.410 1580.080 2791.210 1580.220 ;
        RECT 2520.410 1580.020 2520.730 1580.080 ;
        RECT 2790.890 1580.020 2791.210 1580.080 ;
        RECT 2790.890 427.620 2791.210 427.680 ;
        RECT 2822.170 427.620 2822.490 427.680 ;
        RECT 2790.890 427.480 2822.490 427.620 ;
        RECT 2790.890 427.420 2791.210 427.480 ;
        RECT 2822.170 427.420 2822.490 427.480 ;
      LAYER via ;
        RECT 2520.440 1580.020 2520.700 1580.280 ;
        RECT 2790.920 1580.020 2791.180 1580.280 ;
        RECT 2790.920 427.420 2791.180 427.680 ;
        RECT 2822.200 427.420 2822.460 427.680 ;
      LAYER met2 ;
        RECT 2520.430 1580.475 2520.710 1580.845 ;
        RECT 2520.500 1580.310 2520.640 1580.475 ;
        RECT 2520.440 1579.990 2520.700 1580.310 ;
        RECT 2790.920 1579.990 2791.180 1580.310 ;
        RECT 2790.980 427.710 2791.120 1579.990 ;
        RECT 2790.920 427.390 2791.180 427.710 ;
        RECT 2822.200 427.390 2822.460 427.710 ;
        RECT 2822.260 17.410 2822.400 427.390 ;
        RECT 2822.260 17.270 2827.920 17.410 ;
        RECT 2827.780 2.400 2827.920 17.270 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1580.520 2520.710 1580.800 ;
      LAYER met3 ;
        RECT 2506.000 1580.810 2510.000 1580.960 ;
        RECT 2520.405 1580.810 2520.735 1580.825 ;
        RECT 2506.000 1580.510 2520.735 1580.810 ;
        RECT 2506.000 1580.360 2510.000 1580.510 ;
        RECT 2520.405 1580.495 2520.735 1580.510 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 334.490 1256.540 334.810 1256.600 ;
        RECT 393.370 1256.540 393.690 1256.600 ;
        RECT 334.490 1256.400 393.690 1256.540 ;
        RECT 334.490 1256.340 334.810 1256.400 ;
        RECT 393.370 1256.340 393.690 1256.400 ;
        RECT 334.490 30.840 334.810 30.900 ;
        RECT 2845.170 30.840 2845.490 30.900 ;
        RECT 334.490 30.700 2845.490 30.840 ;
        RECT 334.490 30.640 334.810 30.700 ;
        RECT 2845.170 30.640 2845.490 30.700 ;
      LAYER via ;
        RECT 334.520 1256.340 334.780 1256.600 ;
        RECT 393.400 1256.340 393.660 1256.600 ;
        RECT 334.520 30.640 334.780 30.900 ;
        RECT 2845.200 30.640 2845.460 30.900 ;
      LAYER met2 ;
        RECT 393.390 1262.235 393.670 1262.605 ;
        RECT 393.460 1256.630 393.600 1262.235 ;
        RECT 334.520 1256.310 334.780 1256.630 ;
        RECT 393.400 1256.310 393.660 1256.630 ;
        RECT 334.580 30.930 334.720 1256.310 ;
        RECT 334.520 30.610 334.780 30.930 ;
        RECT 2845.200 30.610 2845.460 30.930 ;
        RECT 2845.260 2.400 2845.400 30.610 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 393.390 1262.280 393.670 1262.560 ;
      LAYER met3 ;
        RECT 393.365 1262.570 393.695 1262.585 ;
        RECT 410.000 1262.570 414.000 1262.720 ;
        RECT 393.365 1262.270 414.000 1262.570 ;
        RECT 393.365 1262.255 393.695 1262.270 ;
        RECT 410.000 1262.120 414.000 1262.270 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2516.730 538.460 2517.050 538.520 ;
        RECT 2659.790 538.460 2660.110 538.520 ;
        RECT 2516.730 538.320 2660.110 538.460 ;
        RECT 2516.730 538.260 2517.050 538.320 ;
        RECT 2659.790 538.260 2660.110 538.320 ;
        RECT 2659.790 32.200 2660.110 32.260 ;
        RECT 2863.110 32.200 2863.430 32.260 ;
        RECT 2659.790 32.060 2863.430 32.200 ;
        RECT 2659.790 32.000 2660.110 32.060 ;
        RECT 2863.110 32.000 2863.430 32.060 ;
      LAYER via ;
        RECT 2516.760 538.260 2517.020 538.520 ;
        RECT 2659.820 538.260 2660.080 538.520 ;
        RECT 2659.820 32.000 2660.080 32.260 ;
        RECT 2863.140 32.000 2863.400 32.260 ;
      LAYER met2 ;
        RECT 2516.750 540.075 2517.030 540.445 ;
        RECT 2516.820 538.550 2516.960 540.075 ;
        RECT 2516.760 538.230 2517.020 538.550 ;
        RECT 2659.820 538.230 2660.080 538.550 ;
        RECT 2659.880 32.290 2660.020 538.230 ;
        RECT 2659.820 31.970 2660.080 32.290 ;
        RECT 2863.140 31.970 2863.400 32.290 ;
        RECT 2863.200 2.400 2863.340 31.970 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
      LAYER via2 ;
        RECT 2516.750 540.120 2517.030 540.400 ;
      LAYER met3 ;
        RECT 2506.000 540.410 2510.000 540.560 ;
        RECT 2516.725 540.410 2517.055 540.425 ;
        RECT 2506.000 540.110 2517.055 540.410 ;
        RECT 2506.000 539.960 2510.000 540.110 ;
        RECT 2516.725 540.095 2517.055 540.110 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2436.000 2519.810 2436.060 ;
        RECT 2859.890 2436.000 2860.210 2436.060 ;
        RECT 2519.490 2435.860 2860.210 2436.000 ;
        RECT 2519.490 2435.800 2519.810 2435.860 ;
        RECT 2859.890 2435.800 2860.210 2435.860 ;
        RECT 2859.890 27.780 2860.210 27.840 ;
        RECT 2881.050 27.780 2881.370 27.840 ;
        RECT 2859.890 27.640 2881.370 27.780 ;
        RECT 2859.890 27.580 2860.210 27.640 ;
        RECT 2881.050 27.580 2881.370 27.640 ;
      LAYER via ;
        RECT 2519.520 2435.800 2519.780 2436.060 ;
        RECT 2859.920 2435.800 2860.180 2436.060 ;
        RECT 2859.920 27.580 2860.180 27.840 ;
        RECT 2881.080 27.580 2881.340 27.840 ;
      LAYER met2 ;
        RECT 2519.510 2438.635 2519.790 2439.005 ;
        RECT 2519.580 2436.090 2519.720 2438.635 ;
        RECT 2519.520 2435.770 2519.780 2436.090 ;
        RECT 2859.920 2435.770 2860.180 2436.090 ;
        RECT 2859.980 27.870 2860.120 2435.770 ;
        RECT 2859.920 27.550 2860.180 27.870 ;
        RECT 2881.080 27.550 2881.340 27.870 ;
        RECT 2881.140 2.400 2881.280 27.550 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2438.680 2519.790 2438.960 ;
      LAYER met3 ;
        RECT 2506.000 2438.970 2510.000 2439.120 ;
        RECT 2519.485 2438.970 2519.815 2438.985 ;
        RECT 2506.000 2438.670 2519.815 2438.970 ;
        RECT 2506.000 2438.520 2510.000 2438.670 ;
        RECT 2519.485 2438.655 2519.815 2438.670 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 3029.980 841.730 3030.040 ;
        RECT 2866.790 3029.980 2867.110 3030.040 ;
        RECT 841.410 3029.840 2867.110 3029.980 ;
        RECT 841.410 3029.780 841.730 3029.840 ;
        RECT 2866.790 3029.780 2867.110 3029.840 ;
        RECT 2866.790 17.240 2867.110 17.300 ;
        RECT 2898.990 17.240 2899.310 17.300 ;
        RECT 2866.790 17.100 2899.310 17.240 ;
        RECT 2866.790 17.040 2867.110 17.100 ;
        RECT 2898.990 17.040 2899.310 17.100 ;
      LAYER via ;
        RECT 841.440 3029.780 841.700 3030.040 ;
        RECT 2866.820 3029.780 2867.080 3030.040 ;
        RECT 2866.820 17.040 2867.080 17.300 ;
        RECT 2899.020 17.040 2899.280 17.300 ;
      LAYER met2 ;
        RECT 841.440 3029.925 841.700 3030.070 ;
        RECT 468.830 3029.555 469.110 3029.925 ;
        RECT 841.430 3029.555 841.710 3029.925 ;
        RECT 2866.820 3029.750 2867.080 3030.070 ;
        RECT 468.900 3010.000 469.040 3029.555 ;
        RECT 468.900 3009.340 469.250 3010.000 ;
        RECT 468.970 3006.000 469.250 3009.340 ;
        RECT 2866.880 17.330 2867.020 3029.750 ;
        RECT 2866.820 17.010 2867.080 17.330 ;
        RECT 2899.020 17.010 2899.280 17.330 ;
        RECT 2899.080 2.400 2899.220 17.010 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 468.830 3029.600 469.110 3029.880 ;
        RECT 841.430 3029.600 841.710 3029.880 ;
      LAYER met3 ;
        RECT 468.805 3029.890 469.135 3029.905 ;
        RECT 841.405 3029.890 841.735 3029.905 ;
        RECT 468.805 3029.590 841.735 3029.890 ;
        RECT 468.805 3029.575 469.135 3029.590 ;
        RECT 841.405 3029.575 841.735 3029.590 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.950 19.875 847.230 20.245 ;
        RECT 847.020 2.400 847.160 19.875 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 846.950 19.920 847.230 20.200 ;
      LAYER met3 ;
        RECT 2506.000 2986.600 2510.000 2987.200 ;
        RECT 2508.230 2982.970 2508.530 2986.600 ;
        RECT 2508.230 2982.670 2509.450 2982.970 ;
        RECT 2509.150 2981.610 2509.450 2982.670 ;
        RECT 2567.070 2981.610 2567.450 2981.620 ;
        RECT 2509.150 2981.310 2567.450 2981.610 ;
        RECT 2567.070 2981.300 2567.450 2981.310 ;
        RECT 1207.310 508.450 1207.690 508.460 ;
        RECT 1255.150 508.450 1255.530 508.460 ;
        RECT 1207.310 508.150 1255.530 508.450 ;
        RECT 1207.310 508.140 1207.690 508.150 ;
        RECT 1255.150 508.140 1255.530 508.150 ;
        RECT 1979.190 505.050 1979.570 505.060 ;
        RECT 2014.150 505.050 2014.530 505.060 ;
        RECT 1979.190 504.750 2014.530 505.050 ;
        RECT 1979.190 504.740 1979.570 504.750 ;
        RECT 2014.150 504.740 2014.530 504.750 ;
        RECT 2018.750 505.050 2019.130 505.060 ;
        RECT 2061.990 505.050 2062.370 505.060 ;
        RECT 2018.750 504.750 2062.370 505.050 ;
        RECT 2018.750 504.740 2019.130 504.750 ;
        RECT 2061.990 504.740 2062.370 504.750 ;
        RECT 2407.910 505.050 2408.290 505.060 ;
        RECT 2475.990 505.050 2476.370 505.060 ;
        RECT 2407.910 504.750 2476.370 505.050 ;
        RECT 2407.910 504.740 2408.290 504.750 ;
        RECT 2475.990 504.740 2476.370 504.750 ;
        RECT 2522.910 505.050 2523.290 505.060 ;
        RECT 2535.790 505.050 2536.170 505.060 ;
        RECT 2522.910 504.750 2536.170 505.050 ;
        RECT 2522.910 504.740 2523.290 504.750 ;
        RECT 2535.790 504.740 2536.170 504.750 ;
        RECT 1159.470 501.650 1159.850 501.660 ;
        RECT 1206.390 501.650 1206.770 501.660 ;
        RECT 1159.470 501.350 1206.770 501.650 ;
        RECT 1159.470 501.340 1159.850 501.350 ;
        RECT 1206.390 501.340 1206.770 501.350 ;
        RECT 1352.670 501.650 1353.050 501.660 ;
        RECT 1369.230 501.650 1369.610 501.660 ;
        RECT 1352.670 501.350 1369.610 501.650 ;
        RECT 1352.670 501.340 1353.050 501.350 ;
        RECT 1369.230 501.340 1369.610 501.350 ;
        RECT 1739.070 501.650 1739.450 501.660 ;
        RECT 1755.630 501.650 1756.010 501.660 ;
        RECT 1739.070 501.350 1756.010 501.650 ;
        RECT 1739.070 501.340 1739.450 501.350 ;
        RECT 1755.630 501.340 1756.010 501.350 ;
        RECT 846.925 20.210 847.255 20.225 ;
        RECT 847.590 20.210 847.970 20.220 ;
        RECT 846.925 19.910 847.970 20.210 ;
        RECT 846.925 19.895 847.255 19.910 ;
        RECT 847.590 19.900 847.970 19.910 ;
      LAYER via3 ;
        RECT 2567.100 2981.300 2567.420 2981.620 ;
        RECT 1207.340 508.140 1207.660 508.460 ;
        RECT 1255.180 508.140 1255.500 508.460 ;
        RECT 1979.220 504.740 1979.540 505.060 ;
        RECT 2014.180 504.740 2014.500 505.060 ;
        RECT 2018.780 504.740 2019.100 505.060 ;
        RECT 2062.020 504.740 2062.340 505.060 ;
        RECT 2407.940 504.740 2408.260 505.060 ;
        RECT 2476.020 504.740 2476.340 505.060 ;
        RECT 2522.940 504.740 2523.260 505.060 ;
        RECT 2535.820 504.740 2536.140 505.060 ;
        RECT 1159.500 501.340 1159.820 501.660 ;
        RECT 1206.420 501.340 1206.740 501.660 ;
        RECT 1352.700 501.340 1353.020 501.660 ;
        RECT 1369.260 501.340 1369.580 501.660 ;
        RECT 1739.100 501.340 1739.420 501.660 ;
        RECT 1755.660 501.340 1755.980 501.660 ;
        RECT 847.620 19.900 847.940 20.220 ;
      LAYER met4 ;
        RECT 2567.095 2981.295 2567.425 2981.625 ;
        RECT 847.190 507.710 848.370 508.890 ;
        RECT 1206.910 507.710 1208.090 508.890 ;
        RECT 1255.175 508.135 1255.505 508.465 ;
        RECT 847.630 20.225 847.930 507.710 ;
        RECT 1205.990 504.310 1207.170 505.490 ;
        RECT 1159.070 500.910 1160.250 502.090 ;
        RECT 1206.430 501.665 1206.730 504.310 ;
        RECT 1255.190 502.090 1255.490 508.135 ;
        RECT 2061.590 507.710 2062.770 508.890 ;
        RECT 2475.590 507.710 2476.770 508.890 ;
        RECT 2522.510 507.710 2523.690 508.890 ;
        RECT 1368.830 504.310 1370.010 505.490 ;
        RECT 1755.230 504.310 1756.410 505.490 ;
        RECT 1978.790 504.310 1979.970 505.490 ;
        RECT 2013.750 504.310 2014.930 505.490 ;
        RECT 2018.350 504.310 2019.530 505.490 ;
        RECT 2062.030 505.065 2062.330 507.710 ;
        RECT 2062.015 504.735 2062.345 505.065 ;
        RECT 2407.510 504.310 2408.690 505.490 ;
        RECT 2476.030 505.065 2476.330 507.710 ;
        RECT 2522.950 505.065 2523.250 507.710 ;
        RECT 2567.110 505.490 2567.410 2981.295 ;
        RECT 2476.015 504.735 2476.345 505.065 ;
        RECT 2522.935 504.735 2523.265 505.065 ;
        RECT 2535.390 504.310 2536.570 505.490 ;
        RECT 2566.670 504.310 2567.850 505.490 ;
        RECT 1206.415 501.335 1206.745 501.665 ;
        RECT 1254.750 500.910 1255.930 502.090 ;
        RECT 1352.270 500.910 1353.450 502.090 ;
        RECT 1369.270 501.665 1369.570 504.310 ;
        RECT 1369.255 501.335 1369.585 501.665 ;
        RECT 1738.670 500.910 1739.850 502.090 ;
        RECT 1755.670 501.665 1755.970 504.310 ;
        RECT 1755.655 501.335 1755.985 501.665 ;
        RECT 847.615 19.895 847.945 20.225 ;
      LAYER met5 ;
        RECT 2475.380 509.100 2480.660 509.780 ;
        RECT 846.980 507.500 908.380 509.100 ;
        RECT 906.780 505.700 908.380 507.500 ;
        RECT 931.620 507.500 1026.140 509.100 ;
        RECT 931.620 505.700 933.220 507.500 ;
        RECT 906.780 504.100 933.220 505.700 ;
        RECT 1024.540 502.300 1026.140 507.500 ;
        RECT 1075.140 505.700 1077.660 509.100 ;
        RECT 1206.700 505.700 1208.300 509.100 ;
        RECT 1075.140 504.100 1124.580 505.700 ;
        RECT 1205.780 504.100 1208.300 505.700 ;
        RECT 1268.340 505.700 1270.860 509.100 ;
        RECT 1434.860 507.500 1484.300 509.100 ;
        RECT 1434.860 505.700 1436.460 507.500 ;
        RECT 1268.340 504.100 1317.780 505.700 ;
        RECT 1368.620 504.100 1436.460 505.700 ;
        RECT 1075.140 502.300 1076.740 504.100 ;
        RECT 1024.540 500.700 1076.740 502.300 ;
        RECT 1122.980 502.300 1124.580 504.100 ;
        RECT 1268.340 502.300 1269.940 504.100 ;
        RECT 1122.980 500.700 1160.460 502.300 ;
        RECT 1254.540 500.700 1269.940 502.300 ;
        RECT 1316.180 502.300 1317.780 504.100 ;
        RECT 1482.700 502.300 1484.300 507.500 ;
        RECT 1558.140 507.500 1581.820 509.100 ;
        RECT 1558.140 502.300 1559.740 507.500 ;
        RECT 1580.220 505.700 1581.820 507.500 ;
        RECT 1628.060 507.500 1677.500 509.100 ;
        RECT 1628.060 505.700 1629.660 507.500 ;
        RECT 1580.220 504.100 1629.660 505.700 ;
        RECT 1316.180 500.700 1353.660 502.300 ;
        RECT 1482.700 500.700 1559.740 502.300 ;
        RECT 1675.900 502.300 1677.500 507.500 ;
        RECT 1821.260 507.500 1871.620 509.100 ;
        RECT 2061.380 507.500 2078.620 509.100 ;
        RECT 1821.260 505.700 1822.860 507.500 ;
        RECT 1755.020 504.100 1822.860 505.700 ;
        RECT 1870.020 505.700 1871.620 507.500 ;
        RECT 1870.020 504.100 1980.180 505.700 ;
        RECT 2013.540 504.100 2019.740 505.700 ;
        RECT 2077.020 502.300 2078.620 507.500 ;
        RECT 2138.660 507.500 2188.100 509.100 ;
        RECT 2138.660 505.700 2140.260 507.500 ;
        RECT 2123.940 504.100 2140.260 505.700 ;
        RECT 2186.500 505.700 2188.100 507.500 ;
        RECT 2235.260 507.500 2285.620 509.100 ;
        RECT 2235.260 505.700 2236.860 507.500 ;
        RECT 2186.500 504.100 2236.860 505.700 ;
        RECT 2284.020 505.700 2285.620 507.500 ;
        RECT 2331.860 507.500 2367.500 509.100 ;
        RECT 2475.380 508.180 2523.900 509.100 ;
        RECT 2475.380 507.500 2476.980 508.180 ;
        RECT 2479.060 507.500 2523.900 508.180 ;
        RECT 2331.860 505.700 2333.460 507.500 ;
        RECT 2284.020 504.100 2333.460 505.700 ;
        RECT 2365.900 505.700 2367.500 507.500 ;
        RECT 2365.900 504.100 2408.900 505.700 ;
        RECT 2535.180 504.100 2568.060 505.700 ;
        RECT 2123.940 502.300 2125.540 504.100 ;
        RECT 1675.900 500.700 1740.060 502.300 ;
        RECT 2077.020 500.700 2125.540 502.300 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 466.720 869.330 466.780 ;
        RECT 980.330 466.720 980.650 466.780 ;
        RECT 869.010 466.580 980.650 466.720 ;
        RECT 869.010 466.520 869.330 466.580 ;
        RECT 980.330 466.520 980.650 466.580 ;
        RECT 864.870 15.540 865.190 15.600 ;
        RECT 869.010 15.540 869.330 15.600 ;
        RECT 864.870 15.400 869.330 15.540 ;
        RECT 864.870 15.340 865.190 15.400 ;
        RECT 869.010 15.340 869.330 15.400 ;
      LAYER via ;
        RECT 869.040 466.520 869.300 466.780 ;
        RECT 980.360 466.520 980.620 466.780 ;
        RECT 864.900 15.340 865.160 15.600 ;
        RECT 869.040 15.340 869.300 15.600 ;
      LAYER met2 ;
        RECT 980.490 510.340 980.770 514.000 ;
        RECT 980.420 510.000 980.770 510.340 ;
        RECT 980.420 466.810 980.560 510.000 ;
        RECT 869.040 466.490 869.300 466.810 ;
        RECT 980.360 466.490 980.620 466.810 ;
        RECT 869.100 15.630 869.240 466.490 ;
        RECT 864.900 15.310 865.160 15.630 ;
        RECT 869.040 15.310 869.300 15.630 ;
        RECT 864.960 2.400 865.100 15.310 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.470 490.180 938.790 490.240 ;
        RECT 942.150 490.180 942.470 490.240 ;
        RECT 938.470 490.040 942.470 490.180 ;
        RECT 938.470 489.980 938.790 490.040 ;
        RECT 942.150 489.980 942.470 490.040 ;
        RECT 882.350 438.160 882.670 438.220 ;
        RECT 938.470 438.160 938.790 438.220 ;
        RECT 882.350 438.020 938.790 438.160 ;
        RECT 882.350 437.960 882.670 438.020 ;
        RECT 938.470 437.960 938.790 438.020 ;
      LAYER via ;
        RECT 938.500 489.980 938.760 490.240 ;
        RECT 942.180 489.980 942.440 490.240 ;
        RECT 882.380 437.960 882.640 438.220 ;
        RECT 938.500 437.960 938.760 438.220 ;
      LAYER met2 ;
        RECT 943.690 510.410 943.970 514.000 ;
        RECT 942.240 510.270 943.970 510.410 ;
        RECT 942.240 490.270 942.380 510.270 ;
        RECT 943.690 510.000 943.970 510.270 ;
        RECT 938.500 489.950 938.760 490.270 ;
        RECT 942.180 489.950 942.440 490.270 ;
        RECT 938.560 438.250 938.700 489.950 ;
        RECT 882.380 437.930 882.640 438.250 ;
        RECT 938.500 437.930 938.760 438.250 ;
        RECT 882.440 15.370 882.580 437.930 ;
        RECT 882.440 15.230 883.040 15.370 ;
        RECT 882.900 2.400 883.040 15.230 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 308.730 3032.020 309.050 3032.080 ;
        RECT 1222.290 3032.020 1222.610 3032.080 ;
        RECT 308.730 3031.880 1222.610 3032.020 ;
        RECT 308.730 3031.820 309.050 3031.880 ;
        RECT 1222.290 3031.820 1222.610 3031.880 ;
        RECT 308.730 494.260 309.050 494.320 ;
        RECT 897.070 494.260 897.390 494.320 ;
        RECT 308.730 494.120 897.390 494.260 ;
        RECT 308.730 494.060 309.050 494.120 ;
        RECT 897.070 494.060 897.390 494.120 ;
        RECT 897.070 20.300 897.390 20.360 ;
        RECT 900.750 20.300 901.070 20.360 ;
        RECT 897.070 20.160 901.070 20.300 ;
        RECT 897.070 20.100 897.390 20.160 ;
        RECT 900.750 20.100 901.070 20.160 ;
      LAYER via ;
        RECT 308.760 3031.820 309.020 3032.080 ;
        RECT 1222.320 3031.820 1222.580 3032.080 ;
        RECT 308.760 494.060 309.020 494.320 ;
        RECT 897.100 494.060 897.360 494.320 ;
        RECT 897.100 20.100 897.360 20.360 ;
        RECT 900.780 20.100 901.040 20.360 ;
      LAYER met2 ;
        RECT 308.760 3031.790 309.020 3032.110 ;
        RECT 1222.320 3031.790 1222.580 3032.110 ;
        RECT 308.820 494.350 308.960 3031.790 ;
        RECT 1222.380 3010.000 1222.520 3031.790 ;
        RECT 1222.380 3009.340 1222.730 3010.000 ;
        RECT 1222.450 3006.000 1222.730 3009.340 ;
        RECT 308.760 494.030 309.020 494.350 ;
        RECT 897.100 494.030 897.360 494.350 ;
        RECT 897.160 20.390 897.300 494.030 ;
        RECT 897.100 20.070 897.360 20.390 ;
        RECT 900.780 20.070 901.040 20.390 ;
        RECT 900.840 2.400 900.980 20.070 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 362.090 635.020 362.410 635.080 ;
        RECT 393.370 635.020 393.690 635.080 ;
        RECT 362.090 634.880 393.690 635.020 ;
        RECT 362.090 634.820 362.410 634.880 ;
        RECT 393.370 634.820 393.690 634.880 ;
        RECT 362.090 33.560 362.410 33.620 ;
        RECT 918.690 33.560 919.010 33.620 ;
        RECT 362.090 33.420 919.010 33.560 ;
        RECT 362.090 33.360 362.410 33.420 ;
        RECT 918.690 33.360 919.010 33.420 ;
      LAYER via ;
        RECT 362.120 634.820 362.380 635.080 ;
        RECT 393.400 634.820 393.660 635.080 ;
        RECT 362.120 33.360 362.380 33.620 ;
        RECT 918.720 33.360 918.980 33.620 ;
      LAYER met2 ;
        RECT 393.390 640.715 393.670 641.085 ;
        RECT 393.460 635.110 393.600 640.715 ;
        RECT 362.120 634.790 362.380 635.110 ;
        RECT 393.400 634.790 393.660 635.110 ;
        RECT 362.180 33.650 362.320 634.790 ;
        RECT 362.120 33.330 362.380 33.650 ;
        RECT 918.720 33.330 918.980 33.650 ;
        RECT 918.780 2.400 918.920 33.330 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 393.390 640.760 393.670 641.040 ;
      LAYER met3 ;
        RECT 393.365 641.050 393.695 641.065 ;
        RECT 410.000 641.050 414.000 641.200 ;
        RECT 393.365 640.750 414.000 641.050 ;
        RECT 393.365 640.735 393.695 640.750 ;
        RECT 410.000 640.600 414.000 640.750 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.770 501.060 573.090 501.120 ;
        RECT 579.210 501.060 579.530 501.120 ;
        RECT 572.770 500.920 579.530 501.060 ;
        RECT 572.770 500.860 573.090 500.920 ;
        RECT 579.210 500.860 579.530 500.920 ;
        RECT 579.210 80.140 579.530 80.200 ;
        RECT 931.570 80.140 931.890 80.200 ;
        RECT 579.210 80.000 931.890 80.140 ;
        RECT 579.210 79.940 579.530 80.000 ;
        RECT 931.570 79.940 931.890 80.000 ;
        RECT 931.570 2.960 931.890 3.020 ;
        RECT 936.170 2.960 936.490 3.020 ;
        RECT 931.570 2.820 936.490 2.960 ;
        RECT 931.570 2.760 931.890 2.820 ;
        RECT 936.170 2.760 936.490 2.820 ;
      LAYER via ;
        RECT 572.800 500.860 573.060 501.120 ;
        RECT 579.240 500.860 579.500 501.120 ;
        RECT 579.240 79.940 579.500 80.200 ;
        RECT 931.600 79.940 931.860 80.200 ;
        RECT 931.600 2.760 931.860 3.020 ;
        RECT 936.200 2.760 936.460 3.020 ;
      LAYER met2 ;
        RECT 572.930 510.340 573.210 514.000 ;
        RECT 572.860 510.000 573.210 510.340 ;
        RECT 572.860 501.150 573.000 510.000 ;
        RECT 572.800 500.830 573.060 501.150 ;
        RECT 579.240 500.830 579.500 501.150 ;
        RECT 579.300 80.230 579.440 500.830 ;
        RECT 579.240 79.910 579.500 80.230 ;
        RECT 931.600 79.910 931.860 80.230 ;
        RECT 931.660 3.050 931.800 79.910 ;
        RECT 931.600 2.730 931.860 3.050 ;
        RECT 936.200 2.730 936.460 3.050 ;
        RECT 936.260 2.400 936.400 2.730 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 3036.440 324.230 3036.500 ;
        RECT 901.210 3036.440 901.530 3036.500 ;
        RECT 323.910 3036.300 901.530 3036.440 ;
        RECT 323.910 3036.240 324.230 3036.300 ;
        RECT 901.210 3036.240 901.530 3036.300 ;
        RECT 323.910 47.840 324.230 47.900 ;
        RECT 954.110 47.840 954.430 47.900 ;
        RECT 323.910 47.700 954.430 47.840 ;
        RECT 323.910 47.640 324.230 47.700 ;
        RECT 954.110 47.640 954.430 47.700 ;
      LAYER via ;
        RECT 323.940 3036.240 324.200 3036.500 ;
        RECT 901.240 3036.240 901.500 3036.500 ;
        RECT 323.940 47.640 324.200 47.900 ;
        RECT 954.140 47.640 954.400 47.900 ;
      LAYER met2 ;
        RECT 323.940 3036.210 324.200 3036.530 ;
        RECT 901.240 3036.210 901.500 3036.530 ;
        RECT 324.000 47.930 324.140 3036.210 ;
        RECT 901.300 3010.000 901.440 3036.210 ;
        RECT 901.300 3009.340 901.650 3010.000 ;
        RECT 901.370 3006.000 901.650 3009.340 ;
        RECT 323.940 47.610 324.200 47.930 ;
        RECT 954.140 47.610 954.400 47.930 ;
        RECT 954.200 2.400 954.340 47.610 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 389.880 972.830 389.940 ;
        RECT 2408.170 389.880 2408.490 389.940 ;
        RECT 972.510 389.740 2408.490 389.880 ;
        RECT 972.510 389.680 972.830 389.740 ;
        RECT 2408.170 389.680 2408.490 389.740 ;
      LAYER via ;
        RECT 972.540 389.680 972.800 389.940 ;
        RECT 2408.200 389.680 2408.460 389.940 ;
      LAYER met2 ;
        RECT 2413.850 510.410 2414.130 514.000 ;
        RECT 2408.260 510.270 2414.130 510.410 ;
        RECT 2408.260 389.970 2408.400 510.270 ;
        RECT 2413.850 510.000 2414.130 510.270 ;
        RECT 972.540 389.650 972.800 389.970 ;
        RECT 2408.200 389.650 2408.460 389.970 ;
        RECT 972.600 17.410 972.740 389.650 ;
        RECT 972.140 17.270 972.740 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.670 16.900 648.990 16.960 ;
        RECT 650.970 16.900 651.290 16.960 ;
        RECT 648.670 16.760 651.290 16.900 ;
        RECT 648.670 16.700 648.990 16.760 ;
        RECT 650.970 16.700 651.290 16.760 ;
      LAYER via ;
        RECT 648.700 16.700 648.960 16.960 ;
        RECT 651.000 16.700 651.260 16.960 ;
      LAYER met2 ;
        RECT 2148.750 3016.635 2149.030 3017.005 ;
        RECT 2148.820 3010.000 2148.960 3016.635 ;
        RECT 2148.820 3009.340 2149.170 3010.000 ;
        RECT 2148.890 3006.000 2149.170 3009.340 ;
        RECT 648.690 493.155 648.970 493.525 ;
        RECT 648.760 16.990 648.900 493.155 ;
        RECT 648.700 16.670 648.960 16.990 ;
        RECT 651.000 16.670 651.260 16.990 ;
        RECT 651.060 2.400 651.200 16.670 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 2148.750 3016.680 2149.030 3016.960 ;
        RECT 648.690 493.200 648.970 493.480 ;
      LAYER met3 ;
        RECT 361.830 3016.970 362.210 3016.980 ;
        RECT 2148.725 3016.970 2149.055 3016.985 ;
        RECT 361.830 3016.670 2149.055 3016.970 ;
        RECT 361.830 3016.660 362.210 3016.670 ;
        RECT 2148.725 3016.655 2149.055 3016.670 ;
        RECT 361.830 493.490 362.210 493.500 ;
        RECT 648.665 493.490 648.995 493.505 ;
        RECT 361.830 493.190 648.995 493.490 ;
        RECT 361.830 493.180 362.210 493.190 ;
        RECT 648.665 493.175 648.995 493.190 ;
      LAYER via3 ;
        RECT 361.860 3016.660 362.180 3016.980 ;
        RECT 361.860 493.180 362.180 493.500 ;
      LAYER met4 ;
        RECT 361.855 3016.655 362.185 3016.985 ;
        RECT 361.870 493.505 362.170 3016.655 ;
        RECT 361.855 493.175 362.185 493.505 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 992.365 386.325 992.535 434.775 ;
        RECT 992.365 338.045 992.535 385.815 ;
        RECT 992.365 241.485 992.535 289.595 ;
        RECT 992.365 158.185 992.535 193.035 ;
      LAYER mcon ;
        RECT 992.365 434.605 992.535 434.775 ;
        RECT 992.365 385.645 992.535 385.815 ;
        RECT 992.365 289.425 992.535 289.595 ;
        RECT 992.365 192.865 992.535 193.035 ;
      LAYER met1 ;
        RECT 2520.410 1118.160 2520.730 1118.220 ;
        RECT 2562.270 1118.160 2562.590 1118.220 ;
        RECT 2520.410 1118.020 2562.590 1118.160 ;
        RECT 2520.410 1117.960 2520.730 1118.020 ;
        RECT 2562.270 1117.960 2562.590 1118.020 ;
        RECT 993.670 507.520 993.990 507.580 ;
        RECT 2562.270 507.520 2562.590 507.580 ;
        RECT 993.670 507.380 2562.590 507.520 ;
        RECT 993.670 507.320 993.990 507.380 ;
        RECT 2562.270 507.320 2562.590 507.380 ;
        RECT 992.305 434.760 992.595 434.805 ;
        RECT 992.750 434.760 993.070 434.820 ;
        RECT 992.305 434.620 993.070 434.760 ;
        RECT 992.305 434.575 992.595 434.620 ;
        RECT 992.750 434.560 993.070 434.620 ;
        RECT 992.290 386.480 992.610 386.540 ;
        RECT 992.095 386.340 992.610 386.480 ;
        RECT 992.290 386.280 992.610 386.340 ;
        RECT 992.290 385.800 992.610 385.860 ;
        RECT 992.095 385.660 992.610 385.800 ;
        RECT 992.290 385.600 992.610 385.660 ;
        RECT 992.305 338.200 992.595 338.245 ;
        RECT 992.750 338.200 993.070 338.260 ;
        RECT 992.305 338.060 993.070 338.200 ;
        RECT 992.305 338.015 992.595 338.060 ;
        RECT 992.750 338.000 993.070 338.060 ;
        RECT 992.750 304.200 993.070 304.260 ;
        RECT 992.380 304.060 993.070 304.200 ;
        RECT 992.380 303.580 992.520 304.060 ;
        RECT 992.750 304.000 993.070 304.060 ;
        RECT 992.290 303.320 992.610 303.580 ;
        RECT 992.290 289.580 992.610 289.640 ;
        RECT 992.095 289.440 992.610 289.580 ;
        RECT 992.290 289.380 992.610 289.440 ;
        RECT 992.305 241.640 992.595 241.685 ;
        RECT 992.750 241.640 993.070 241.700 ;
        RECT 992.305 241.500 993.070 241.640 ;
        RECT 992.305 241.455 992.595 241.500 ;
        RECT 992.750 241.440 993.070 241.500 ;
        RECT 992.750 207.300 993.070 207.360 ;
        RECT 992.380 207.160 993.070 207.300 ;
        RECT 992.380 207.020 992.520 207.160 ;
        RECT 992.750 207.100 993.070 207.160 ;
        RECT 992.290 206.760 992.610 207.020 ;
        RECT 992.290 193.020 992.610 193.080 ;
        RECT 992.095 192.880 992.610 193.020 ;
        RECT 992.290 192.820 992.610 192.880 ;
        RECT 992.305 158.340 992.595 158.385 ;
        RECT 992.750 158.340 993.070 158.400 ;
        RECT 992.305 158.200 993.070 158.340 ;
        RECT 992.305 158.155 992.595 158.200 ;
        RECT 992.750 158.140 993.070 158.200 ;
        RECT 989.990 20.300 990.310 20.360 ;
        RECT 993.210 20.300 993.530 20.360 ;
        RECT 989.990 20.160 993.530 20.300 ;
        RECT 989.990 20.100 990.310 20.160 ;
        RECT 993.210 20.100 993.530 20.160 ;
      LAYER via ;
        RECT 2520.440 1117.960 2520.700 1118.220 ;
        RECT 2562.300 1117.960 2562.560 1118.220 ;
        RECT 993.700 507.320 993.960 507.580 ;
        RECT 2562.300 507.320 2562.560 507.580 ;
        RECT 992.780 434.560 993.040 434.820 ;
        RECT 992.320 386.280 992.580 386.540 ;
        RECT 992.320 385.600 992.580 385.860 ;
        RECT 992.780 338.000 993.040 338.260 ;
        RECT 992.780 304.000 993.040 304.260 ;
        RECT 992.320 303.320 992.580 303.580 ;
        RECT 992.320 289.380 992.580 289.640 ;
        RECT 992.780 241.440 993.040 241.700 ;
        RECT 992.780 207.100 993.040 207.360 ;
        RECT 992.320 206.760 992.580 207.020 ;
        RECT 992.320 192.820 992.580 193.080 ;
        RECT 992.780 158.140 993.040 158.400 ;
        RECT 990.020 20.100 990.280 20.360 ;
        RECT 993.240 20.100 993.500 20.360 ;
      LAYER met2 ;
        RECT 2520.430 1123.515 2520.710 1123.885 ;
        RECT 2520.500 1118.250 2520.640 1123.515 ;
        RECT 2520.440 1117.930 2520.700 1118.250 ;
        RECT 2562.300 1117.930 2562.560 1118.250 ;
        RECT 2562.360 507.610 2562.500 1117.930 ;
        RECT 993.700 507.290 993.960 507.610 ;
        RECT 2562.300 507.290 2562.560 507.610 ;
        RECT 993.760 483.325 993.900 507.290 ;
        RECT 991.850 482.955 992.130 483.325 ;
        RECT 993.690 482.955 993.970 483.325 ;
        RECT 991.920 448.530 992.060 482.955 ;
        RECT 991.920 448.390 992.980 448.530 ;
        RECT 992.840 434.850 992.980 448.390 ;
        RECT 992.780 434.530 993.040 434.850 ;
        RECT 992.320 386.250 992.580 386.570 ;
        RECT 992.380 385.890 992.520 386.250 ;
        RECT 992.320 385.570 992.580 385.890 ;
        RECT 992.780 337.970 993.040 338.290 ;
        RECT 992.840 304.290 992.980 337.970 ;
        RECT 992.780 303.970 993.040 304.290 ;
        RECT 992.320 303.290 992.580 303.610 ;
        RECT 992.380 289.670 992.520 303.290 ;
        RECT 992.320 289.350 992.580 289.670 ;
        RECT 992.780 241.410 993.040 241.730 ;
        RECT 992.840 207.390 992.980 241.410 ;
        RECT 992.780 207.070 993.040 207.390 ;
        RECT 992.320 206.730 992.580 207.050 ;
        RECT 992.380 193.110 992.520 206.730 ;
        RECT 992.320 192.790 992.580 193.110 ;
        RECT 992.780 158.110 993.040 158.430 ;
        RECT 992.840 109.890 992.980 158.110 ;
        RECT 992.840 109.750 993.440 109.890 ;
        RECT 993.300 20.390 993.440 109.750 ;
        RECT 990.020 20.070 990.280 20.390 ;
        RECT 993.240 20.070 993.500 20.390 ;
        RECT 990.080 2.400 990.220 20.070 ;
        RECT 989.870 -4.800 990.430 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1123.560 2520.710 1123.840 ;
        RECT 991.850 483.000 992.130 483.280 ;
        RECT 993.690 483.000 993.970 483.280 ;
      LAYER met3 ;
        RECT 2506.000 1123.850 2510.000 1124.000 ;
        RECT 2520.405 1123.850 2520.735 1123.865 ;
        RECT 2506.000 1123.550 2520.735 1123.850 ;
        RECT 2506.000 1123.400 2510.000 1123.550 ;
        RECT 2520.405 1123.535 2520.735 1123.550 ;
        RECT 991.825 483.290 992.155 483.305 ;
        RECT 993.665 483.290 993.995 483.305 ;
        RECT 991.825 482.990 993.995 483.290 ;
        RECT 991.825 482.975 992.155 482.990 ;
        RECT 993.665 482.975 993.995 482.990 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1013.910 80.480 1014.230 80.540 ;
        RECT 1842.370 80.480 1842.690 80.540 ;
        RECT 1013.910 80.340 1842.690 80.480 ;
        RECT 1013.910 80.280 1014.230 80.340 ;
        RECT 1842.370 80.280 1842.690 80.340 ;
        RECT 1007.470 20.300 1007.790 20.360 ;
        RECT 1013.910 20.300 1014.230 20.360 ;
        RECT 1007.470 20.160 1014.230 20.300 ;
        RECT 1007.470 20.100 1007.790 20.160 ;
        RECT 1013.910 20.100 1014.230 20.160 ;
      LAYER via ;
        RECT 1013.940 80.280 1014.200 80.540 ;
        RECT 1842.400 80.280 1842.660 80.540 ;
        RECT 1007.500 20.100 1007.760 20.360 ;
        RECT 1013.940 20.100 1014.200 20.360 ;
      LAYER met2 ;
        RECT 1845.290 510.410 1845.570 514.000 ;
        RECT 1842.460 510.270 1845.570 510.410 ;
        RECT 1842.460 80.570 1842.600 510.270 ;
        RECT 1845.290 510.000 1845.570 510.270 ;
        RECT 1013.940 80.250 1014.200 80.570 ;
        RECT 1842.400 80.250 1842.660 80.570 ;
        RECT 1014.000 20.390 1014.140 80.250 ;
        RECT 1007.500 20.070 1007.760 20.390 ;
        RECT 1013.940 20.070 1014.200 20.390 ;
        RECT 1007.560 2.400 1007.700 20.070 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 375.940 600.230 376.000 ;
        RECT 1021.270 375.940 1021.590 376.000 ;
        RECT 599.910 375.800 1021.590 375.940 ;
        RECT 599.910 375.740 600.230 375.800 ;
        RECT 1021.270 375.740 1021.590 375.800 ;
        RECT 1021.270 62.120 1021.590 62.180 ;
        RECT 1025.410 62.120 1025.730 62.180 ;
        RECT 1021.270 61.980 1025.730 62.120 ;
        RECT 1021.270 61.920 1021.590 61.980 ;
        RECT 1025.410 61.920 1025.730 61.980 ;
      LAYER via ;
        RECT 599.940 375.740 600.200 376.000 ;
        RECT 1021.300 375.740 1021.560 376.000 ;
        RECT 1021.300 61.920 1021.560 62.180 ;
        RECT 1025.440 61.920 1025.700 62.180 ;
      LAYER met2 ;
        RECT 597.770 510.410 598.050 514.000 ;
        RECT 597.770 510.270 600.140 510.410 ;
        RECT 597.770 510.000 598.050 510.270 ;
        RECT 600.000 376.030 600.140 510.270 ;
        RECT 599.940 375.710 600.200 376.030 ;
        RECT 1021.300 375.710 1021.560 376.030 ;
        RECT 1021.360 62.210 1021.500 375.710 ;
        RECT 1021.300 61.890 1021.560 62.210 ;
        RECT 1025.440 61.890 1025.700 62.210 ;
        RECT 1025.500 2.400 1025.640 61.890 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 20.300 1043.670 20.360 ;
        RECT 1048.410 20.300 1048.730 20.360 ;
        RECT 1043.350 20.160 1048.730 20.300 ;
        RECT 1043.350 20.100 1043.670 20.160 ;
        RECT 1048.410 20.100 1048.730 20.160 ;
      LAYER via ;
        RECT 1043.380 20.100 1043.640 20.360 ;
        RECT 1048.440 20.100 1048.700 20.360 ;
      LAYER met2 ;
        RECT 1048.430 438.075 1048.710 438.445 ;
        RECT 1048.500 20.390 1048.640 438.075 ;
        RECT 1043.380 20.070 1043.640 20.390 ;
        RECT 1048.440 20.070 1048.700 20.390 ;
        RECT 1043.440 2.400 1043.580 20.070 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1048.430 438.120 1048.710 438.400 ;
      LAYER met3 ;
        RECT 2506.000 2785.770 2510.000 2785.920 ;
        RECT 2532.110 2785.770 2532.490 2785.780 ;
        RECT 2506.000 2785.470 2532.490 2785.770 ;
        RECT 2506.000 2785.320 2510.000 2785.470 ;
        RECT 2532.110 2785.460 2532.490 2785.470 ;
        RECT 2532.110 439.090 2532.490 439.100 ;
        RECT 2500.870 438.790 2532.490 439.090 ;
        RECT 1048.405 438.410 1048.735 438.425 ;
        RECT 2500.870 438.410 2501.170 438.790 ;
        RECT 2532.110 438.780 2532.490 438.790 ;
        RECT 1048.405 438.110 2501.170 438.410 ;
        RECT 1048.405 438.095 1048.735 438.110 ;
      LAYER via3 ;
        RECT 2532.140 2785.460 2532.460 2785.780 ;
        RECT 2532.140 438.780 2532.460 439.100 ;
      LAYER met4 ;
        RECT 2532.135 2785.455 2532.465 2785.785 ;
        RECT 2532.150 439.105 2532.450 2785.455 ;
        RECT 2532.135 438.775 2532.465 439.105 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1062.285 241.485 1062.455 289.595 ;
        RECT 1062.285 48.365 1062.455 96.475 ;
      LAYER mcon ;
        RECT 1062.285 289.425 1062.455 289.595 ;
        RECT 1062.285 96.305 1062.455 96.475 ;
      LAYER met1 ;
        RECT 2519.950 1814.820 2520.270 1814.880 ;
        RECT 2582.970 1814.820 2583.290 1814.880 ;
        RECT 2519.950 1814.680 2583.290 1814.820 ;
        RECT 2519.950 1814.620 2520.270 1814.680 ;
        RECT 2582.970 1814.620 2583.290 1814.680 ;
        RECT 1061.290 483.380 1061.610 483.440 ;
        RECT 1061.750 483.380 1062.070 483.440 ;
        RECT 1061.290 483.240 1062.070 483.380 ;
        RECT 1061.290 483.180 1061.610 483.240 ;
        RECT 1061.750 483.180 1062.070 483.240 ;
        RECT 1062.210 289.580 1062.530 289.640 ;
        RECT 1062.015 289.440 1062.530 289.580 ;
        RECT 1062.210 289.380 1062.530 289.440 ;
        RECT 1062.210 241.640 1062.530 241.700 ;
        RECT 1062.015 241.500 1062.530 241.640 ;
        RECT 1062.210 241.440 1062.530 241.500 ;
        RECT 1062.210 96.460 1062.530 96.520 ;
        RECT 1062.015 96.320 1062.530 96.460 ;
        RECT 1062.210 96.260 1062.530 96.320 ;
        RECT 1062.210 48.520 1062.530 48.580 ;
        RECT 1062.015 48.380 1062.530 48.520 ;
        RECT 1062.210 48.320 1062.530 48.380 ;
        RECT 1062.210 14.180 1062.530 14.240 ;
        RECT 1061.380 14.040 1062.530 14.180 ;
        RECT 1061.380 13.900 1061.520 14.040 ;
        RECT 1062.210 13.980 1062.530 14.040 ;
        RECT 1061.290 13.640 1061.610 13.900 ;
      LAYER via ;
        RECT 2519.980 1814.620 2520.240 1814.880 ;
        RECT 2583.000 1814.620 2583.260 1814.880 ;
        RECT 1061.320 483.180 1061.580 483.440 ;
        RECT 1061.780 483.180 1062.040 483.440 ;
        RECT 1062.240 289.380 1062.500 289.640 ;
        RECT 1062.240 241.440 1062.500 241.700 ;
        RECT 1062.240 96.260 1062.500 96.520 ;
        RECT 1062.240 48.320 1062.500 48.580 ;
        RECT 1062.240 13.980 1062.500 14.240 ;
        RECT 1061.320 13.640 1061.580 13.900 ;
      LAYER met2 ;
        RECT 2519.970 1818.475 2520.250 1818.845 ;
        RECT 2520.040 1814.910 2520.180 1818.475 ;
        RECT 2519.980 1814.590 2520.240 1814.910 ;
        RECT 2583.000 1814.590 2583.260 1814.910 ;
        RECT 2583.060 507.805 2583.200 1814.590 ;
        RECT 1061.310 507.435 1061.590 507.805 ;
        RECT 2582.990 507.435 2583.270 507.805 ;
        RECT 1061.380 483.470 1061.520 507.435 ;
        RECT 1061.320 483.150 1061.580 483.470 ;
        RECT 1061.780 483.210 1062.040 483.470 ;
        RECT 1061.780 483.150 1062.440 483.210 ;
        RECT 1061.840 483.070 1062.440 483.150 ;
        RECT 1062.300 482.530 1062.440 483.070 ;
        RECT 1061.840 482.390 1062.440 482.530 ;
        RECT 1061.840 458.730 1061.980 482.390 ;
        RECT 1061.840 458.590 1062.440 458.730 ;
        RECT 1062.300 289.670 1062.440 458.590 ;
        RECT 1062.240 289.350 1062.500 289.670 ;
        RECT 1062.240 241.410 1062.500 241.730 ;
        RECT 1062.300 96.550 1062.440 241.410 ;
        RECT 1062.240 96.230 1062.500 96.550 ;
        RECT 1062.240 48.290 1062.500 48.610 ;
        RECT 1062.300 14.270 1062.440 48.290 ;
        RECT 1062.240 13.950 1062.500 14.270 ;
        RECT 1061.320 13.610 1061.580 13.930 ;
        RECT 1061.380 2.400 1061.520 13.610 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
      LAYER via2 ;
        RECT 2519.970 1818.520 2520.250 1818.800 ;
        RECT 1061.310 507.480 1061.590 507.760 ;
        RECT 2582.990 507.480 2583.270 507.760 ;
      LAYER met3 ;
        RECT 2506.000 1818.810 2510.000 1818.960 ;
        RECT 2519.945 1818.810 2520.275 1818.825 ;
        RECT 2506.000 1818.510 2520.275 1818.810 ;
        RECT 2506.000 1818.360 2510.000 1818.510 ;
        RECT 2519.945 1818.495 2520.275 1818.510 ;
        RECT 1061.285 507.770 1061.615 507.785 ;
        RECT 2582.965 507.770 2583.295 507.785 ;
        RECT 1061.285 507.470 2583.295 507.770 ;
        RECT 1061.285 507.455 1061.615 507.470 ;
        RECT 2582.965 507.455 2583.295 507.470 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2180.660 2519.810 2180.720 ;
        RECT 2595.390 2180.660 2595.710 2180.720 ;
        RECT 2519.490 2180.520 2595.710 2180.660 ;
        RECT 2519.490 2180.460 2519.810 2180.520 ;
        RECT 2595.390 2180.460 2595.710 2180.520 ;
        RECT 1082.910 493.240 1083.230 493.300 ;
        RECT 2595.390 493.240 2595.710 493.300 ;
        RECT 1082.910 493.100 2595.710 493.240 ;
        RECT 1082.910 493.040 1083.230 493.100 ;
        RECT 2595.390 493.040 2595.710 493.100 ;
        RECT 1079.230 15.880 1079.550 15.940 ;
        RECT 1082.910 15.880 1083.230 15.940 ;
        RECT 1079.230 15.740 1083.230 15.880 ;
        RECT 1079.230 15.680 1079.550 15.740 ;
        RECT 1082.910 15.680 1083.230 15.740 ;
      LAYER via ;
        RECT 2519.520 2180.460 2519.780 2180.720 ;
        RECT 2595.420 2180.460 2595.680 2180.720 ;
        RECT 1082.940 493.040 1083.200 493.300 ;
        RECT 2595.420 493.040 2595.680 493.300 ;
        RECT 1079.260 15.680 1079.520 15.940 ;
        RECT 1082.940 15.680 1083.200 15.940 ;
      LAYER met2 ;
        RECT 2519.510 2182.955 2519.790 2183.325 ;
        RECT 2519.580 2180.750 2519.720 2182.955 ;
        RECT 2519.520 2180.430 2519.780 2180.750 ;
        RECT 2595.420 2180.430 2595.680 2180.750 ;
        RECT 2595.480 493.330 2595.620 2180.430 ;
        RECT 1082.940 493.010 1083.200 493.330 ;
        RECT 2595.420 493.010 2595.680 493.330 ;
        RECT 1083.000 15.970 1083.140 493.010 ;
        RECT 1079.260 15.650 1079.520 15.970 ;
        RECT 1082.940 15.650 1083.200 15.970 ;
        RECT 1079.320 2.400 1079.460 15.650 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2183.000 2519.790 2183.280 ;
      LAYER met3 ;
        RECT 2506.000 2183.290 2510.000 2183.440 ;
        RECT 2519.485 2183.290 2519.815 2183.305 ;
        RECT 2506.000 2182.990 2519.815 2183.290 ;
        RECT 2506.000 2182.840 2510.000 2182.990 ;
        RECT 2519.485 2182.975 2519.815 2182.990 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 336.330 3024.880 336.650 3024.940 ;
        RECT 1110.970 3024.880 1111.290 3024.940 ;
        RECT 336.330 3024.740 1111.290 3024.880 ;
        RECT 336.330 3024.680 336.650 3024.740 ;
        RECT 1110.970 3024.680 1111.290 3024.740 ;
        RECT 336.330 493.580 336.650 493.640 ;
        RECT 1090.270 493.580 1090.590 493.640 ;
        RECT 336.330 493.440 1090.590 493.580 ;
        RECT 336.330 493.380 336.650 493.440 ;
        RECT 1090.270 493.380 1090.590 493.440 ;
        RECT 1090.270 20.300 1090.590 20.360 ;
        RECT 1096.710 20.300 1097.030 20.360 ;
        RECT 1090.270 20.160 1097.030 20.300 ;
        RECT 1090.270 20.100 1090.590 20.160 ;
        RECT 1096.710 20.100 1097.030 20.160 ;
      LAYER via ;
        RECT 336.360 3024.680 336.620 3024.940 ;
        RECT 1111.000 3024.680 1111.260 3024.940 ;
        RECT 336.360 493.380 336.620 493.640 ;
        RECT 1090.300 493.380 1090.560 493.640 ;
        RECT 1090.300 20.100 1090.560 20.360 ;
        RECT 1096.740 20.100 1097.000 20.360 ;
      LAYER met2 ;
        RECT 336.360 3024.650 336.620 3024.970 ;
        RECT 1111.000 3024.650 1111.260 3024.970 ;
        RECT 336.420 493.670 336.560 3024.650 ;
        RECT 1111.060 3010.000 1111.200 3024.650 ;
        RECT 1111.060 3009.340 1111.410 3010.000 ;
        RECT 1111.130 3006.000 1111.410 3009.340 ;
        RECT 336.360 493.350 336.620 493.670 ;
        RECT 1090.300 493.350 1090.560 493.670 ;
        RECT 1090.360 20.390 1090.500 493.350 ;
        RECT 1090.300 20.070 1090.560 20.390 ;
        RECT 1096.740 20.070 1097.000 20.390 ;
        RECT 1096.800 2.400 1096.940 20.070 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 316.090 2028.680 316.410 2028.740 ;
        RECT 393.370 2028.680 393.690 2028.740 ;
        RECT 316.090 2028.540 393.690 2028.680 ;
        RECT 316.090 2028.480 316.410 2028.540 ;
        RECT 393.370 2028.480 393.690 2028.540 ;
        RECT 316.090 18.260 316.410 18.320 ;
        RECT 1114.650 18.260 1114.970 18.320 ;
        RECT 316.090 18.120 1114.970 18.260 ;
        RECT 316.090 18.060 316.410 18.120 ;
        RECT 1114.650 18.060 1114.970 18.120 ;
      LAYER via ;
        RECT 316.120 2028.480 316.380 2028.740 ;
        RECT 393.400 2028.480 393.660 2028.740 ;
        RECT 316.120 18.060 316.380 18.320 ;
        RECT 1114.680 18.060 1114.940 18.320 ;
      LAYER met2 ;
        RECT 393.390 2029.275 393.670 2029.645 ;
        RECT 393.460 2028.770 393.600 2029.275 ;
        RECT 316.120 2028.450 316.380 2028.770 ;
        RECT 393.400 2028.450 393.660 2028.770 ;
        RECT 316.180 18.350 316.320 2028.450 ;
        RECT 316.120 18.030 316.380 18.350 ;
        RECT 1114.680 18.030 1114.940 18.350 ;
        RECT 1114.740 2.400 1114.880 18.030 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 393.390 2029.320 393.670 2029.600 ;
      LAYER met3 ;
        RECT 393.365 2029.610 393.695 2029.625 ;
        RECT 410.000 2029.610 414.000 2029.760 ;
        RECT 393.365 2029.310 414.000 2029.610 ;
        RECT 393.365 2029.295 393.695 2029.310 ;
        RECT 410.000 2029.160 414.000 2029.310 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1104.560 2520.730 1104.620 ;
        RECT 2548.470 1104.560 2548.790 1104.620 ;
        RECT 2520.410 1104.420 2548.790 1104.560 ;
        RECT 2520.410 1104.360 2520.730 1104.420 ;
        RECT 2548.470 1104.360 2548.790 1104.420 ;
        RECT 1138.110 493.580 1138.430 493.640 ;
        RECT 2548.470 493.580 2548.790 493.640 ;
        RECT 1138.110 493.440 2548.790 493.580 ;
        RECT 1138.110 493.380 1138.430 493.440 ;
        RECT 2548.470 493.380 2548.790 493.440 ;
        RECT 1132.590 16.900 1132.910 16.960 ;
        RECT 1138.110 16.900 1138.430 16.960 ;
        RECT 1132.590 16.760 1138.430 16.900 ;
        RECT 1132.590 16.700 1132.910 16.760 ;
        RECT 1138.110 16.700 1138.430 16.760 ;
      LAYER via ;
        RECT 2520.440 1104.360 2520.700 1104.620 ;
        RECT 2548.500 1104.360 2548.760 1104.620 ;
        RECT 1138.140 493.380 1138.400 493.640 ;
        RECT 2548.500 493.380 2548.760 493.640 ;
        RECT 1132.620 16.700 1132.880 16.960 ;
        RECT 1138.140 16.700 1138.400 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1105.835 2520.710 1106.205 ;
        RECT 2520.500 1104.650 2520.640 1105.835 ;
        RECT 2520.440 1104.330 2520.700 1104.650 ;
        RECT 2548.500 1104.330 2548.760 1104.650 ;
        RECT 2548.560 493.670 2548.700 1104.330 ;
        RECT 1138.140 493.350 1138.400 493.670 ;
        RECT 2548.500 493.350 2548.760 493.670 ;
        RECT 1138.200 16.990 1138.340 493.350 ;
        RECT 1132.620 16.670 1132.880 16.990 ;
        RECT 1138.140 16.670 1138.400 16.990 ;
        RECT 1132.680 2.400 1132.820 16.670 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1105.880 2520.710 1106.160 ;
      LAYER met3 ;
        RECT 2506.000 1106.170 2510.000 1106.320 ;
        RECT 2520.405 1106.170 2520.735 1106.185 ;
        RECT 2506.000 1105.870 2520.735 1106.170 ;
        RECT 2506.000 1105.720 2510.000 1105.870 ;
        RECT 2520.405 1105.855 2520.735 1105.870 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.250 3036.100 406.570 3036.160 ;
        RECT 1024.490 3036.100 1024.810 3036.160 ;
        RECT 406.250 3035.960 1024.810 3036.100 ;
        RECT 406.250 3035.900 406.570 3035.960 ;
        RECT 1024.490 3035.900 1024.810 3035.960 ;
        RECT 406.250 61.780 406.570 61.840 ;
        RECT 1145.470 61.780 1145.790 61.840 ;
        RECT 406.250 61.640 1145.790 61.780 ;
        RECT 406.250 61.580 406.570 61.640 ;
        RECT 1145.470 61.580 1145.790 61.640 ;
      LAYER via ;
        RECT 406.280 3035.900 406.540 3036.160 ;
        RECT 1024.520 3035.900 1024.780 3036.160 ;
        RECT 406.280 61.580 406.540 61.840 ;
        RECT 1145.500 61.580 1145.760 61.840 ;
      LAYER met2 ;
        RECT 406.280 3035.870 406.540 3036.190 ;
        RECT 1024.520 3035.870 1024.780 3036.190 ;
        RECT 406.340 61.870 406.480 3035.870 ;
        RECT 1024.580 3010.000 1024.720 3035.870 ;
        RECT 1024.580 3009.340 1024.930 3010.000 ;
        RECT 1024.650 3006.000 1024.930 3009.340 ;
        RECT 406.280 61.550 406.540 61.870 ;
        RECT 1145.500 61.550 1145.760 61.870 ;
        RECT 1145.560 17.410 1145.700 61.550 ;
        RECT 1145.560 17.270 1150.760 17.410 ;
        RECT 1150.620 2.400 1150.760 17.270 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 322.070 2208.200 322.390 2208.260 ;
        RECT 393.370 2208.200 393.690 2208.260 ;
        RECT 322.070 2208.060 393.690 2208.200 ;
        RECT 322.070 2208.000 322.390 2208.060 ;
        RECT 393.370 2208.000 393.690 2208.060 ;
        RECT 322.070 20.640 322.390 20.700 ;
        RECT 668.910 20.640 669.230 20.700 ;
        RECT 322.070 20.500 669.230 20.640 ;
        RECT 322.070 20.440 322.390 20.500 ;
        RECT 668.910 20.440 669.230 20.500 ;
      LAYER via ;
        RECT 322.100 2208.000 322.360 2208.260 ;
        RECT 393.400 2208.000 393.660 2208.260 ;
        RECT 322.100 20.440 322.360 20.700 ;
        RECT 668.940 20.440 669.200 20.700 ;
      LAYER met2 ;
        RECT 393.390 2211.515 393.670 2211.885 ;
        RECT 393.460 2208.290 393.600 2211.515 ;
        RECT 322.100 2207.970 322.360 2208.290 ;
        RECT 393.400 2207.970 393.660 2208.290 ;
        RECT 322.160 20.730 322.300 2207.970 ;
        RECT 322.100 20.410 322.360 20.730 ;
        RECT 668.940 20.410 669.200 20.730 ;
        RECT 669.000 2.400 669.140 20.410 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 393.390 2211.560 393.670 2211.840 ;
      LAYER met3 ;
        RECT 393.365 2211.850 393.695 2211.865 ;
        RECT 410.000 2211.850 414.000 2212.000 ;
        RECT 393.365 2211.550 414.000 2211.850 ;
        RECT 393.365 2211.535 393.695 2211.550 ;
        RECT 410.000 2211.400 414.000 2211.550 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1082.450 120.940 1082.770 121.000 ;
        RECT 1166.630 120.940 1166.950 121.000 ;
        RECT 1082.450 120.800 1166.950 120.940 ;
        RECT 1082.450 120.740 1082.770 120.800 ;
        RECT 1166.630 120.740 1166.950 120.800 ;
      LAYER via ;
        RECT 1082.480 120.740 1082.740 121.000 ;
        RECT 1166.660 120.740 1166.920 121.000 ;
      LAYER met2 ;
        RECT 1079.850 510.410 1080.130 514.000 ;
        RECT 1079.850 510.270 1082.680 510.410 ;
        RECT 1079.850 510.000 1080.130 510.270 ;
        RECT 1082.540 121.030 1082.680 510.270 ;
        RECT 1082.480 120.710 1082.740 121.030 ;
        RECT 1166.660 120.710 1166.920 121.030 ;
        RECT 1166.720 16.730 1166.860 120.710 ;
        RECT 1166.720 16.590 1168.700 16.730 ;
        RECT 1168.560 2.400 1168.700 16.590 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2836.180 2519.810 2836.240 ;
        RECT 2589.870 2836.180 2590.190 2836.240 ;
        RECT 2519.490 2836.040 2590.190 2836.180 ;
        RECT 2519.490 2835.980 2519.810 2836.040 ;
        RECT 2589.870 2835.980 2590.190 2836.040 ;
      LAYER via ;
        RECT 2519.520 2835.980 2519.780 2836.240 ;
        RECT 2589.900 2835.980 2590.160 2836.240 ;
      LAYER met2 ;
        RECT 2519.510 2841.195 2519.790 2841.565 ;
        RECT 2519.580 2836.270 2519.720 2841.195 ;
        RECT 2519.520 2835.950 2519.780 2836.270 ;
        RECT 2589.900 2835.950 2590.160 2836.270 ;
        RECT 2589.960 493.525 2590.100 2835.950 ;
        RECT 1186.430 493.155 1186.710 493.525 ;
        RECT 2589.890 493.155 2590.170 493.525 ;
        RECT 1186.500 17.410 1186.640 493.155 ;
        RECT 1186.040 17.270 1186.640 17.410 ;
        RECT 1186.040 2.400 1186.180 17.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2841.240 2519.790 2841.520 ;
        RECT 1186.430 493.200 1186.710 493.480 ;
        RECT 2589.890 493.200 2590.170 493.480 ;
      LAYER met3 ;
        RECT 2506.000 2841.530 2510.000 2841.680 ;
        RECT 2519.485 2841.530 2519.815 2841.545 ;
        RECT 2506.000 2841.230 2519.815 2841.530 ;
        RECT 2506.000 2841.080 2510.000 2841.230 ;
        RECT 2519.485 2841.215 2519.815 2841.230 ;
        RECT 1186.405 493.490 1186.735 493.505 ;
        RECT 2589.865 493.490 2590.195 493.505 ;
        RECT 1186.405 493.190 2590.195 493.490 ;
        RECT 1186.405 493.175 1186.735 493.190 ;
        RECT 2589.865 493.175 2590.195 493.190 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1594.160 2520.730 1594.220 ;
        RECT 2575.610 1594.160 2575.930 1594.220 ;
        RECT 2520.410 1594.020 2575.930 1594.160 ;
        RECT 2520.410 1593.960 2520.730 1594.020 ;
        RECT 2575.610 1593.960 2575.930 1594.020 ;
        RECT 1207.110 493.920 1207.430 493.980 ;
        RECT 2575.610 493.920 2575.930 493.980 ;
        RECT 1207.110 493.780 2575.930 493.920 ;
        RECT 1207.110 493.720 1207.430 493.780 ;
        RECT 2575.610 493.720 2575.930 493.780 ;
        RECT 1203.890 16.900 1204.210 16.960 ;
        RECT 1207.110 16.900 1207.430 16.960 ;
        RECT 1203.890 16.760 1207.430 16.900 ;
        RECT 1203.890 16.700 1204.210 16.760 ;
        RECT 1207.110 16.700 1207.430 16.760 ;
      LAYER via ;
        RECT 2520.440 1593.960 2520.700 1594.220 ;
        RECT 2575.640 1593.960 2575.900 1594.220 ;
        RECT 1207.140 493.720 1207.400 493.980 ;
        RECT 2575.640 493.720 2575.900 493.980 ;
        RECT 1203.920 16.700 1204.180 16.960 ;
        RECT 1207.140 16.700 1207.400 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1599.515 2520.710 1599.885 ;
        RECT 2520.500 1594.250 2520.640 1599.515 ;
        RECT 2520.440 1593.930 2520.700 1594.250 ;
        RECT 2575.640 1593.930 2575.900 1594.250 ;
        RECT 2575.700 494.010 2575.840 1593.930 ;
        RECT 1207.140 493.690 1207.400 494.010 ;
        RECT 2575.640 493.690 2575.900 494.010 ;
        RECT 1207.200 16.990 1207.340 493.690 ;
        RECT 1203.920 16.670 1204.180 16.990 ;
        RECT 1207.140 16.670 1207.400 16.990 ;
        RECT 1203.980 2.400 1204.120 16.670 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1599.560 2520.710 1599.840 ;
      LAYER met3 ;
        RECT 2506.000 1599.850 2510.000 1600.000 ;
        RECT 2520.405 1599.850 2520.735 1599.865 ;
        RECT 2506.000 1599.550 2520.735 1599.850 ;
        RECT 2506.000 1599.400 2510.000 1599.550 ;
        RECT 2520.405 1599.535 2520.735 1599.550 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 328.050 855.680 328.370 855.740 ;
        RECT 393.370 855.680 393.690 855.740 ;
        RECT 328.050 855.540 393.690 855.680 ;
        RECT 328.050 855.480 328.370 855.540 ;
        RECT 393.370 855.480 393.690 855.540 ;
        RECT 328.050 46.140 328.370 46.200 ;
        RECT 1221.830 46.140 1222.150 46.200 ;
        RECT 328.050 46.000 1222.150 46.140 ;
        RECT 328.050 45.940 328.370 46.000 ;
        RECT 1221.830 45.940 1222.150 46.000 ;
      LAYER via ;
        RECT 328.080 855.480 328.340 855.740 ;
        RECT 393.400 855.480 393.660 855.740 ;
        RECT 328.080 45.940 328.340 46.200 ;
        RECT 1221.860 45.940 1222.120 46.200 ;
      LAYER met2 ;
        RECT 393.390 861.035 393.670 861.405 ;
        RECT 393.460 855.770 393.600 861.035 ;
        RECT 328.080 855.450 328.340 855.770 ;
        RECT 393.400 855.450 393.660 855.770 ;
        RECT 328.140 46.230 328.280 855.450 ;
        RECT 328.080 45.910 328.340 46.230 ;
        RECT 1221.860 45.910 1222.120 46.230 ;
        RECT 1221.920 2.400 1222.060 45.910 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
      LAYER via2 ;
        RECT 393.390 861.080 393.670 861.360 ;
      LAYER met3 ;
        RECT 393.365 861.370 393.695 861.385 ;
        RECT 410.000 861.370 414.000 861.520 ;
        RECT 393.365 861.070 414.000 861.370 ;
        RECT 393.365 861.055 393.695 861.070 ;
        RECT 410.000 860.920 414.000 861.070 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1239.770 2.960 1240.090 3.020 ;
        RECT 1241.610 2.960 1241.930 3.020 ;
        RECT 1239.770 2.820 1241.930 2.960 ;
        RECT 1239.770 2.760 1240.090 2.820 ;
        RECT 1241.610 2.760 1241.930 2.820 ;
      LAYER via ;
        RECT 1239.800 2.760 1240.060 3.020 ;
        RECT 1241.640 2.760 1241.900 3.020 ;
      LAYER met2 ;
        RECT 1241.630 361.915 1241.910 362.285 ;
        RECT 1241.700 3.050 1241.840 361.915 ;
        RECT 1239.800 2.730 1240.060 3.050 ;
        RECT 1241.640 2.730 1241.900 3.050 ;
        RECT 1239.860 2.400 1240.000 2.730 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1241.630 361.960 1241.910 362.240 ;
      LAYER met3 ;
        RECT 2506.000 2402.250 2510.000 2402.400 ;
        RECT 2529.350 2402.250 2529.730 2402.260 ;
        RECT 2506.000 2401.950 2529.730 2402.250 ;
        RECT 2506.000 2401.800 2510.000 2401.950 ;
        RECT 2529.350 2401.940 2529.730 2401.950 ;
        RECT 1241.605 362.250 1241.935 362.265 ;
        RECT 2529.350 362.250 2529.730 362.260 ;
        RECT 1241.605 361.950 2529.730 362.250 ;
        RECT 1241.605 361.935 1241.935 361.950 ;
        RECT 2529.350 361.940 2529.730 361.950 ;
      LAYER via3 ;
        RECT 2529.380 2401.940 2529.700 2402.260 ;
        RECT 2529.380 361.940 2529.700 362.260 ;
      LAYER met4 ;
        RECT 2529.375 2401.935 2529.705 2402.265 ;
        RECT 2529.390 362.265 2529.690 2401.935 ;
        RECT 2529.375 361.935 2529.705 362.265 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1269.745 16.745 1269.915 18.275 ;
      LAYER mcon ;
        RECT 1269.745 18.105 1269.915 18.275 ;
      LAYER met1 ;
        RECT 1877.330 3043.240 1877.650 3043.300 ;
        RECT 2601.830 3043.240 2602.150 3043.300 ;
        RECT 1877.330 3043.100 2602.150 3043.240 ;
        RECT 1877.330 3043.040 1877.650 3043.100 ;
        RECT 2601.830 3043.040 2602.150 3043.100 ;
        RECT 1269.685 18.260 1269.975 18.305 ;
        RECT 2601.830 18.260 2602.150 18.320 ;
        RECT 1269.685 18.120 2602.150 18.260 ;
        RECT 1269.685 18.075 1269.975 18.120 ;
        RECT 2601.830 18.060 2602.150 18.120 ;
        RECT 1257.250 16.900 1257.570 16.960 ;
        RECT 1269.685 16.900 1269.975 16.945 ;
        RECT 1257.250 16.760 1269.975 16.900 ;
        RECT 1257.250 16.700 1257.570 16.760 ;
        RECT 1269.685 16.715 1269.975 16.760 ;
      LAYER via ;
        RECT 1877.360 3043.040 1877.620 3043.300 ;
        RECT 2601.860 3043.040 2602.120 3043.300 ;
        RECT 2601.860 18.060 2602.120 18.320 ;
        RECT 1257.280 16.700 1257.540 16.960 ;
      LAYER met2 ;
        RECT 1877.360 3043.010 1877.620 3043.330 ;
        RECT 2601.860 3043.010 2602.120 3043.330 ;
        RECT 1877.420 3010.000 1877.560 3043.010 ;
        RECT 1877.420 3009.340 1877.770 3010.000 ;
        RECT 1877.490 3006.000 1877.770 3009.340 ;
        RECT 2601.920 18.350 2602.060 3043.010 ;
        RECT 2601.860 18.030 2602.120 18.350 ;
        RECT 1257.280 16.670 1257.540 16.990 ;
        RECT 1257.340 2.400 1257.480 16.670 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 385.550 2500.260 385.870 2500.320 ;
        RECT 395.210 2500.260 395.530 2500.320 ;
        RECT 385.550 2500.120 395.530 2500.260 ;
        RECT 385.550 2500.060 385.870 2500.120 ;
        RECT 395.210 2500.060 395.530 2500.120 ;
        RECT 385.550 52.260 385.870 52.320 ;
        RECT 1269.670 52.260 1269.990 52.320 ;
        RECT 385.550 52.120 1269.990 52.260 ;
        RECT 385.550 52.060 385.870 52.120 ;
        RECT 1269.670 52.060 1269.990 52.120 ;
      LAYER via ;
        RECT 385.580 2500.060 385.840 2500.320 ;
        RECT 395.240 2500.060 395.500 2500.320 ;
        RECT 385.580 52.060 385.840 52.320 ;
        RECT 1269.700 52.060 1269.960 52.320 ;
      LAYER met2 ;
        RECT 395.230 2503.915 395.510 2504.285 ;
        RECT 395.300 2500.350 395.440 2503.915 ;
        RECT 385.580 2500.030 385.840 2500.350 ;
        RECT 395.240 2500.030 395.500 2500.350 ;
        RECT 385.640 52.350 385.780 2500.030 ;
        RECT 385.580 52.030 385.840 52.350 ;
        RECT 1269.700 52.030 1269.960 52.350 ;
        RECT 1269.760 17.410 1269.900 52.030 ;
        RECT 1269.760 17.270 1275.420 17.410 ;
        RECT 1275.280 2.400 1275.420 17.270 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 395.230 2503.960 395.510 2504.240 ;
      LAYER met3 ;
        RECT 395.205 2504.250 395.535 2504.265 ;
        RECT 410.000 2504.250 414.000 2504.400 ;
        RECT 395.205 2503.950 414.000 2504.250 ;
        RECT 395.205 2503.935 395.535 2503.950 ;
        RECT 410.000 2503.800 414.000 2503.950 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 336.790 2808.640 337.110 2808.700 ;
        RECT 393.370 2808.640 393.690 2808.700 ;
        RECT 336.790 2808.500 393.690 2808.640 ;
        RECT 336.790 2808.440 337.110 2808.500 ;
        RECT 393.370 2808.440 393.690 2808.500 ;
        RECT 336.790 32.540 337.110 32.600 ;
        RECT 1293.130 32.540 1293.450 32.600 ;
        RECT 336.790 32.400 1293.450 32.540 ;
        RECT 336.790 32.340 337.110 32.400 ;
        RECT 1293.130 32.340 1293.450 32.400 ;
      LAYER via ;
        RECT 336.820 2808.440 337.080 2808.700 ;
        RECT 393.400 2808.440 393.660 2808.700 ;
        RECT 336.820 32.340 337.080 32.600 ;
        RECT 1293.160 32.340 1293.420 32.600 ;
      LAYER met2 ;
        RECT 393.390 2813.995 393.670 2814.365 ;
        RECT 393.460 2808.730 393.600 2813.995 ;
        RECT 336.820 2808.410 337.080 2808.730 ;
        RECT 393.400 2808.410 393.660 2808.730 ;
        RECT 336.880 32.630 337.020 2808.410 ;
        RECT 336.820 32.310 337.080 32.630 ;
        RECT 1293.160 32.310 1293.420 32.630 ;
        RECT 1293.220 2.400 1293.360 32.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
      LAYER via2 ;
        RECT 393.390 2814.040 393.670 2814.320 ;
      LAYER met3 ;
        RECT 393.365 2814.330 393.695 2814.345 ;
        RECT 410.000 2814.330 414.000 2814.480 ;
        RECT 393.365 2814.030 414.000 2814.330 ;
        RECT 393.365 2814.015 393.695 2814.030 ;
        RECT 410.000 2813.880 414.000 2814.030 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 16.900 1311.390 16.960 ;
        RECT 1317.050 16.900 1317.370 16.960 ;
        RECT 1311.070 16.760 1317.370 16.900 ;
        RECT 1311.070 16.700 1311.390 16.760 ;
        RECT 1317.050 16.700 1317.370 16.760 ;
      LAYER via ;
        RECT 1311.100 16.700 1311.360 16.960 ;
        RECT 1317.080 16.700 1317.340 16.960 ;
      LAYER met2 ;
        RECT 1317.070 431.275 1317.350 431.645 ;
        RECT 1317.140 16.990 1317.280 431.275 ;
        RECT 1311.100 16.670 1311.360 16.990 ;
        RECT 1317.080 16.670 1317.340 16.990 ;
        RECT 1311.160 2.400 1311.300 16.670 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1317.070 431.320 1317.350 431.600 ;
      LAYER met3 ;
        RECT 2506.000 2566.810 2510.000 2566.960 ;
        RECT 2528.430 2566.810 2528.810 2566.820 ;
        RECT 2506.000 2566.510 2528.810 2566.810 ;
        RECT 2506.000 2566.360 2510.000 2566.510 ;
        RECT 2528.430 2566.500 2528.810 2566.510 ;
        RECT 1317.045 431.610 1317.375 431.625 ;
        RECT 2528.430 431.610 2528.810 431.620 ;
        RECT 1317.045 431.310 2528.810 431.610 ;
        RECT 1317.045 431.295 1317.375 431.310 ;
        RECT 2528.430 431.300 2528.810 431.310 ;
      LAYER via3 ;
        RECT 2528.460 2566.500 2528.780 2566.820 ;
        RECT 2528.460 431.300 2528.780 431.620 ;
      LAYER met4 ;
        RECT 2528.455 2566.495 2528.785 2566.825 ;
        RECT 2528.470 431.625 2528.770 2566.495 ;
        RECT 2528.455 431.295 2528.785 431.625 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2508.010 1606.995 2508.290 1607.365 ;
        RECT 2508.080 1560.445 2508.220 1606.995 ;
        RECT 2508.010 1560.075 2508.290 1560.445 ;
        RECT 1330.870 355.795 1331.150 356.165 ;
        RECT 1330.940 17.410 1331.080 355.795 ;
        RECT 1329.100 17.270 1331.080 17.410 ;
        RECT 1329.100 2.400 1329.240 17.270 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 2508.010 1607.040 2508.290 1607.320 ;
        RECT 2508.010 1560.120 2508.290 1560.400 ;
        RECT 1330.870 355.840 1331.150 356.120 ;
      LAYER met3 ;
        RECT 2506.000 2293.000 2510.000 2293.600 ;
        RECT 2508.230 2291.420 2508.530 2293.000 ;
        RECT 2508.190 2291.100 2508.570 2291.420 ;
        RECT 2507.270 1608.380 2507.650 1608.700 ;
        RECT 2507.310 1607.330 2507.610 1608.380 ;
        RECT 2507.985 1607.330 2508.315 1607.345 ;
        RECT 2507.310 1607.030 2508.315 1607.330 ;
        RECT 2507.985 1607.015 2508.315 1607.030 ;
        RECT 2507.985 1560.410 2508.315 1560.425 ;
        RECT 2507.310 1560.110 2508.315 1560.410 ;
        RECT 2507.310 1559.740 2507.610 1560.110 ;
        RECT 2507.985 1560.095 2508.315 1560.110 ;
        RECT 2507.270 1559.420 2507.650 1559.740 ;
        RECT 2506.350 1280.250 2506.730 1280.260 ;
        RECT 2507.270 1280.250 2507.650 1280.260 ;
        RECT 2506.350 1279.950 2507.650 1280.250 ;
        RECT 2506.350 1279.940 2506.730 1279.950 ;
        RECT 2507.270 1279.940 2507.650 1279.950 ;
        RECT 2507.270 1145.980 2507.650 1146.300 ;
        RECT 2507.310 1144.940 2507.610 1145.980 ;
        RECT 2507.270 1144.620 2507.650 1144.940 ;
        RECT 2506.350 1098.010 2506.730 1098.020 ;
        RECT 2506.350 1097.710 2507.610 1098.010 ;
        RECT 2506.350 1097.700 2506.730 1097.710 ;
        RECT 2507.310 1097.340 2507.610 1097.710 ;
        RECT 2507.270 1097.020 2507.650 1097.340 ;
        RECT 2507.270 607.730 2507.650 607.740 ;
        RECT 2507.270 607.430 2508.530 607.730 ;
        RECT 2507.270 607.420 2507.650 607.430 ;
        RECT 2508.230 606.380 2508.530 607.430 ;
        RECT 2508.190 606.060 2508.570 606.380 ;
        RECT 1330.845 356.130 1331.175 356.145 ;
        RECT 2508.190 356.130 2508.570 356.140 ;
        RECT 1330.845 355.830 2508.570 356.130 ;
        RECT 1330.845 355.815 1331.175 355.830 ;
        RECT 2508.190 355.820 2508.570 355.830 ;
      LAYER via3 ;
        RECT 2508.220 2291.100 2508.540 2291.420 ;
        RECT 2507.300 1608.380 2507.620 1608.700 ;
        RECT 2507.300 1559.420 2507.620 1559.740 ;
        RECT 2506.380 1279.940 2506.700 1280.260 ;
        RECT 2507.300 1279.940 2507.620 1280.260 ;
        RECT 2507.300 1145.980 2507.620 1146.300 ;
        RECT 2507.300 1144.620 2507.620 1144.940 ;
        RECT 2506.380 1097.700 2506.700 1098.020 ;
        RECT 2507.300 1097.020 2507.620 1097.340 ;
        RECT 2507.300 607.420 2507.620 607.740 ;
        RECT 2508.220 606.060 2508.540 606.380 ;
        RECT 2508.220 355.820 2508.540 356.140 ;
      LAYER met4 ;
        RECT 2508.215 2291.095 2508.545 2291.425 ;
        RECT 2508.230 2222.050 2508.530 2291.095 ;
        RECT 2506.390 2221.750 2508.530 2222.050 ;
        RECT 2506.390 2058.850 2506.690 2221.750 ;
        RECT 2506.390 2058.550 2508.530 2058.850 ;
        RECT 2508.230 2007.850 2508.530 2058.550 ;
        RECT 2507.310 2007.550 2508.530 2007.850 ;
        RECT 2507.310 1984.050 2507.610 2007.550 ;
        RECT 2506.390 1983.750 2507.610 1984.050 ;
        RECT 2506.390 1912.650 2506.690 1983.750 ;
        RECT 2505.470 1912.350 2506.690 1912.650 ;
        RECT 2505.470 1817.450 2505.770 1912.350 ;
        RECT 2505.470 1817.150 2506.690 1817.450 ;
        RECT 2506.390 1712.050 2506.690 1817.150 ;
        RECT 2506.390 1711.750 2507.610 1712.050 ;
        RECT 2507.310 1608.705 2507.610 1711.750 ;
        RECT 2507.295 1608.375 2507.625 1608.705 ;
        RECT 2507.295 1559.415 2507.625 1559.745 ;
        RECT 2507.310 1440.050 2507.610 1559.415 ;
        RECT 2504.550 1439.750 2507.610 1440.050 ;
        RECT 2504.550 1280.250 2504.850 1439.750 ;
        RECT 2506.375 1280.250 2506.705 1280.265 ;
        RECT 2504.550 1279.950 2506.705 1280.250 ;
        RECT 2506.375 1279.935 2506.705 1279.950 ;
        RECT 2507.295 1279.935 2507.625 1280.265 ;
        RECT 2507.310 1146.305 2507.610 1279.935 ;
        RECT 2507.295 1145.975 2507.625 1146.305 ;
        RECT 2507.295 1144.615 2507.625 1144.945 ;
        RECT 2507.310 1144.250 2507.610 1144.615 ;
        RECT 2506.390 1143.950 2507.610 1144.250 ;
        RECT 2506.390 1098.025 2506.690 1143.950 ;
        RECT 2506.375 1097.695 2506.705 1098.025 ;
        RECT 2507.295 1097.015 2507.625 1097.345 ;
        RECT 2507.310 1049.050 2507.610 1097.015 ;
        RECT 2507.310 1048.750 2508.530 1049.050 ;
        RECT 2508.230 899.450 2508.530 1048.750 ;
        RECT 2505.470 899.150 2508.530 899.450 ;
        RECT 2505.470 896.050 2505.770 899.150 ;
        RECT 2504.550 895.750 2505.770 896.050 ;
        RECT 2504.550 637.650 2504.850 895.750 ;
        RECT 2504.550 637.350 2506.690 637.650 ;
        RECT 2506.390 634.250 2506.690 637.350 ;
        RECT 2506.390 633.950 2507.610 634.250 ;
        RECT 2507.310 607.745 2507.610 633.950 ;
        RECT 2507.295 607.415 2507.625 607.745 ;
        RECT 2508.215 606.055 2508.545 606.385 ;
        RECT 2508.230 356.145 2508.530 606.055 ;
        RECT 2508.215 355.815 2508.545 356.145 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 93.740 586.430 93.800 ;
        RECT 683.170 93.740 683.490 93.800 ;
        RECT 586.110 93.600 683.490 93.740 ;
        RECT 586.110 93.540 586.430 93.600 ;
        RECT 683.170 93.540 683.490 93.600 ;
      LAYER via ;
        RECT 586.140 93.540 586.400 93.800 ;
        RECT 683.200 93.540 683.460 93.800 ;
      LAYER met2 ;
        RECT 584.890 510.410 585.170 514.000 ;
        RECT 584.890 510.270 586.340 510.410 ;
        RECT 584.890 510.000 585.170 510.270 ;
        RECT 586.200 93.830 586.340 510.270 ;
        RECT 586.140 93.510 586.400 93.830 ;
        RECT 683.200 93.510 683.460 93.830 ;
        RECT 683.260 17.410 683.400 93.510 ;
        RECT 683.260 17.270 686.620 17.410 ;
        RECT 686.480 2.400 686.620 17.270 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 316.550 2553.300 316.870 2553.360 ;
        RECT 393.370 2553.300 393.690 2553.360 ;
        RECT 316.550 2553.160 393.690 2553.300 ;
        RECT 316.550 2553.100 316.870 2553.160 ;
        RECT 393.370 2553.100 393.690 2553.160 ;
        RECT 316.550 61.100 316.870 61.160 ;
        RECT 1345.570 61.100 1345.890 61.160 ;
        RECT 316.550 60.960 1345.890 61.100 ;
        RECT 316.550 60.900 316.870 60.960 ;
        RECT 1345.570 60.900 1345.890 60.960 ;
      LAYER via ;
        RECT 316.580 2553.100 316.840 2553.360 ;
        RECT 393.400 2553.100 393.660 2553.360 ;
        RECT 316.580 60.900 316.840 61.160 ;
        RECT 1345.600 60.900 1345.860 61.160 ;
      LAYER met2 ;
        RECT 393.390 2558.315 393.670 2558.685 ;
        RECT 393.460 2553.390 393.600 2558.315 ;
        RECT 316.580 2553.070 316.840 2553.390 ;
        RECT 393.400 2553.070 393.660 2553.390 ;
        RECT 316.640 61.190 316.780 2553.070 ;
        RECT 316.580 60.870 316.840 61.190 ;
        RECT 1345.600 60.870 1345.860 61.190 ;
        RECT 1345.660 17.410 1345.800 60.870 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 393.390 2558.360 393.670 2558.640 ;
      LAYER met3 ;
        RECT 393.365 2558.650 393.695 2558.665 ;
        RECT 410.000 2558.650 414.000 2558.800 ;
        RECT 393.365 2558.350 414.000 2558.650 ;
        RECT 393.365 2558.335 393.695 2558.350 ;
        RECT 410.000 2558.200 414.000 2558.350 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1704.370 3036.100 1704.690 3036.160 ;
        RECT 2528.690 3036.100 2529.010 3036.160 ;
        RECT 1704.370 3035.960 2529.010 3036.100 ;
        RECT 1704.370 3035.900 1704.690 3035.960 ;
        RECT 2528.690 3035.900 2529.010 3035.960 ;
        RECT 2528.690 1776.740 2529.010 1776.800 ;
        RECT 2598.150 1776.740 2598.470 1776.800 ;
        RECT 2528.690 1776.600 2598.470 1776.740 ;
        RECT 2528.690 1776.540 2529.010 1776.600 ;
        RECT 2598.150 1776.540 2598.470 1776.600 ;
        RECT 2598.150 1157.260 2598.470 1157.320 ;
        RECT 2604.590 1157.260 2604.910 1157.320 ;
        RECT 2598.150 1157.120 2604.910 1157.260 ;
        RECT 2598.150 1157.060 2598.470 1157.120 ;
        RECT 2604.590 1157.060 2604.910 1157.120 ;
        RECT 2566.410 503.780 2566.730 503.840 ;
        RECT 2604.590 503.780 2604.910 503.840 ;
        RECT 2566.410 503.640 2604.910 503.780 ;
        RECT 2566.410 503.580 2566.730 503.640 ;
        RECT 2604.590 503.580 2604.910 503.640 ;
        RECT 2515.350 496.640 2515.670 496.700 ;
        RECT 2566.410 496.640 2566.730 496.700 ;
        RECT 2515.350 496.500 2566.730 496.640 ;
        RECT 2515.350 496.440 2515.670 496.500 ;
        RECT 2566.410 496.440 2566.730 496.500 ;
        RECT 2456.470 488.140 2456.790 488.200 ;
        RECT 2515.350 488.140 2515.670 488.200 ;
        RECT 2456.470 488.000 2515.670 488.140 ;
        RECT 2456.470 487.940 2456.790 488.000 ;
        RECT 2515.350 487.940 2515.670 488.000 ;
        RECT 2438.990 469.440 2439.310 469.500 ;
        RECT 2456.470 469.440 2456.790 469.500 ;
        RECT 2438.990 469.300 2456.790 469.440 ;
        RECT 2438.990 469.240 2439.310 469.300 ;
        RECT 2456.470 469.240 2456.790 469.300 ;
        RECT 2422.430 443.260 2422.750 443.320 ;
        RECT 2438.990 443.260 2439.310 443.320 ;
        RECT 2422.430 443.120 2439.310 443.260 ;
        RECT 2422.430 443.060 2422.750 443.120 ;
        RECT 2438.990 443.060 2439.310 443.120 ;
        RECT 2418.750 434.760 2419.070 434.820 ;
        RECT 2422.430 434.760 2422.750 434.820 ;
        RECT 2418.750 434.620 2422.750 434.760 ;
        RECT 2418.750 434.560 2419.070 434.620 ;
        RECT 2422.430 434.560 2422.750 434.620 ;
        RECT 2405.410 414.360 2405.730 414.420 ;
        RECT 2418.750 414.360 2419.070 414.420 ;
        RECT 2405.410 414.220 2419.070 414.360 ;
        RECT 2405.410 414.160 2405.730 414.220 ;
        RECT 2418.750 414.160 2419.070 414.220 ;
        RECT 2394.370 407.220 2394.690 407.280 ;
        RECT 2405.410 407.220 2405.730 407.280 ;
        RECT 2394.370 407.080 2405.730 407.220 ;
        RECT 2394.370 407.020 2394.690 407.080 ;
        RECT 2405.410 407.020 2405.730 407.080 ;
        RECT 2376.890 387.840 2377.210 387.900 ;
        RECT 2394.370 387.840 2394.690 387.900 ;
        RECT 2376.890 387.700 2394.690 387.840 ;
        RECT 2376.890 387.640 2377.210 387.700 ;
        RECT 2394.370 387.640 2394.690 387.700 ;
        RECT 2362.170 353.160 2362.490 353.220 ;
        RECT 2376.890 353.160 2377.210 353.220 ;
        RECT 2362.170 353.020 2377.210 353.160 ;
        RECT 2362.170 352.960 2362.490 353.020 ;
        RECT 2376.890 352.960 2377.210 353.020 ;
        RECT 2349.290 346.360 2349.610 346.420 ;
        RECT 2362.170 346.360 2362.490 346.420 ;
        RECT 2349.290 346.220 2362.490 346.360 ;
        RECT 2349.290 346.160 2349.610 346.220 ;
        RECT 2362.170 346.160 2362.490 346.220 ;
        RECT 2339.170 288.900 2339.490 288.960 ;
        RECT 2349.290 288.900 2349.610 288.960 ;
        RECT 2339.170 288.760 2349.610 288.900 ;
        RECT 2339.170 288.700 2339.490 288.760 ;
        RECT 2349.290 288.700 2349.610 288.760 ;
        RECT 2321.690 269.180 2322.010 269.240 ;
        RECT 2339.170 269.180 2339.490 269.240 ;
        RECT 2321.690 269.040 2339.490 269.180 ;
        RECT 2321.690 268.980 2322.010 269.040 ;
        RECT 2339.170 268.980 2339.490 269.040 ;
        RECT 2313.410 217.840 2313.730 217.900 ;
        RECT 2321.690 217.840 2322.010 217.900 ;
        RECT 2313.410 217.700 2322.010 217.840 ;
        RECT 2313.410 217.640 2313.730 217.700 ;
        RECT 2321.690 217.640 2322.010 217.700 ;
        RECT 2300.990 207.300 2301.310 207.360 ;
        RECT 2313.410 207.300 2313.730 207.360 ;
        RECT 2300.990 207.160 2313.730 207.300 ;
        RECT 2300.990 207.100 2301.310 207.160 ;
        RECT 2313.410 207.100 2313.730 207.160 ;
        RECT 1364.430 24.040 1364.750 24.100 ;
        RECT 2300.990 24.040 2301.310 24.100 ;
        RECT 1364.430 23.900 2301.310 24.040 ;
        RECT 1364.430 23.840 1364.750 23.900 ;
        RECT 2300.990 23.840 2301.310 23.900 ;
      LAYER via ;
        RECT 1704.400 3035.900 1704.660 3036.160 ;
        RECT 2528.720 3035.900 2528.980 3036.160 ;
        RECT 2528.720 1776.540 2528.980 1776.800 ;
        RECT 2598.180 1776.540 2598.440 1776.800 ;
        RECT 2598.180 1157.060 2598.440 1157.320 ;
        RECT 2604.620 1157.060 2604.880 1157.320 ;
        RECT 2566.440 503.580 2566.700 503.840 ;
        RECT 2604.620 503.580 2604.880 503.840 ;
        RECT 2515.380 496.440 2515.640 496.700 ;
        RECT 2566.440 496.440 2566.700 496.700 ;
        RECT 2456.500 487.940 2456.760 488.200 ;
        RECT 2515.380 487.940 2515.640 488.200 ;
        RECT 2439.020 469.240 2439.280 469.500 ;
        RECT 2456.500 469.240 2456.760 469.500 ;
        RECT 2422.460 443.060 2422.720 443.320 ;
        RECT 2439.020 443.060 2439.280 443.320 ;
        RECT 2418.780 434.560 2419.040 434.820 ;
        RECT 2422.460 434.560 2422.720 434.820 ;
        RECT 2405.440 414.160 2405.700 414.420 ;
        RECT 2418.780 414.160 2419.040 414.420 ;
        RECT 2394.400 407.020 2394.660 407.280 ;
        RECT 2405.440 407.020 2405.700 407.280 ;
        RECT 2376.920 387.640 2377.180 387.900 ;
        RECT 2394.400 387.640 2394.660 387.900 ;
        RECT 2362.200 352.960 2362.460 353.220 ;
        RECT 2376.920 352.960 2377.180 353.220 ;
        RECT 2349.320 346.160 2349.580 346.420 ;
        RECT 2362.200 346.160 2362.460 346.420 ;
        RECT 2339.200 288.700 2339.460 288.960 ;
        RECT 2349.320 288.700 2349.580 288.960 ;
        RECT 2321.720 268.980 2321.980 269.240 ;
        RECT 2339.200 268.980 2339.460 269.240 ;
        RECT 2313.440 217.640 2313.700 217.900 ;
        RECT 2321.720 217.640 2321.980 217.900 ;
        RECT 2301.020 207.100 2301.280 207.360 ;
        RECT 2313.440 207.100 2313.700 207.360 ;
        RECT 1364.460 23.840 1364.720 24.100 ;
        RECT 2301.020 23.840 2301.280 24.100 ;
      LAYER met2 ;
        RECT 1704.400 3035.870 1704.660 3036.190 ;
        RECT 2528.720 3035.870 2528.980 3036.190 ;
        RECT 1704.460 3010.000 1704.600 3035.870 ;
        RECT 1704.460 3009.340 1704.810 3010.000 ;
        RECT 1704.530 3006.000 1704.810 3009.340 ;
        RECT 2528.780 1776.830 2528.920 3035.870 ;
        RECT 2528.720 1776.510 2528.980 1776.830 ;
        RECT 2598.180 1776.510 2598.440 1776.830 ;
        RECT 2598.240 1157.350 2598.380 1776.510 ;
        RECT 2598.180 1157.030 2598.440 1157.350 ;
        RECT 2604.620 1157.030 2604.880 1157.350 ;
        RECT 2604.680 503.870 2604.820 1157.030 ;
        RECT 2566.440 503.550 2566.700 503.870 ;
        RECT 2604.620 503.550 2604.880 503.870 ;
        RECT 2566.500 496.730 2566.640 503.550 ;
        RECT 2515.380 496.410 2515.640 496.730 ;
        RECT 2566.440 496.410 2566.700 496.730 ;
        RECT 2515.440 488.230 2515.580 496.410 ;
        RECT 2456.500 487.910 2456.760 488.230 ;
        RECT 2515.380 487.910 2515.640 488.230 ;
        RECT 2456.560 469.530 2456.700 487.910 ;
        RECT 2439.020 469.210 2439.280 469.530 ;
        RECT 2456.500 469.210 2456.760 469.530 ;
        RECT 2439.080 443.350 2439.220 469.210 ;
        RECT 2422.460 443.030 2422.720 443.350 ;
        RECT 2439.020 443.030 2439.280 443.350 ;
        RECT 2422.520 434.850 2422.660 443.030 ;
        RECT 2418.780 434.530 2419.040 434.850 ;
        RECT 2422.460 434.530 2422.720 434.850 ;
        RECT 2418.840 414.450 2418.980 434.530 ;
        RECT 2405.440 414.130 2405.700 414.450 ;
        RECT 2418.780 414.130 2419.040 414.450 ;
        RECT 2405.500 407.310 2405.640 414.130 ;
        RECT 2394.400 406.990 2394.660 407.310 ;
        RECT 2405.440 406.990 2405.700 407.310 ;
        RECT 2394.460 387.930 2394.600 406.990 ;
        RECT 2376.920 387.610 2377.180 387.930 ;
        RECT 2394.400 387.610 2394.660 387.930 ;
        RECT 2376.980 353.250 2377.120 387.610 ;
        RECT 2362.200 352.930 2362.460 353.250 ;
        RECT 2376.920 352.930 2377.180 353.250 ;
        RECT 2362.260 346.450 2362.400 352.930 ;
        RECT 2349.320 346.130 2349.580 346.450 ;
        RECT 2362.200 346.130 2362.460 346.450 ;
        RECT 2349.380 288.990 2349.520 346.130 ;
        RECT 2339.200 288.670 2339.460 288.990 ;
        RECT 2349.320 288.670 2349.580 288.990 ;
        RECT 2339.260 269.270 2339.400 288.670 ;
        RECT 2321.720 268.950 2321.980 269.270 ;
        RECT 2339.200 268.950 2339.460 269.270 ;
        RECT 2321.780 217.930 2321.920 268.950 ;
        RECT 2313.440 217.610 2313.700 217.930 ;
        RECT 2321.720 217.610 2321.980 217.930 ;
        RECT 2313.500 207.390 2313.640 217.610 ;
        RECT 2301.020 207.070 2301.280 207.390 ;
        RECT 2313.440 207.070 2313.700 207.390 ;
        RECT 2301.080 24.130 2301.220 207.070 ;
        RECT 1364.460 23.810 1364.720 24.130 ;
        RECT 2301.020 23.810 2301.280 24.130 ;
        RECT 1364.520 2.400 1364.660 23.810 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 342.310 766.260 342.630 766.320 ;
        RECT 393.370 766.260 393.690 766.320 ;
        RECT 342.310 766.120 393.690 766.260 ;
        RECT 342.310 766.060 342.630 766.120 ;
        RECT 393.370 766.060 393.690 766.120 ;
        RECT 342.310 60.760 342.630 60.820 ;
        RECT 1382.370 60.760 1382.690 60.820 ;
        RECT 342.310 60.620 1382.690 60.760 ;
        RECT 342.310 60.560 342.630 60.620 ;
        RECT 1382.370 60.560 1382.690 60.620 ;
      LAYER via ;
        RECT 342.340 766.060 342.600 766.320 ;
        RECT 393.400 766.060 393.660 766.320 ;
        RECT 342.340 60.560 342.600 60.820 ;
        RECT 1382.400 60.560 1382.660 60.820 ;
      LAYER met2 ;
        RECT 393.390 768.555 393.670 768.925 ;
        RECT 393.460 766.350 393.600 768.555 ;
        RECT 342.340 766.030 342.600 766.350 ;
        RECT 393.400 766.030 393.660 766.350 ;
        RECT 342.400 60.850 342.540 766.030 ;
        RECT 342.340 60.530 342.600 60.850 ;
        RECT 1382.400 60.530 1382.660 60.850 ;
        RECT 1382.460 2.400 1382.600 60.530 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 393.390 768.600 393.670 768.880 ;
      LAYER met3 ;
        RECT 393.365 768.890 393.695 768.905 ;
        RECT 410.000 768.890 414.000 769.040 ;
        RECT 393.365 768.590 414.000 768.890 ;
        RECT 393.365 768.575 393.695 768.590 ;
        RECT 410.000 768.440 414.000 768.590 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.010 2773.960 317.330 2774.020 ;
        RECT 393.370 2773.960 393.690 2774.020 ;
        RECT 317.010 2773.820 393.690 2773.960 ;
        RECT 317.010 2773.760 317.330 2773.820 ;
        RECT 393.370 2773.760 393.690 2773.820 ;
        RECT 317.010 47.160 317.330 47.220 ;
        RECT 1399.850 47.160 1400.170 47.220 ;
        RECT 317.010 47.020 1400.170 47.160 ;
        RECT 317.010 46.960 317.330 47.020 ;
        RECT 1399.850 46.960 1400.170 47.020 ;
      LAYER via ;
        RECT 317.040 2773.760 317.300 2774.020 ;
        RECT 393.400 2773.760 393.660 2774.020 ;
        RECT 317.040 46.960 317.300 47.220 ;
        RECT 1399.880 46.960 1400.140 47.220 ;
      LAYER met2 ;
        RECT 393.390 2778.635 393.670 2779.005 ;
        RECT 393.460 2774.050 393.600 2778.635 ;
        RECT 317.040 2773.730 317.300 2774.050 ;
        RECT 393.400 2773.730 393.660 2774.050 ;
        RECT 317.100 47.250 317.240 2773.730 ;
        RECT 317.040 46.930 317.300 47.250 ;
        RECT 1399.880 46.930 1400.140 47.250 ;
        RECT 1399.940 19.450 1400.080 46.930 ;
        RECT 1399.940 19.310 1400.540 19.450 ;
        RECT 1400.400 2.400 1400.540 19.310 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 393.390 2778.680 393.670 2778.960 ;
      LAYER met3 ;
        RECT 393.365 2778.970 393.695 2778.985 ;
        RECT 410.000 2778.970 414.000 2779.120 ;
        RECT 393.365 2778.670 414.000 2778.970 ;
        RECT 393.365 2778.655 393.695 2778.670 ;
        RECT 410.000 2778.520 414.000 2778.670 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1049.140 2520.730 1049.200 ;
        RECT 2562.730 1049.140 2563.050 1049.200 ;
        RECT 2520.410 1049.000 2563.050 1049.140 ;
        RECT 2520.410 1048.940 2520.730 1049.000 ;
        RECT 2562.730 1048.940 2563.050 1049.000 ;
        RECT 1421.010 494.600 1421.330 494.660 ;
        RECT 2562.730 494.600 2563.050 494.660 ;
        RECT 1421.010 494.460 2563.050 494.600 ;
        RECT 1421.010 494.400 1421.330 494.460 ;
        RECT 2562.730 494.400 2563.050 494.460 ;
        RECT 1418.250 16.900 1418.570 16.960 ;
        RECT 1421.010 16.900 1421.330 16.960 ;
        RECT 1418.250 16.760 1421.330 16.900 ;
        RECT 1418.250 16.700 1418.570 16.760 ;
        RECT 1421.010 16.700 1421.330 16.760 ;
      LAYER via ;
        RECT 2520.440 1048.940 2520.700 1049.200 ;
        RECT 2562.760 1048.940 2563.020 1049.200 ;
        RECT 1421.040 494.400 1421.300 494.660 ;
        RECT 2562.760 494.400 2563.020 494.660 ;
        RECT 1418.280 16.700 1418.540 16.960 ;
        RECT 1421.040 16.700 1421.300 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1051.435 2520.710 1051.805 ;
        RECT 2520.500 1049.230 2520.640 1051.435 ;
        RECT 2520.440 1048.910 2520.700 1049.230 ;
        RECT 2562.760 1048.910 2563.020 1049.230 ;
        RECT 2562.820 494.690 2562.960 1048.910 ;
        RECT 1421.040 494.370 1421.300 494.690 ;
        RECT 2562.760 494.370 2563.020 494.690 ;
        RECT 1421.100 16.990 1421.240 494.370 ;
        RECT 1418.280 16.670 1418.540 16.990 ;
        RECT 1421.040 16.670 1421.300 16.990 ;
        RECT 1418.340 2.400 1418.480 16.670 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1051.480 2520.710 1051.760 ;
      LAYER met3 ;
        RECT 2506.000 1051.770 2510.000 1051.920 ;
        RECT 2520.405 1051.770 2520.735 1051.785 ;
        RECT 2506.000 1051.470 2520.735 1051.770 ;
        RECT 2506.000 1051.320 2510.000 1051.470 ;
        RECT 2520.405 1051.455 2520.735 1051.470 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1729.210 3019.780 1729.530 3019.840 ;
        RECT 2463.370 3019.780 2463.690 3019.840 ;
        RECT 1729.210 3019.640 2463.690 3019.780 ;
        RECT 1729.210 3019.580 1729.530 3019.640 ;
        RECT 2463.370 3019.580 2463.690 3019.640 ;
        RECT 2463.370 3014.000 2463.690 3014.060 ;
        RECT 2490.970 3014.000 2491.290 3014.060 ;
        RECT 2463.370 3013.860 2491.290 3014.000 ;
        RECT 2463.370 3013.800 2463.690 3013.860 ;
        RECT 2490.970 3013.800 2491.290 3013.860 ;
        RECT 2490.970 3006.520 2491.290 3006.580 ;
        RECT 2519.950 3006.520 2520.270 3006.580 ;
        RECT 2490.970 3006.380 2520.270 3006.520 ;
        RECT 2490.970 3006.320 2491.290 3006.380 ;
        RECT 2519.950 3006.320 2520.270 3006.380 ;
        RECT 2519.950 2991.560 2520.270 2991.620 ;
        RECT 2615.630 2991.560 2615.950 2991.620 ;
        RECT 2519.950 2991.420 2615.950 2991.560 ;
        RECT 2519.950 2991.360 2520.270 2991.420 ;
        RECT 2615.630 2991.360 2615.950 2991.420 ;
        RECT 2463.830 473.520 2464.150 473.580 ;
        RECT 2615.630 473.520 2615.950 473.580 ;
        RECT 2463.830 473.380 2615.950 473.520 ;
        RECT 2463.830 473.320 2464.150 473.380 ;
        RECT 2615.630 473.320 2615.950 473.380 ;
        RECT 2442.670 459.920 2442.990 459.980 ;
        RECT 2463.830 459.920 2464.150 459.980 ;
        RECT 2442.670 459.780 2464.150 459.920 ;
        RECT 2442.670 459.720 2442.990 459.780 ;
        RECT 2463.830 459.720 2464.150 459.780 ;
        RECT 2436.230 433.400 2436.550 433.460 ;
        RECT 2442.670 433.400 2442.990 433.460 ;
        RECT 2436.230 433.260 2442.990 433.400 ;
        RECT 2436.230 433.200 2436.550 433.260 ;
        RECT 2442.670 433.200 2442.990 433.260 ;
        RECT 2427.490 414.360 2427.810 414.420 ;
        RECT 2436.230 414.360 2436.550 414.420 ;
        RECT 2427.490 414.220 2436.550 414.360 ;
        RECT 2427.490 414.160 2427.810 414.220 ;
        RECT 2436.230 414.160 2436.550 414.220 ;
        RECT 2418.290 391.240 2418.610 391.300 ;
        RECT 2427.490 391.240 2427.810 391.300 ;
        RECT 2418.290 391.100 2427.810 391.240 ;
        RECT 2418.290 391.040 2418.610 391.100 ;
        RECT 2427.490 391.040 2427.810 391.100 ;
        RECT 2410.010 303.860 2410.330 303.920 ;
        RECT 2418.290 303.860 2418.610 303.920 ;
        RECT 2410.010 303.720 2418.610 303.860 ;
        RECT 2410.010 303.660 2410.330 303.720 ;
        RECT 2418.290 303.660 2418.610 303.720 ;
        RECT 2394.370 280.060 2394.690 280.120 ;
        RECT 2410.010 280.060 2410.330 280.120 ;
        RECT 2394.370 279.920 2410.330 280.060 ;
        RECT 2394.370 279.860 2394.690 279.920 ;
        RECT 2410.010 279.860 2410.330 279.920 ;
        RECT 2364.470 269.520 2364.790 269.580 ;
        RECT 2394.370 269.520 2394.690 269.580 ;
        RECT 2364.470 269.380 2394.690 269.520 ;
        RECT 2364.470 269.320 2364.790 269.380 ;
        RECT 2394.370 269.320 2394.690 269.380 ;
        RECT 2339.170 262.380 2339.490 262.440 ;
        RECT 2364.470 262.380 2364.790 262.440 ;
        RECT 2339.170 262.240 2364.790 262.380 ;
        RECT 2339.170 262.180 2339.490 262.240 ;
        RECT 2364.470 262.180 2364.790 262.240 ;
        RECT 2329.050 239.600 2329.370 239.660 ;
        RECT 2339.170 239.600 2339.490 239.660 ;
        RECT 2329.050 239.460 2339.490 239.600 ;
        RECT 2329.050 239.400 2329.370 239.460 ;
        RECT 2339.170 239.400 2339.490 239.460 ;
        RECT 2318.930 214.100 2319.250 214.160 ;
        RECT 2329.050 214.100 2329.370 214.160 ;
        RECT 2318.930 213.960 2329.370 214.100 ;
        RECT 2318.930 213.900 2319.250 213.960 ;
        RECT 2329.050 213.900 2329.370 213.960 ;
        RECT 2307.890 199.480 2308.210 199.540 ;
        RECT 2318.930 199.480 2319.250 199.540 ;
        RECT 2307.890 199.340 2319.250 199.480 ;
        RECT 2307.890 199.280 2308.210 199.340 ;
        RECT 2318.930 199.280 2319.250 199.340 ;
        RECT 2291.330 172.620 2291.650 172.680 ;
        RECT 2307.890 172.620 2308.210 172.680 ;
        RECT 2291.330 172.480 2308.210 172.620 ;
        RECT 2291.330 172.420 2291.650 172.480 ;
        RECT 2307.890 172.420 2308.210 172.480 ;
        RECT 2287.190 151.200 2287.510 151.260 ;
        RECT 2291.330 151.200 2291.650 151.260 ;
        RECT 2287.190 151.060 2291.650 151.200 ;
        RECT 2287.190 151.000 2287.510 151.060 ;
        RECT 2291.330 151.000 2291.650 151.060 ;
        RECT 2277.070 110.740 2277.390 110.800 ;
        RECT 2287.190 110.740 2287.510 110.800 ;
        RECT 2277.070 110.600 2287.510 110.740 ;
        RECT 2277.070 110.540 2277.390 110.600 ;
        RECT 2287.190 110.540 2287.510 110.600 ;
        RECT 2252.690 86.940 2253.010 87.000 ;
        RECT 2276.610 86.940 2276.930 87.000 ;
        RECT 2252.690 86.800 2276.930 86.940 ;
        RECT 2252.690 86.740 2253.010 86.800 ;
        RECT 2276.610 86.740 2276.930 86.800 ;
        RECT 1435.730 24.380 1436.050 24.440 ;
        RECT 2252.690 24.380 2253.010 24.440 ;
        RECT 1435.730 24.240 2253.010 24.380 ;
        RECT 1435.730 24.180 1436.050 24.240 ;
        RECT 2252.690 24.180 2253.010 24.240 ;
      LAYER via ;
        RECT 1729.240 3019.580 1729.500 3019.840 ;
        RECT 2463.400 3019.580 2463.660 3019.840 ;
        RECT 2463.400 3013.800 2463.660 3014.060 ;
        RECT 2491.000 3013.800 2491.260 3014.060 ;
        RECT 2491.000 3006.320 2491.260 3006.580 ;
        RECT 2519.980 3006.320 2520.240 3006.580 ;
        RECT 2519.980 2991.360 2520.240 2991.620 ;
        RECT 2615.660 2991.360 2615.920 2991.620 ;
        RECT 2463.860 473.320 2464.120 473.580 ;
        RECT 2615.660 473.320 2615.920 473.580 ;
        RECT 2442.700 459.720 2442.960 459.980 ;
        RECT 2463.860 459.720 2464.120 459.980 ;
        RECT 2436.260 433.200 2436.520 433.460 ;
        RECT 2442.700 433.200 2442.960 433.460 ;
        RECT 2427.520 414.160 2427.780 414.420 ;
        RECT 2436.260 414.160 2436.520 414.420 ;
        RECT 2418.320 391.040 2418.580 391.300 ;
        RECT 2427.520 391.040 2427.780 391.300 ;
        RECT 2410.040 303.660 2410.300 303.920 ;
        RECT 2418.320 303.660 2418.580 303.920 ;
        RECT 2394.400 279.860 2394.660 280.120 ;
        RECT 2410.040 279.860 2410.300 280.120 ;
        RECT 2364.500 269.320 2364.760 269.580 ;
        RECT 2394.400 269.320 2394.660 269.580 ;
        RECT 2339.200 262.180 2339.460 262.440 ;
        RECT 2364.500 262.180 2364.760 262.440 ;
        RECT 2329.080 239.400 2329.340 239.660 ;
        RECT 2339.200 239.400 2339.460 239.660 ;
        RECT 2318.960 213.900 2319.220 214.160 ;
        RECT 2329.080 213.900 2329.340 214.160 ;
        RECT 2307.920 199.280 2308.180 199.540 ;
        RECT 2318.960 199.280 2319.220 199.540 ;
        RECT 2291.360 172.420 2291.620 172.680 ;
        RECT 2307.920 172.420 2308.180 172.680 ;
        RECT 2287.220 151.000 2287.480 151.260 ;
        RECT 2291.360 151.000 2291.620 151.260 ;
        RECT 2277.100 110.540 2277.360 110.800 ;
        RECT 2287.220 110.540 2287.480 110.800 ;
        RECT 2252.720 86.740 2252.980 87.000 ;
        RECT 2276.640 86.740 2276.900 87.000 ;
        RECT 1435.760 24.180 1436.020 24.440 ;
        RECT 2252.720 24.180 2252.980 24.440 ;
      LAYER met2 ;
        RECT 1729.240 3019.550 1729.500 3019.870 ;
        RECT 2463.400 3019.550 2463.660 3019.870 ;
        RECT 1729.300 3010.000 1729.440 3019.550 ;
        RECT 2463.460 3014.090 2463.600 3019.550 ;
        RECT 2463.400 3013.770 2463.660 3014.090 ;
        RECT 2491.000 3013.770 2491.260 3014.090 ;
        RECT 1729.300 3009.340 1729.650 3010.000 ;
        RECT 1729.370 3006.000 1729.650 3009.340 ;
        RECT 2491.060 3006.610 2491.200 3013.770 ;
        RECT 2491.000 3006.290 2491.260 3006.610 ;
        RECT 2519.980 3006.290 2520.240 3006.610 ;
        RECT 2520.040 2991.650 2520.180 3006.290 ;
        RECT 2519.980 2991.330 2520.240 2991.650 ;
        RECT 2615.660 2991.330 2615.920 2991.650 ;
        RECT 2615.720 473.610 2615.860 2991.330 ;
        RECT 2463.860 473.290 2464.120 473.610 ;
        RECT 2615.660 473.290 2615.920 473.610 ;
        RECT 2463.920 460.010 2464.060 473.290 ;
        RECT 2442.700 459.690 2442.960 460.010 ;
        RECT 2463.860 459.690 2464.120 460.010 ;
        RECT 2442.760 433.490 2442.900 459.690 ;
        RECT 2436.260 433.170 2436.520 433.490 ;
        RECT 2442.700 433.170 2442.960 433.490 ;
        RECT 2436.320 414.450 2436.460 433.170 ;
        RECT 2427.520 414.130 2427.780 414.450 ;
        RECT 2436.260 414.130 2436.520 414.450 ;
        RECT 2427.580 391.330 2427.720 414.130 ;
        RECT 2418.320 391.010 2418.580 391.330 ;
        RECT 2427.520 391.010 2427.780 391.330 ;
        RECT 2418.380 303.950 2418.520 391.010 ;
        RECT 2410.040 303.630 2410.300 303.950 ;
        RECT 2418.320 303.630 2418.580 303.950 ;
        RECT 2410.100 280.150 2410.240 303.630 ;
        RECT 2394.400 279.830 2394.660 280.150 ;
        RECT 2410.040 279.830 2410.300 280.150 ;
        RECT 2394.460 269.610 2394.600 279.830 ;
        RECT 2364.500 269.290 2364.760 269.610 ;
        RECT 2394.400 269.290 2394.660 269.610 ;
        RECT 2364.560 262.470 2364.700 269.290 ;
        RECT 2339.200 262.150 2339.460 262.470 ;
        RECT 2364.500 262.150 2364.760 262.470 ;
        RECT 2339.260 239.690 2339.400 262.150 ;
        RECT 2329.080 239.370 2329.340 239.690 ;
        RECT 2339.200 239.370 2339.460 239.690 ;
        RECT 2329.140 214.190 2329.280 239.370 ;
        RECT 2318.960 213.870 2319.220 214.190 ;
        RECT 2329.080 213.870 2329.340 214.190 ;
        RECT 2319.020 199.570 2319.160 213.870 ;
        RECT 2307.920 199.250 2308.180 199.570 ;
        RECT 2318.960 199.250 2319.220 199.570 ;
        RECT 2307.980 172.710 2308.120 199.250 ;
        RECT 2291.360 172.390 2291.620 172.710 ;
        RECT 2307.920 172.390 2308.180 172.710 ;
        RECT 2291.420 151.290 2291.560 172.390 ;
        RECT 2287.220 150.970 2287.480 151.290 ;
        RECT 2291.360 150.970 2291.620 151.290 ;
        RECT 2287.280 110.830 2287.420 150.970 ;
        RECT 2277.100 110.510 2277.360 110.830 ;
        RECT 2287.220 110.510 2287.480 110.830 ;
        RECT 2277.160 103.770 2277.300 110.510 ;
        RECT 2276.700 103.630 2277.300 103.770 ;
        RECT 2276.700 87.030 2276.840 103.630 ;
        RECT 2252.720 86.710 2252.980 87.030 ;
        RECT 2276.640 86.710 2276.900 87.030 ;
        RECT 2252.780 24.470 2252.920 86.710 ;
        RECT 1435.760 24.150 1436.020 24.470 ;
        RECT 2252.720 24.150 2252.980 24.470 ;
        RECT 1435.820 2.400 1435.960 24.150 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 302.290 2960.280 302.610 2960.340 ;
        RECT 393.370 2960.280 393.690 2960.340 ;
        RECT 302.290 2960.140 393.690 2960.280 ;
        RECT 302.290 2960.080 302.610 2960.140 ;
        RECT 393.370 2960.080 393.690 2960.140 ;
        RECT 302.290 46.480 302.610 46.540 ;
        RECT 1453.670 46.480 1453.990 46.540 ;
        RECT 302.290 46.340 1453.990 46.480 ;
        RECT 302.290 46.280 302.610 46.340 ;
        RECT 1453.670 46.280 1453.990 46.340 ;
      LAYER via ;
        RECT 302.320 2960.080 302.580 2960.340 ;
        RECT 393.400 2960.080 393.660 2960.340 ;
        RECT 302.320 46.280 302.580 46.540 ;
        RECT 1453.700 46.280 1453.960 46.540 ;
      LAYER met2 ;
        RECT 393.390 2960.875 393.670 2961.245 ;
        RECT 393.460 2960.370 393.600 2960.875 ;
        RECT 302.320 2960.050 302.580 2960.370 ;
        RECT 393.400 2960.050 393.660 2960.370 ;
        RECT 302.380 46.570 302.520 2960.050 ;
        RECT 302.320 46.250 302.580 46.570 ;
        RECT 1453.700 46.250 1453.960 46.570 ;
        RECT 1453.760 2.400 1453.900 46.250 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 393.390 2960.920 393.670 2961.200 ;
      LAYER met3 ;
        RECT 393.365 2961.210 393.695 2961.225 ;
        RECT 410.000 2961.210 414.000 2961.360 ;
        RECT 393.365 2960.910 414.000 2961.210 ;
        RECT 393.365 2960.895 393.695 2960.910 ;
        RECT 410.000 2960.760 414.000 2960.910 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1091.650 502.420 1091.970 502.480 ;
        RECT 1096.710 502.420 1097.030 502.480 ;
        RECT 1091.650 502.280 1097.030 502.420 ;
        RECT 1091.650 502.220 1091.970 502.280 ;
        RECT 1096.710 502.220 1097.030 502.280 ;
        RECT 1096.710 162.420 1097.030 162.480 ;
        RECT 1470.230 162.420 1470.550 162.480 ;
        RECT 1096.710 162.280 1470.550 162.420 ;
        RECT 1096.710 162.220 1097.030 162.280 ;
        RECT 1470.230 162.220 1470.550 162.280 ;
      LAYER via ;
        RECT 1091.680 502.220 1091.940 502.480 ;
        RECT 1096.740 502.220 1097.000 502.480 ;
        RECT 1096.740 162.220 1097.000 162.480 ;
        RECT 1470.260 162.220 1470.520 162.480 ;
      LAYER met2 ;
        RECT 1091.810 510.340 1092.090 514.000 ;
        RECT 1091.740 510.000 1092.090 510.340 ;
        RECT 1091.740 502.510 1091.880 510.000 ;
        RECT 1091.680 502.190 1091.940 502.510 ;
        RECT 1096.740 502.190 1097.000 502.510 ;
        RECT 1096.800 162.510 1096.940 502.190 ;
        RECT 1096.740 162.190 1097.000 162.510 ;
        RECT 1470.260 162.190 1470.520 162.510 ;
        RECT 1470.320 17.410 1470.460 162.190 ;
        RECT 1470.320 17.270 1471.840 17.410 ;
        RECT 1471.700 2.400 1471.840 17.270 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1489.090 148.820 1489.410 148.880 ;
        RECT 2152.870 148.820 2153.190 148.880 ;
        RECT 1489.090 148.680 2153.190 148.820 ;
        RECT 1489.090 148.620 1489.410 148.680 ;
        RECT 2152.870 148.620 2153.190 148.680 ;
      LAYER via ;
        RECT 1489.120 148.620 1489.380 148.880 ;
        RECT 2152.900 148.620 2153.160 148.880 ;
      LAYER met2 ;
        RECT 2154.410 510.410 2154.690 514.000 ;
        RECT 2152.960 510.270 2154.690 510.410 ;
        RECT 2152.960 148.910 2153.100 510.270 ;
        RECT 2154.410 510.000 2154.690 510.270 ;
        RECT 1489.120 148.590 1489.380 148.910 ;
        RECT 2152.900 148.590 2153.160 148.910 ;
        RECT 1489.180 17.410 1489.320 148.590 ;
        RECT 1489.180 17.270 1489.780 17.410 ;
        RECT 1489.640 2.400 1489.780 17.270 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1902.170 3043.580 1902.490 3043.640 ;
        RECT 2609.190 3043.580 2609.510 3043.640 ;
        RECT 1902.170 3043.440 2609.510 3043.580 ;
        RECT 1902.170 3043.380 1902.490 3043.440 ;
        RECT 2609.190 3043.380 2609.510 3043.440 ;
        RECT 1510.710 500.040 1511.030 500.100 ;
        RECT 2609.190 500.040 2609.510 500.100 ;
        RECT 1510.710 499.900 2609.510 500.040 ;
        RECT 1510.710 499.840 1511.030 499.900 ;
        RECT 2609.190 499.840 2609.510 499.900 ;
        RECT 1507.030 16.900 1507.350 16.960 ;
        RECT 1510.710 16.900 1511.030 16.960 ;
        RECT 1507.030 16.760 1511.030 16.900 ;
        RECT 1507.030 16.700 1507.350 16.760 ;
        RECT 1510.710 16.700 1511.030 16.760 ;
      LAYER via ;
        RECT 1902.200 3043.380 1902.460 3043.640 ;
        RECT 2609.220 3043.380 2609.480 3043.640 ;
        RECT 1510.740 499.840 1511.000 500.100 ;
        RECT 2609.220 499.840 2609.480 500.100 ;
        RECT 1507.060 16.700 1507.320 16.960 ;
        RECT 1510.740 16.700 1511.000 16.960 ;
      LAYER met2 ;
        RECT 1902.200 3043.350 1902.460 3043.670 ;
        RECT 2609.220 3043.350 2609.480 3043.670 ;
        RECT 1902.260 3010.000 1902.400 3043.350 ;
        RECT 1902.260 3009.340 1902.610 3010.000 ;
        RECT 1902.330 3006.000 1902.610 3009.340 ;
        RECT 2609.280 500.130 2609.420 3043.350 ;
        RECT 1510.740 499.810 1511.000 500.130 ;
        RECT 2609.220 499.810 2609.480 500.130 ;
        RECT 1510.800 16.990 1510.940 499.810 ;
        RECT 1507.060 16.670 1507.320 16.990 ;
        RECT 1510.740 16.670 1511.000 16.990 ;
        RECT 1507.120 2.400 1507.260 16.670 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 703.485 234.685 703.655 282.795 ;
        RECT 703.945 179.605 704.115 227.715 ;
        RECT 703.945 48.365 704.115 113.475 ;
      LAYER mcon ;
        RECT 703.485 282.625 703.655 282.795 ;
        RECT 703.945 227.545 704.115 227.715 ;
        RECT 703.945 113.305 704.115 113.475 ;
      LAYER met1 ;
        RECT 412.690 502.760 413.010 502.820 ;
        RECT 424.650 502.760 424.970 502.820 ;
        RECT 412.690 502.620 424.970 502.760 ;
        RECT 412.690 502.560 413.010 502.620 ;
        RECT 424.650 502.560 424.970 502.620 ;
        RECT 424.650 438.160 424.970 438.220 ;
        RECT 690.070 438.160 690.390 438.220 ;
        RECT 424.650 438.020 690.390 438.160 ;
        RECT 424.650 437.960 424.970 438.020 ;
        RECT 690.070 437.960 690.390 438.020 ;
        RECT 703.870 337.860 704.190 337.920 ;
        RECT 704.330 337.860 704.650 337.920 ;
        RECT 703.870 337.720 704.650 337.860 ;
        RECT 703.870 337.660 704.190 337.720 ;
        RECT 704.330 337.660 704.650 337.720 ;
        RECT 703.410 289.580 703.730 289.640 ;
        RECT 703.870 289.580 704.190 289.640 ;
        RECT 703.410 289.440 704.190 289.580 ;
        RECT 703.410 289.380 703.730 289.440 ;
        RECT 703.870 289.380 704.190 289.440 ;
        RECT 703.410 282.780 703.730 282.840 ;
        RECT 703.215 282.640 703.730 282.780 ;
        RECT 703.410 282.580 703.730 282.640 ;
        RECT 703.425 234.840 703.715 234.885 ;
        RECT 703.870 234.840 704.190 234.900 ;
        RECT 703.425 234.700 704.190 234.840 ;
        RECT 703.425 234.655 703.715 234.700 ;
        RECT 703.870 234.640 704.190 234.700 ;
        RECT 703.870 227.700 704.190 227.760 ;
        RECT 703.675 227.560 704.190 227.700 ;
        RECT 703.870 227.500 704.190 227.560 ;
        RECT 703.885 179.760 704.175 179.805 ;
        RECT 704.330 179.760 704.650 179.820 ;
        RECT 703.885 179.620 704.650 179.760 ;
        RECT 703.885 179.575 704.175 179.620 ;
        RECT 704.330 179.560 704.650 179.620 ;
        RECT 703.885 113.460 704.175 113.505 ;
        RECT 704.330 113.460 704.650 113.520 ;
        RECT 703.885 113.320 704.650 113.460 ;
        RECT 703.885 113.275 704.175 113.320 ;
        RECT 704.330 113.260 704.650 113.320 ;
        RECT 703.870 48.520 704.190 48.580 ;
        RECT 703.675 48.380 704.190 48.520 ;
        RECT 703.870 48.320 704.190 48.380 ;
      LAYER via ;
        RECT 412.720 502.560 412.980 502.820 ;
        RECT 424.680 502.560 424.940 502.820 ;
        RECT 424.680 437.960 424.940 438.220 ;
        RECT 690.100 437.960 690.360 438.220 ;
        RECT 703.900 337.660 704.160 337.920 ;
        RECT 704.360 337.660 704.620 337.920 ;
        RECT 703.440 289.380 703.700 289.640 ;
        RECT 703.900 289.380 704.160 289.640 ;
        RECT 703.440 282.580 703.700 282.840 ;
        RECT 703.900 234.640 704.160 234.900 ;
        RECT 703.900 227.500 704.160 227.760 ;
        RECT 704.360 179.560 704.620 179.820 ;
        RECT 704.360 113.260 704.620 113.520 ;
        RECT 703.900 48.320 704.160 48.580 ;
      LAYER met2 ;
        RECT 412.850 510.340 413.130 514.000 ;
        RECT 412.780 510.000 413.130 510.340 ;
        RECT 412.780 502.850 412.920 510.000 ;
        RECT 412.720 502.530 412.980 502.850 ;
        RECT 424.680 502.530 424.940 502.850 ;
        RECT 424.740 438.250 424.880 502.530 ;
        RECT 424.680 437.930 424.940 438.250 ;
        RECT 690.100 437.930 690.360 438.250 ;
        RECT 690.160 435.045 690.300 437.930 ;
        RECT 690.090 434.675 690.370 435.045 ;
        RECT 703.890 434.675 704.170 435.045 ;
        RECT 703.960 386.085 704.100 434.675 ;
        RECT 702.510 385.715 702.790 386.085 ;
        RECT 703.890 385.715 704.170 386.085 ;
        RECT 702.580 338.485 702.720 385.715 ;
        RECT 702.510 338.115 702.790 338.485 ;
        RECT 703.890 338.115 704.170 338.485 ;
        RECT 703.960 337.950 704.100 338.115 ;
        RECT 703.900 337.630 704.160 337.950 ;
        RECT 704.360 337.630 704.620 337.950 ;
        RECT 704.420 290.090 704.560 337.630 ;
        RECT 703.960 289.950 704.560 290.090 ;
        RECT 703.960 289.670 704.100 289.950 ;
        RECT 703.440 289.350 703.700 289.670 ;
        RECT 703.900 289.350 704.160 289.670 ;
        RECT 703.500 282.870 703.640 289.350 ;
        RECT 703.440 282.550 703.700 282.870 ;
        RECT 703.900 234.610 704.160 234.930 ;
        RECT 703.960 227.790 704.100 234.610 ;
        RECT 703.900 227.470 704.160 227.790 ;
        RECT 704.360 179.530 704.620 179.850 ;
        RECT 704.420 146.610 704.560 179.530 ;
        RECT 704.420 146.470 705.020 146.610 ;
        RECT 704.880 144.570 705.020 146.470 ;
        RECT 703.960 144.430 705.020 144.570 ;
        RECT 703.960 137.770 704.100 144.430 ;
        RECT 703.960 137.630 704.560 137.770 ;
        RECT 704.420 113.550 704.560 137.630 ;
        RECT 704.360 113.230 704.620 113.550 ;
        RECT 703.900 48.290 704.160 48.610 ;
        RECT 703.960 24.210 704.100 48.290 ;
        RECT 703.960 24.070 704.560 24.210 ;
        RECT 704.420 2.400 704.560 24.070 ;
        RECT 704.210 -4.800 704.770 2.400 ;
      LAYER via2 ;
        RECT 690.090 434.720 690.370 435.000 ;
        RECT 703.890 434.720 704.170 435.000 ;
        RECT 702.510 385.760 702.790 386.040 ;
        RECT 703.890 385.760 704.170 386.040 ;
        RECT 702.510 338.160 702.790 338.440 ;
        RECT 703.890 338.160 704.170 338.440 ;
      LAYER met3 ;
        RECT 690.065 435.010 690.395 435.025 ;
        RECT 703.865 435.010 704.195 435.025 ;
        RECT 690.065 434.710 704.195 435.010 ;
        RECT 690.065 434.695 690.395 434.710 ;
        RECT 703.865 434.695 704.195 434.710 ;
        RECT 702.485 386.050 702.815 386.065 ;
        RECT 703.865 386.050 704.195 386.065 ;
        RECT 702.485 385.750 704.195 386.050 ;
        RECT 702.485 385.735 702.815 385.750 ;
        RECT 703.865 385.735 704.195 385.750 ;
        RECT 702.485 338.450 702.815 338.465 ;
        RECT 703.865 338.450 704.195 338.465 ;
        RECT 702.485 338.150 704.195 338.450 ;
        RECT 702.485 338.135 702.815 338.150 ;
        RECT 703.865 338.135 704.195 338.150 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2346.240 2519.810 2346.300 ;
        RECT 2553.990 2346.240 2554.310 2346.300 ;
        RECT 2519.490 2346.100 2554.310 2346.240 ;
        RECT 2519.490 2346.040 2519.810 2346.100 ;
        RECT 2553.990 2346.040 2554.310 2346.100 ;
        RECT 1531.410 494.940 1531.730 495.000 ;
        RECT 2553.990 494.940 2554.310 495.000 ;
        RECT 1531.410 494.800 2554.310 494.940 ;
        RECT 1531.410 494.740 1531.730 494.800 ;
        RECT 2553.990 494.740 2554.310 494.800 ;
        RECT 1524.970 16.220 1525.290 16.280 ;
        RECT 1531.410 16.220 1531.730 16.280 ;
        RECT 1524.970 16.080 1531.730 16.220 ;
        RECT 1524.970 16.020 1525.290 16.080 ;
        RECT 1531.410 16.020 1531.730 16.080 ;
      LAYER via ;
        RECT 2519.520 2346.040 2519.780 2346.300 ;
        RECT 2554.020 2346.040 2554.280 2346.300 ;
        RECT 1531.440 494.740 1531.700 495.000 ;
        RECT 2554.020 494.740 2554.280 495.000 ;
        RECT 1525.000 16.020 1525.260 16.280 ;
        RECT 1531.440 16.020 1531.700 16.280 ;
      LAYER met2 ;
        RECT 2519.510 2347.515 2519.790 2347.885 ;
        RECT 2519.580 2346.330 2519.720 2347.515 ;
        RECT 2519.520 2346.010 2519.780 2346.330 ;
        RECT 2554.020 2346.010 2554.280 2346.330 ;
        RECT 2554.080 495.030 2554.220 2346.010 ;
        RECT 1531.440 494.710 1531.700 495.030 ;
        RECT 2554.020 494.710 2554.280 495.030 ;
        RECT 1531.500 16.310 1531.640 494.710 ;
        RECT 1525.000 15.990 1525.260 16.310 ;
        RECT 1531.440 15.990 1531.700 16.310 ;
        RECT 1525.060 2.400 1525.200 15.990 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2347.560 2519.790 2347.840 ;
      LAYER met3 ;
        RECT 2506.000 2347.850 2510.000 2348.000 ;
        RECT 2519.485 2347.850 2519.815 2347.865 ;
        RECT 2506.000 2347.550 2519.815 2347.850 ;
        RECT 2506.000 2347.400 2510.000 2347.550 ;
        RECT 2519.485 2347.535 2519.815 2347.550 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 342.770 1462.920 343.090 1462.980 ;
        RECT 393.370 1462.920 393.690 1462.980 ;
        RECT 342.770 1462.780 393.690 1462.920 ;
        RECT 342.770 1462.720 343.090 1462.780 ;
        RECT 393.370 1462.720 393.690 1462.780 ;
        RECT 342.770 45.800 343.090 45.860 ;
        RECT 1542.910 45.800 1543.230 45.860 ;
        RECT 342.770 45.660 1543.230 45.800 ;
        RECT 342.770 45.600 343.090 45.660 ;
        RECT 1542.910 45.600 1543.230 45.660 ;
      LAYER via ;
        RECT 342.800 1462.720 343.060 1462.980 ;
        RECT 393.400 1462.720 393.660 1462.980 ;
        RECT 342.800 45.600 343.060 45.860 ;
        RECT 1542.940 45.600 1543.200 45.860 ;
      LAYER met2 ;
        RECT 393.390 1463.515 393.670 1463.885 ;
        RECT 393.460 1463.010 393.600 1463.515 ;
        RECT 342.800 1462.690 343.060 1463.010 ;
        RECT 393.400 1462.690 393.660 1463.010 ;
        RECT 342.860 45.890 343.000 1462.690 ;
        RECT 342.800 45.570 343.060 45.890 ;
        RECT 1542.940 45.570 1543.200 45.890 ;
        RECT 1543.000 2.400 1543.140 45.570 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 393.390 1463.560 393.670 1463.840 ;
      LAYER met3 ;
        RECT 393.365 1463.850 393.695 1463.865 ;
        RECT 410.000 1463.850 414.000 1464.000 ;
        RECT 393.365 1463.550 414.000 1463.850 ;
        RECT 393.365 1463.535 393.695 1463.550 ;
        RECT 410.000 1463.400 414.000 1463.550 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 307.600 537.670 307.660 ;
        RECT 1559.930 307.600 1560.250 307.660 ;
        RECT 537.350 307.460 1560.250 307.600 ;
        RECT 537.350 307.400 537.670 307.460 ;
        RECT 1559.930 307.400 1560.250 307.460 ;
      LAYER via ;
        RECT 537.380 307.400 537.640 307.660 ;
        RECT 1559.960 307.400 1560.220 307.660 ;
      LAYER met2 ;
        RECT 536.130 510.410 536.410 514.000 ;
        RECT 536.130 510.270 537.580 510.410 ;
        RECT 536.130 510.000 536.410 510.270 ;
        RECT 537.440 307.690 537.580 510.270 ;
        RECT 537.380 307.370 537.640 307.690 ;
        RECT 1559.960 307.370 1560.220 307.690 ;
        RECT 1560.020 17.410 1560.160 307.370 ;
        RECT 1560.020 17.270 1561.080 17.410 ;
        RECT 1560.940 2.400 1561.080 17.270 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 328.000 1580.030 328.060 ;
        RECT 2526.390 328.000 2526.710 328.060 ;
        RECT 1579.710 327.860 2526.710 328.000 ;
        RECT 1579.710 327.800 1580.030 327.860 ;
        RECT 2526.390 327.800 2526.710 327.860 ;
      LAYER via ;
        RECT 1579.740 327.800 1580.000 328.060 ;
        RECT 2526.420 327.800 2526.680 328.060 ;
      LAYER met2 ;
        RECT 2526.410 1781.755 2526.690 1782.125 ;
        RECT 2526.480 328.090 2526.620 1781.755 ;
        RECT 1579.740 327.770 1580.000 328.090 ;
        RECT 2526.420 327.770 2526.680 328.090 ;
        RECT 1579.800 17.410 1579.940 327.770 ;
        RECT 1578.880 17.270 1579.940 17.410 ;
        RECT 1578.880 2.400 1579.020 17.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
      LAYER via2 ;
        RECT 2526.410 1781.800 2526.690 1782.080 ;
      LAYER met3 ;
        RECT 2506.000 1782.090 2510.000 1782.240 ;
        RECT 2526.385 1782.090 2526.715 1782.105 ;
        RECT 2506.000 1781.790 2526.715 1782.090 ;
        RECT 2506.000 1781.640 2510.000 1781.790 ;
        RECT 2526.385 1781.775 2526.715 1781.790 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1596.270 15.200 1596.590 15.260 ;
        RECT 1599.950 15.200 1600.270 15.260 ;
        RECT 1596.270 15.060 1600.270 15.200 ;
        RECT 1596.270 15.000 1596.590 15.060 ;
        RECT 1599.950 15.000 1600.270 15.060 ;
      LAYER via ;
        RECT 1596.300 15.000 1596.560 15.260 ;
        RECT 1599.980 15.000 1600.240 15.260 ;
      LAYER met2 ;
        RECT 1963.830 3024.795 1964.110 3025.165 ;
        RECT 1963.900 3010.000 1964.040 3024.795 ;
        RECT 1963.900 3009.340 1964.250 3010.000 ;
        RECT 1963.970 3006.000 1964.250 3009.340 ;
        RECT 1599.970 479.555 1600.250 479.925 ;
        RECT 1600.040 15.290 1600.180 479.555 ;
        RECT 1596.300 14.970 1596.560 15.290 ;
        RECT 1599.980 14.970 1600.240 15.290 ;
        RECT 1596.360 2.400 1596.500 14.970 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
      LAYER via2 ;
        RECT 1963.830 3024.840 1964.110 3025.120 ;
        RECT 1599.970 479.600 1600.250 479.880 ;
      LAYER met3 ;
        RECT 1963.805 3025.130 1964.135 3025.145 ;
        RECT 2464.030 3025.130 2464.410 3025.140 ;
        RECT 1963.805 3024.830 2464.410 3025.130 ;
        RECT 1963.805 3024.815 1964.135 3024.830 ;
        RECT 2464.030 3024.820 2464.410 3024.830 ;
        RECT 2464.030 512.220 2464.410 512.540 ;
        RECT 2464.070 511.180 2464.370 512.220 ;
        RECT 2464.030 510.860 2464.410 511.180 ;
        RECT 1599.945 479.890 1600.275 479.905 ;
        RECT 2464.030 479.890 2464.410 479.900 ;
        RECT 1599.945 479.590 2464.410 479.890 ;
        RECT 1599.945 479.575 1600.275 479.590 ;
        RECT 2464.030 479.580 2464.410 479.590 ;
      LAYER via3 ;
        RECT 2464.060 3024.820 2464.380 3025.140 ;
        RECT 2464.060 512.220 2464.380 512.540 ;
        RECT 2464.060 510.860 2464.380 511.180 ;
        RECT 2464.060 479.580 2464.380 479.900 ;
      LAYER met4 ;
        RECT 2464.055 3024.815 2464.385 3025.145 ;
        RECT 2464.070 512.545 2464.370 3024.815 ;
        RECT 2464.055 512.215 2464.385 512.545 ;
        RECT 2464.055 510.855 2464.385 511.185 ;
        RECT 2464.070 479.905 2464.370 510.855 ;
        RECT 2464.055 479.575 2464.385 479.905 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2421.050 3017.400 2421.370 3017.460 ;
        RECT 2588.030 3017.400 2588.350 3017.460 ;
        RECT 2421.050 3017.260 2588.350 3017.400 ;
        RECT 2421.050 3017.200 2421.370 3017.260 ;
        RECT 2588.030 3017.200 2588.350 3017.260 ;
        RECT 1614.670 17.920 1614.990 17.980 ;
        RECT 2588.030 17.920 2588.350 17.980 ;
        RECT 1614.670 17.780 2588.350 17.920 ;
        RECT 1614.670 17.720 1614.990 17.780 ;
        RECT 2588.030 17.720 2588.350 17.780 ;
      LAYER via ;
        RECT 2421.080 3017.200 2421.340 3017.460 ;
        RECT 2588.060 3017.200 2588.320 3017.460 ;
        RECT 1614.700 17.720 1614.960 17.980 ;
        RECT 2588.060 17.720 2588.320 17.980 ;
      LAYER met2 ;
        RECT 2421.080 3017.170 2421.340 3017.490 ;
        RECT 2588.060 3017.170 2588.320 3017.490 ;
        RECT 2421.140 3010.000 2421.280 3017.170 ;
        RECT 2421.140 3009.340 2421.490 3010.000 ;
        RECT 2421.210 3006.000 2421.490 3009.340 ;
        RECT 2588.120 18.010 2588.260 3017.170 ;
        RECT 1614.700 17.690 1614.960 18.010 ;
        RECT 2588.060 17.690 2588.320 18.010 ;
        RECT 1614.760 17.410 1614.900 17.690 ;
        RECT 1614.300 17.270 1614.900 17.410 ;
        RECT 1614.300 2.400 1614.440 17.270 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2726.020 2519.810 2726.080 ;
        RECT 2575.150 2726.020 2575.470 2726.080 ;
        RECT 2519.490 2725.880 2575.470 2726.020 ;
        RECT 2519.490 2725.820 2519.810 2725.880 ;
        RECT 2575.150 2725.820 2575.470 2725.880 ;
        RECT 1634.910 480.660 1635.230 480.720 ;
        RECT 2575.150 480.660 2575.470 480.720 ;
        RECT 1634.910 480.520 2575.470 480.660 ;
        RECT 1634.910 480.460 1635.230 480.520 ;
        RECT 2575.150 480.460 2575.470 480.520 ;
        RECT 1632.150 16.900 1632.470 16.960 ;
        RECT 1634.910 16.900 1635.230 16.960 ;
        RECT 1632.150 16.760 1635.230 16.900 ;
        RECT 1632.150 16.700 1632.470 16.760 ;
        RECT 1634.910 16.700 1635.230 16.760 ;
      LAYER via ;
        RECT 2519.520 2725.820 2519.780 2726.080 ;
        RECT 2575.180 2725.820 2575.440 2726.080 ;
        RECT 1634.940 480.460 1635.200 480.720 ;
        RECT 2575.180 480.460 2575.440 480.720 ;
        RECT 1632.180 16.700 1632.440 16.960 ;
        RECT 1634.940 16.700 1635.200 16.960 ;
      LAYER met2 ;
        RECT 2519.510 2731.035 2519.790 2731.405 ;
        RECT 2519.580 2726.110 2519.720 2731.035 ;
        RECT 2519.520 2725.790 2519.780 2726.110 ;
        RECT 2575.180 2725.790 2575.440 2726.110 ;
        RECT 2575.240 480.750 2575.380 2725.790 ;
        RECT 1634.940 480.430 1635.200 480.750 ;
        RECT 2575.180 480.430 2575.440 480.750 ;
        RECT 1635.000 16.990 1635.140 480.430 ;
        RECT 1632.180 16.670 1632.440 16.990 ;
        RECT 1634.940 16.670 1635.200 16.990 ;
        RECT 1632.240 2.400 1632.380 16.670 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2731.080 2519.790 2731.360 ;
      LAYER met3 ;
        RECT 2506.000 2731.370 2510.000 2731.520 ;
        RECT 2519.485 2731.370 2519.815 2731.385 ;
        RECT 2506.000 2731.070 2519.815 2731.370 ;
        RECT 2506.000 2730.920 2510.000 2731.070 ;
        RECT 2519.485 2731.055 2519.815 2731.070 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2801.500 2519.810 2801.560 ;
        RECT 2603.210 2801.500 2603.530 2801.560 ;
        RECT 2519.490 2801.360 2603.530 2801.500 ;
        RECT 2519.490 2801.300 2519.810 2801.360 ;
        RECT 2603.210 2801.300 2603.530 2801.360 ;
        RECT 1655.610 495.280 1655.930 495.340 ;
        RECT 2603.210 495.280 2603.530 495.340 ;
        RECT 1655.610 495.140 2603.530 495.280 ;
        RECT 1655.610 495.080 1655.930 495.140 ;
        RECT 2603.210 495.080 2603.530 495.140 ;
        RECT 1650.090 16.900 1650.410 16.960 ;
        RECT 1655.610 16.900 1655.930 16.960 ;
        RECT 1650.090 16.760 1655.930 16.900 ;
        RECT 1650.090 16.700 1650.410 16.760 ;
        RECT 1655.610 16.700 1655.930 16.760 ;
      LAYER via ;
        RECT 2519.520 2801.300 2519.780 2801.560 ;
        RECT 2603.240 2801.300 2603.500 2801.560 ;
        RECT 1655.640 495.080 1655.900 495.340 ;
        RECT 2603.240 495.080 2603.500 495.340 ;
        RECT 1650.120 16.700 1650.380 16.960 ;
        RECT 1655.640 16.700 1655.900 16.960 ;
      LAYER met2 ;
        RECT 2519.510 2804.475 2519.790 2804.845 ;
        RECT 2519.580 2801.590 2519.720 2804.475 ;
        RECT 2519.520 2801.270 2519.780 2801.590 ;
        RECT 2603.240 2801.270 2603.500 2801.590 ;
        RECT 2603.300 495.370 2603.440 2801.270 ;
        RECT 1655.640 495.050 1655.900 495.370 ;
        RECT 2603.240 495.050 2603.500 495.370 ;
        RECT 1655.700 16.990 1655.840 495.050 ;
        RECT 1650.120 16.670 1650.380 16.990 ;
        RECT 1655.640 16.670 1655.900 16.990 ;
        RECT 1650.180 2.400 1650.320 16.670 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2804.520 2519.790 2804.800 ;
      LAYER met3 ;
        RECT 2506.000 2804.810 2510.000 2804.960 ;
        RECT 2519.485 2804.810 2519.815 2804.825 ;
        RECT 2506.000 2804.510 2519.815 2804.810 ;
        RECT 2506.000 2804.360 2510.000 2804.510 ;
        RECT 2519.485 2804.495 2519.815 2804.510 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1669.485 241.485 1669.655 289.595 ;
        RECT 1669.485 48.365 1669.655 96.475 ;
      LAYER mcon ;
        RECT 1669.485 289.425 1669.655 289.595 ;
        RECT 1669.485 96.305 1669.655 96.475 ;
      LAYER met1 ;
        RECT 1669.410 300.800 1669.730 300.860 ;
        RECT 2283.970 300.800 2284.290 300.860 ;
        RECT 1669.410 300.660 2284.290 300.800 ;
        RECT 1669.410 300.600 1669.730 300.660 ;
        RECT 2283.970 300.600 2284.290 300.660 ;
        RECT 1669.410 289.580 1669.730 289.640 ;
        RECT 1669.215 289.440 1669.730 289.580 ;
        RECT 1669.410 289.380 1669.730 289.440 ;
        RECT 1669.410 241.640 1669.730 241.700 ;
        RECT 1669.215 241.500 1669.730 241.640 ;
        RECT 1669.410 241.440 1669.730 241.500 ;
        RECT 1669.410 96.460 1669.730 96.520 ;
        RECT 1669.215 96.320 1669.730 96.460 ;
        RECT 1669.410 96.260 1669.730 96.320 ;
        RECT 1669.410 48.520 1669.730 48.580 ;
        RECT 1669.215 48.380 1669.730 48.520 ;
        RECT 1669.410 48.320 1669.730 48.380 ;
        RECT 1669.410 14.180 1669.730 14.240 ;
        RECT 1668.120 14.040 1669.730 14.180 ;
        RECT 1668.120 13.900 1668.260 14.040 ;
        RECT 1669.410 13.980 1669.730 14.040 ;
        RECT 1668.030 13.640 1668.350 13.900 ;
      LAYER via ;
        RECT 1669.440 300.600 1669.700 300.860 ;
        RECT 2284.000 300.600 2284.260 300.860 ;
        RECT 1669.440 289.380 1669.700 289.640 ;
        RECT 1669.440 241.440 1669.700 241.700 ;
        RECT 1669.440 96.260 1669.700 96.520 ;
        RECT 1669.440 48.320 1669.700 48.580 ;
        RECT 1669.440 13.980 1669.700 14.240 ;
        RECT 1668.060 13.640 1668.320 13.900 ;
      LAYER met2 ;
        RECT 2290.570 510.410 2290.850 514.000 ;
        RECT 2284.060 510.270 2290.850 510.410 ;
        RECT 2284.060 300.890 2284.200 510.270 ;
        RECT 2290.570 510.000 2290.850 510.270 ;
        RECT 1669.440 300.570 1669.700 300.890 ;
        RECT 2284.000 300.570 2284.260 300.890 ;
        RECT 1669.500 289.670 1669.640 300.570 ;
        RECT 1669.440 289.350 1669.700 289.670 ;
        RECT 1669.440 241.410 1669.700 241.730 ;
        RECT 1669.500 96.550 1669.640 241.410 ;
        RECT 1669.440 96.230 1669.700 96.550 ;
        RECT 1669.440 48.290 1669.700 48.610 ;
        RECT 1669.500 14.270 1669.640 48.290 ;
        RECT 1669.440 13.950 1669.700 14.270 ;
        RECT 1668.060 13.610 1668.320 13.930 ;
        RECT 1668.120 2.400 1668.260 13.610 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.110 348.740 1690.430 348.800 ;
        RECT 2484.070 348.740 2484.390 348.800 ;
        RECT 1690.110 348.600 2484.390 348.740 ;
        RECT 1690.110 348.540 1690.430 348.600 ;
        RECT 2484.070 348.540 2484.390 348.600 ;
        RECT 1685.510 20.300 1685.830 20.360 ;
        RECT 1690.110 20.300 1690.430 20.360 ;
        RECT 1685.510 20.160 1690.430 20.300 ;
        RECT 1685.510 20.100 1685.830 20.160 ;
        RECT 1690.110 20.100 1690.430 20.160 ;
      LAYER via ;
        RECT 1690.140 348.540 1690.400 348.800 ;
        RECT 2484.100 348.540 2484.360 348.800 ;
        RECT 1685.540 20.100 1685.800 20.360 ;
        RECT 1690.140 20.100 1690.400 20.360 ;
      LAYER met2 ;
        RECT 2487.450 510.410 2487.730 514.000 ;
        RECT 2484.160 510.270 2487.730 510.410 ;
        RECT 2484.160 348.830 2484.300 510.270 ;
        RECT 2487.450 510.000 2487.730 510.270 ;
        RECT 1690.140 348.510 1690.400 348.830 ;
        RECT 2484.100 348.510 2484.360 348.830 ;
        RECT 1690.200 20.390 1690.340 348.510 ;
        RECT 1685.540 20.070 1685.800 20.390 ;
        RECT 1690.140 20.070 1690.400 20.390 ;
        RECT 1685.600 2.400 1685.740 20.070 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 723.725 241.485 723.895 289.595 ;
        RECT 723.725 144.925 723.895 193.035 ;
        RECT 723.725 48.365 723.895 96.475 ;
      LAYER mcon ;
        RECT 723.725 289.425 723.895 289.595 ;
        RECT 723.725 192.865 723.895 193.035 ;
        RECT 723.725 96.305 723.895 96.475 ;
      LAYER met1 ;
        RECT 723.190 294.000 723.510 294.060 ;
        RECT 1980.830 294.000 1981.150 294.060 ;
        RECT 723.190 293.860 1981.150 294.000 ;
        RECT 723.190 293.800 723.510 293.860 ;
        RECT 1980.830 293.800 1981.150 293.860 ;
        RECT 723.650 289.580 723.970 289.640 ;
        RECT 723.455 289.440 723.970 289.580 ;
        RECT 723.650 289.380 723.970 289.440 ;
        RECT 723.650 241.640 723.970 241.700 ;
        RECT 723.455 241.500 723.970 241.640 ;
        RECT 723.650 241.440 723.970 241.500 ;
        RECT 723.650 193.020 723.970 193.080 ;
        RECT 723.455 192.880 723.970 193.020 ;
        RECT 723.650 192.820 723.970 192.880 ;
        RECT 723.650 145.080 723.970 145.140 ;
        RECT 723.455 144.940 723.970 145.080 ;
        RECT 723.650 144.880 723.970 144.940 ;
        RECT 723.650 96.460 723.970 96.520 ;
        RECT 723.455 96.320 723.970 96.460 ;
        RECT 723.650 96.260 723.970 96.320 ;
        RECT 723.650 48.520 723.970 48.580 ;
        RECT 723.455 48.380 723.970 48.520 ;
        RECT 723.650 48.320 723.970 48.380 ;
        RECT 723.650 14.180 723.970 14.240 ;
        RECT 722.360 14.040 723.970 14.180 ;
        RECT 722.360 13.900 722.500 14.040 ;
        RECT 723.650 13.980 723.970 14.040 ;
        RECT 722.270 13.640 722.590 13.900 ;
      LAYER via ;
        RECT 723.220 293.800 723.480 294.060 ;
        RECT 1980.860 293.800 1981.120 294.060 ;
        RECT 723.680 289.380 723.940 289.640 ;
        RECT 723.680 241.440 723.940 241.700 ;
        RECT 723.680 192.820 723.940 193.080 ;
        RECT 723.680 144.880 723.940 145.140 ;
        RECT 723.680 96.260 723.940 96.520 ;
        RECT 723.680 48.320 723.940 48.580 ;
        RECT 723.680 13.980 723.940 14.240 ;
        RECT 722.300 13.640 722.560 13.900 ;
      LAYER met2 ;
        RECT 1981.450 510.410 1981.730 514.000 ;
        RECT 1980.920 510.270 1981.730 510.410 ;
        RECT 1980.920 294.090 1981.060 510.270 ;
        RECT 1981.450 510.000 1981.730 510.270 ;
        RECT 723.220 293.770 723.480 294.090 ;
        RECT 1980.860 293.770 1981.120 294.090 ;
        RECT 723.280 290.090 723.420 293.770 ;
        RECT 723.280 289.950 723.880 290.090 ;
        RECT 723.740 289.670 723.880 289.950 ;
        RECT 723.680 289.350 723.940 289.670 ;
        RECT 723.680 241.410 723.940 241.730 ;
        RECT 723.740 193.110 723.880 241.410 ;
        RECT 723.680 192.790 723.940 193.110 ;
        RECT 723.680 144.850 723.940 145.170 ;
        RECT 723.740 96.550 723.880 144.850 ;
        RECT 723.680 96.230 723.940 96.550 ;
        RECT 723.680 48.290 723.940 48.610 ;
        RECT 723.740 14.270 723.880 48.290 ;
        RECT 723.680 13.950 723.940 14.270 ;
        RECT 722.300 13.610 722.560 13.930 ;
        RECT 722.360 2.400 722.500 13.610 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 350.130 1366.360 350.450 1366.420 ;
        RECT 393.370 1366.360 393.690 1366.420 ;
        RECT 350.130 1366.220 393.690 1366.360 ;
        RECT 350.130 1366.160 350.450 1366.220 ;
        RECT 393.370 1366.160 393.690 1366.220 ;
        RECT 350.130 45.120 350.450 45.180 ;
        RECT 1703.450 45.120 1703.770 45.180 ;
        RECT 350.130 44.980 1703.770 45.120 ;
        RECT 350.130 44.920 350.450 44.980 ;
        RECT 1703.450 44.920 1703.770 44.980 ;
      LAYER via ;
        RECT 350.160 1366.160 350.420 1366.420 ;
        RECT 393.400 1366.160 393.660 1366.420 ;
        RECT 350.160 44.920 350.420 45.180 ;
        RECT 1703.480 44.920 1703.740 45.180 ;
      LAYER met2 ;
        RECT 393.390 1372.395 393.670 1372.765 ;
        RECT 393.460 1366.450 393.600 1372.395 ;
        RECT 350.160 1366.130 350.420 1366.450 ;
        RECT 393.400 1366.130 393.660 1366.450 ;
        RECT 350.220 45.210 350.360 1366.130 ;
        RECT 350.160 44.890 350.420 45.210 ;
        RECT 1703.480 44.890 1703.740 45.210 ;
        RECT 1703.540 2.400 1703.680 44.890 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
      LAYER via2 ;
        RECT 393.390 1372.440 393.670 1372.720 ;
      LAYER met3 ;
        RECT 393.365 1372.730 393.695 1372.745 ;
        RECT 410.000 1372.730 414.000 1372.880 ;
        RECT 393.365 1372.430 414.000 1372.730 ;
        RECT 393.365 1372.415 393.695 1372.430 ;
        RECT 410.000 1372.280 414.000 1372.430 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1721.390 16.900 1721.710 16.960 ;
        RECT 1724.610 16.900 1724.930 16.960 ;
        RECT 1721.390 16.760 1724.930 16.900 ;
        RECT 1721.390 16.700 1721.710 16.760 ;
        RECT 1724.610 16.700 1724.930 16.760 ;
      LAYER via ;
        RECT 1721.420 16.700 1721.680 16.960 ;
        RECT 1724.640 16.700 1724.900 16.960 ;
      LAYER met2 ;
        RECT 2609.670 2897.635 2609.950 2898.005 ;
        RECT 2609.740 2851.085 2609.880 2897.635 ;
        RECT 2609.670 2850.715 2609.950 2851.085 ;
        RECT 2610.590 2801.075 2610.870 2801.445 ;
        RECT 2610.660 2753.845 2610.800 2801.075 ;
        RECT 2610.590 2753.475 2610.870 2753.845 ;
        RECT 2610.130 2704.515 2610.410 2704.885 ;
        RECT 2610.200 2657.965 2610.340 2704.515 ;
        RECT 2610.130 2657.595 2610.410 2657.965 ;
        RECT 2610.130 2607.955 2610.410 2608.325 ;
        RECT 2610.200 2561.405 2610.340 2607.955 ;
        RECT 2610.130 2561.035 2610.410 2561.405 ;
        RECT 2610.130 2511.395 2610.410 2511.765 ;
        RECT 2610.200 2463.485 2610.340 2511.395 ;
        RECT 2610.130 2463.115 2610.410 2463.485 ;
        RECT 2610.590 2316.915 2610.870 2317.285 ;
        RECT 2610.660 2270.365 2610.800 2316.915 ;
        RECT 2610.590 2269.995 2610.870 2270.365 ;
        RECT 2611.050 2124.475 2611.330 2124.845 ;
        RECT 2611.120 2077.245 2611.260 2124.475 ;
        RECT 2611.050 2076.875 2611.330 2077.245 ;
        RECT 2611.050 2027.235 2611.330 2027.605 ;
        RECT 2611.120 1980.685 2611.260 2027.235 ;
        RECT 2611.050 1980.315 2611.330 1980.685 ;
        RECT 2611.050 1930.675 2611.330 1931.045 ;
        RECT 2611.120 1884.125 2611.260 1930.675 ;
        RECT 2611.050 1883.755 2611.330 1884.125 ;
        RECT 2611.050 1786.515 2611.330 1786.885 ;
        RECT 2611.120 1752.885 2611.260 1786.515 ;
        RECT 2611.050 1752.515 2611.330 1752.885 ;
        RECT 2611.050 1737.555 2611.330 1737.925 ;
        RECT 2611.120 1691.005 2611.260 1737.555 ;
        RECT 2611.050 1690.635 2611.330 1691.005 ;
        RECT 2611.050 1641.675 2611.330 1642.045 ;
        RECT 2611.120 1595.125 2611.260 1641.675 ;
        RECT 2611.050 1594.755 2611.330 1595.125 ;
        RECT 2611.050 1544.435 2611.330 1544.805 ;
        RECT 2611.120 1510.805 2611.260 1544.435 ;
        RECT 2611.050 1510.435 2611.330 1510.805 ;
        RECT 2611.050 1447.875 2611.330 1448.245 ;
        RECT 2611.120 1402.005 2611.260 1447.875 ;
        RECT 2611.050 1401.635 2611.330 1402.005 ;
        RECT 2611.050 1351.995 2611.330 1352.365 ;
        RECT 2611.120 1305.445 2611.260 1351.995 ;
        RECT 2611.050 1305.075 2611.330 1305.445 ;
        RECT 2611.050 1255.435 2611.330 1255.805 ;
        RECT 2611.120 1208.885 2611.260 1255.435 ;
        RECT 2611.050 1208.515 2611.330 1208.885 ;
        RECT 2611.050 1110.595 2611.330 1110.965 ;
        RECT 2611.120 1063.365 2611.260 1110.595 ;
        RECT 2611.050 1062.995 2611.330 1063.365 ;
        RECT 2611.050 1062.315 2611.330 1062.685 ;
        RECT 2611.120 1031.405 2611.260 1062.315 ;
        RECT 2611.050 1031.035 2611.330 1031.405 ;
        RECT 2607.830 999.755 2608.110 1000.125 ;
        RECT 2607.900 952.525 2608.040 999.755 ;
        RECT 2607.830 952.155 2608.110 952.525 ;
        RECT 2611.050 869.195 2611.330 869.565 ;
        RECT 2611.120 821.285 2611.260 869.195 ;
        RECT 2611.050 820.915 2611.330 821.285 ;
        RECT 2611.510 675.395 2611.790 675.765 ;
        RECT 2611.580 628.165 2611.720 675.395 ;
        RECT 2611.510 627.795 2611.790 628.165 ;
        RECT 2611.050 578.835 2611.330 579.205 ;
        RECT 2611.120 531.605 2611.260 578.835 ;
        RECT 2611.050 531.235 2611.330 531.605 ;
        RECT 1724.630 493.835 1724.910 494.205 ;
        RECT 1724.700 16.990 1724.840 493.835 ;
        RECT 1721.420 16.670 1721.680 16.990 ;
        RECT 1724.640 16.670 1724.900 16.990 ;
        RECT 1721.480 2.400 1721.620 16.670 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
      LAYER via2 ;
        RECT 2609.670 2897.680 2609.950 2897.960 ;
        RECT 2609.670 2850.760 2609.950 2851.040 ;
        RECT 2610.590 2801.120 2610.870 2801.400 ;
        RECT 2610.590 2753.520 2610.870 2753.800 ;
        RECT 2610.130 2704.560 2610.410 2704.840 ;
        RECT 2610.130 2657.640 2610.410 2657.920 ;
        RECT 2610.130 2608.000 2610.410 2608.280 ;
        RECT 2610.130 2561.080 2610.410 2561.360 ;
        RECT 2610.130 2511.440 2610.410 2511.720 ;
        RECT 2610.130 2463.160 2610.410 2463.440 ;
        RECT 2610.590 2316.960 2610.870 2317.240 ;
        RECT 2610.590 2270.040 2610.870 2270.320 ;
        RECT 2611.050 2124.520 2611.330 2124.800 ;
        RECT 2611.050 2076.920 2611.330 2077.200 ;
        RECT 2611.050 2027.280 2611.330 2027.560 ;
        RECT 2611.050 1980.360 2611.330 1980.640 ;
        RECT 2611.050 1930.720 2611.330 1931.000 ;
        RECT 2611.050 1883.800 2611.330 1884.080 ;
        RECT 2611.050 1786.560 2611.330 1786.840 ;
        RECT 2611.050 1752.560 2611.330 1752.840 ;
        RECT 2611.050 1737.600 2611.330 1737.880 ;
        RECT 2611.050 1690.680 2611.330 1690.960 ;
        RECT 2611.050 1641.720 2611.330 1642.000 ;
        RECT 2611.050 1594.800 2611.330 1595.080 ;
        RECT 2611.050 1544.480 2611.330 1544.760 ;
        RECT 2611.050 1510.480 2611.330 1510.760 ;
        RECT 2611.050 1447.920 2611.330 1448.200 ;
        RECT 2611.050 1401.680 2611.330 1401.960 ;
        RECT 2611.050 1352.040 2611.330 1352.320 ;
        RECT 2611.050 1305.120 2611.330 1305.400 ;
        RECT 2611.050 1255.480 2611.330 1255.760 ;
        RECT 2611.050 1208.560 2611.330 1208.840 ;
        RECT 2611.050 1110.640 2611.330 1110.920 ;
        RECT 2611.050 1063.040 2611.330 1063.320 ;
        RECT 2611.050 1062.360 2611.330 1062.640 ;
        RECT 2611.050 1031.080 2611.330 1031.360 ;
        RECT 2607.830 999.800 2608.110 1000.080 ;
        RECT 2607.830 952.200 2608.110 952.480 ;
        RECT 2611.050 869.240 2611.330 869.520 ;
        RECT 2611.050 820.960 2611.330 821.240 ;
        RECT 2611.510 675.440 2611.790 675.720 ;
        RECT 2611.510 627.840 2611.790 628.120 ;
        RECT 2611.050 578.880 2611.330 579.160 ;
        RECT 2611.050 531.280 2611.330 531.560 ;
        RECT 1724.630 493.880 1724.910 494.160 ;
      LAYER met3 ;
        RECT 2455.750 2999.970 2456.130 2999.980 ;
        RECT 2465.870 2999.970 2466.250 2999.980 ;
        RECT 2455.750 2999.670 2466.250 2999.970 ;
        RECT 2455.750 2999.660 2456.130 2999.670 ;
        RECT 2465.870 2999.660 2466.250 2999.670 ;
        RECT 2557.870 2990.450 2558.250 2990.460 ;
        RECT 2576.270 2990.450 2576.650 2990.460 ;
        RECT 2557.870 2990.150 2576.650 2990.450 ;
        RECT 2557.870 2990.140 2558.250 2990.150 ;
        RECT 2576.270 2990.140 2576.650 2990.150 ;
        RECT 2610.310 2960.530 2610.690 2960.540 ;
        RECT 2609.430 2960.230 2610.690 2960.530 ;
        RECT 2609.430 2959.180 2609.730 2960.230 ;
        RECT 2610.310 2960.220 2610.690 2960.230 ;
        RECT 2609.390 2958.860 2609.770 2959.180 ;
        RECT 2609.390 2911.940 2609.770 2912.260 ;
        RECT 2609.430 2910.890 2609.730 2911.940 ;
        RECT 2610.310 2910.890 2610.690 2910.900 ;
        RECT 2609.430 2910.590 2610.690 2910.890 ;
        RECT 2610.310 2910.580 2610.690 2910.590 ;
        RECT 2609.645 2897.970 2609.975 2897.985 ;
        RECT 2610.310 2897.970 2610.690 2897.980 ;
        RECT 2609.645 2897.670 2610.690 2897.970 ;
        RECT 2609.645 2897.655 2609.975 2897.670 ;
        RECT 2610.310 2897.660 2610.690 2897.670 ;
        RECT 2609.645 2851.050 2609.975 2851.065 ;
        RECT 2609.430 2850.735 2609.975 2851.050 ;
        RECT 2609.430 2850.380 2609.730 2850.735 ;
        RECT 2609.390 2850.060 2609.770 2850.380 ;
        RECT 2609.390 2815.380 2609.770 2815.700 ;
        RECT 2609.430 2814.330 2609.730 2815.380 ;
        RECT 2610.310 2814.330 2610.690 2814.340 ;
        RECT 2609.430 2814.030 2610.690 2814.330 ;
        RECT 2610.310 2814.020 2610.690 2814.030 ;
        RECT 2610.565 2801.420 2610.895 2801.425 ;
        RECT 2610.310 2801.410 2610.895 2801.420 ;
        RECT 2610.110 2801.110 2610.895 2801.410 ;
        RECT 2610.310 2801.100 2610.895 2801.110 ;
        RECT 2610.565 2801.095 2610.895 2801.100 ;
        RECT 2610.565 2753.810 2610.895 2753.825 ;
        RECT 2611.230 2753.810 2611.610 2753.820 ;
        RECT 2610.565 2753.510 2611.610 2753.810 ;
        RECT 2610.565 2753.495 2610.895 2753.510 ;
        RECT 2611.230 2753.500 2611.610 2753.510 ;
        RECT 2611.230 2719.810 2611.610 2719.820 ;
        RECT 2610.350 2719.510 2611.610 2719.810 ;
        RECT 2610.350 2718.460 2610.650 2719.510 ;
        RECT 2611.230 2719.500 2611.610 2719.510 ;
        RECT 2610.310 2718.140 2610.690 2718.460 ;
        RECT 2610.105 2704.860 2610.435 2704.865 ;
        RECT 2610.105 2704.850 2610.690 2704.860 ;
        RECT 2609.880 2704.550 2610.690 2704.850 ;
        RECT 2610.105 2704.540 2610.690 2704.550 ;
        RECT 2610.105 2704.535 2610.435 2704.540 ;
        RECT 2610.105 2657.930 2610.435 2657.945 ;
        RECT 2609.430 2657.630 2610.435 2657.930 ;
        RECT 2609.430 2657.260 2609.730 2657.630 ;
        RECT 2610.105 2657.615 2610.435 2657.630 ;
        RECT 2609.390 2656.940 2609.770 2657.260 ;
        RECT 2609.390 2622.260 2609.770 2622.580 ;
        RECT 2609.430 2621.210 2609.730 2622.260 ;
        RECT 2610.310 2621.210 2610.690 2621.220 ;
        RECT 2609.430 2620.910 2610.690 2621.210 ;
        RECT 2610.310 2620.900 2610.690 2620.910 ;
        RECT 2610.105 2608.300 2610.435 2608.305 ;
        RECT 2610.105 2608.290 2610.690 2608.300 ;
        RECT 2609.880 2607.990 2610.690 2608.290 ;
        RECT 2610.105 2607.980 2610.690 2607.990 ;
        RECT 2610.105 2607.975 2610.435 2607.980 ;
        RECT 2610.105 2561.370 2610.435 2561.385 ;
        RECT 2609.430 2561.070 2610.435 2561.370 ;
        RECT 2609.430 2560.700 2609.730 2561.070 ;
        RECT 2610.105 2561.055 2610.435 2561.070 ;
        RECT 2609.390 2560.380 2609.770 2560.700 ;
        RECT 2609.390 2526.010 2609.770 2526.020 ;
        RECT 2608.510 2525.710 2609.770 2526.010 ;
        RECT 2608.510 2524.660 2608.810 2525.710 ;
        RECT 2609.390 2525.700 2609.770 2525.710 ;
        RECT 2608.470 2524.340 2608.850 2524.660 ;
        RECT 2608.470 2511.730 2608.850 2511.740 ;
        RECT 2610.105 2511.730 2610.435 2511.745 ;
        RECT 2608.470 2511.430 2610.435 2511.730 ;
        RECT 2608.470 2511.420 2608.850 2511.430 ;
        RECT 2610.105 2511.415 2610.435 2511.430 ;
        RECT 2609.390 2463.450 2609.770 2463.460 ;
        RECT 2610.105 2463.450 2610.435 2463.465 ;
        RECT 2609.390 2463.150 2610.435 2463.450 ;
        RECT 2609.390 2463.140 2609.770 2463.150 ;
        RECT 2610.105 2463.135 2610.435 2463.150 ;
        RECT 2609.390 2429.450 2609.770 2429.460 ;
        RECT 2608.510 2429.150 2609.770 2429.450 ;
        RECT 2608.510 2428.100 2608.810 2429.150 ;
        RECT 2609.390 2429.140 2609.770 2429.150 ;
        RECT 2608.470 2427.780 2608.850 2428.100 ;
        RECT 2608.470 2380.490 2608.850 2380.500 ;
        RECT 2612.150 2380.490 2612.530 2380.500 ;
        RECT 2608.470 2380.190 2612.530 2380.490 ;
        RECT 2608.470 2380.180 2608.850 2380.190 ;
        RECT 2612.150 2380.180 2612.530 2380.190 ;
        RECT 2612.150 2332.890 2612.530 2332.900 ;
        RECT 2611.270 2332.590 2612.530 2332.890 ;
        RECT 2611.270 2331.540 2611.570 2332.590 ;
        RECT 2612.150 2332.580 2612.530 2332.590 ;
        RECT 2611.230 2331.220 2611.610 2331.540 ;
        RECT 2611.230 2317.620 2611.610 2317.940 ;
        RECT 2610.565 2317.250 2610.895 2317.265 ;
        RECT 2611.270 2317.250 2611.570 2317.620 ;
        RECT 2610.565 2316.950 2611.570 2317.250 ;
        RECT 2610.565 2316.935 2610.895 2316.950 ;
        RECT 2609.390 2270.330 2609.770 2270.340 ;
        RECT 2610.565 2270.330 2610.895 2270.345 ;
        RECT 2609.390 2270.030 2610.895 2270.330 ;
        RECT 2609.390 2270.020 2609.770 2270.030 ;
        RECT 2610.565 2270.015 2610.895 2270.030 ;
        RECT 2609.390 2236.020 2609.770 2236.340 ;
        RECT 2609.430 2234.970 2609.730 2236.020 ;
        RECT 2610.310 2234.970 2610.690 2234.980 ;
        RECT 2609.430 2234.670 2610.690 2234.970 ;
        RECT 2610.310 2234.660 2610.690 2234.670 ;
        RECT 2608.470 2187.370 2608.850 2187.380 ;
        RECT 2611.230 2187.370 2611.610 2187.380 ;
        RECT 2608.470 2187.070 2611.610 2187.370 ;
        RECT 2608.470 2187.060 2608.850 2187.070 ;
        RECT 2611.230 2187.060 2611.610 2187.070 ;
        RECT 2611.230 2139.770 2611.610 2139.780 ;
        RECT 2610.350 2139.470 2611.610 2139.770 ;
        RECT 2610.350 2138.420 2610.650 2139.470 ;
        RECT 2611.230 2139.460 2611.610 2139.470 ;
        RECT 2610.310 2138.100 2610.690 2138.420 ;
        RECT 2610.310 2124.810 2610.690 2124.820 ;
        RECT 2611.025 2124.810 2611.355 2124.825 ;
        RECT 2610.310 2124.510 2611.355 2124.810 ;
        RECT 2610.310 2124.500 2610.690 2124.510 ;
        RECT 2611.025 2124.495 2611.355 2124.510 ;
        RECT 2609.390 2077.210 2609.770 2077.220 ;
        RECT 2611.025 2077.210 2611.355 2077.225 ;
        RECT 2609.390 2076.910 2611.355 2077.210 ;
        RECT 2609.390 2076.900 2609.770 2076.910 ;
        RECT 2611.025 2076.895 2611.355 2076.910 ;
        RECT 2609.390 2043.210 2609.770 2043.220 ;
        RECT 2608.510 2042.910 2609.770 2043.210 ;
        RECT 2608.510 2041.860 2608.810 2042.910 ;
        RECT 2609.390 2042.900 2609.770 2042.910 ;
        RECT 2608.470 2041.540 2608.850 2041.860 ;
        RECT 2608.470 2027.940 2608.850 2028.260 ;
        RECT 2608.510 2027.570 2608.810 2027.940 ;
        RECT 2611.025 2027.570 2611.355 2027.585 ;
        RECT 2608.510 2027.270 2611.355 2027.570 ;
        RECT 2611.025 2027.255 2611.355 2027.270 ;
        RECT 2609.390 1980.650 2609.770 1980.660 ;
        RECT 2611.025 1980.650 2611.355 1980.665 ;
        RECT 2609.390 1980.350 2611.355 1980.650 ;
        RECT 2609.390 1980.340 2609.770 1980.350 ;
        RECT 2611.025 1980.335 2611.355 1980.350 ;
        RECT 2609.390 1946.340 2609.770 1946.660 ;
        RECT 2609.430 1945.290 2609.730 1946.340 ;
        RECT 2610.310 1945.290 2610.690 1945.300 ;
        RECT 2609.430 1944.990 2610.690 1945.290 ;
        RECT 2610.310 1944.980 2610.690 1944.990 ;
        RECT 2610.310 1931.380 2610.690 1931.700 ;
        RECT 2610.350 1931.010 2610.650 1931.380 ;
        RECT 2611.025 1931.010 2611.355 1931.025 ;
        RECT 2610.350 1930.710 2611.355 1931.010 ;
        RECT 2611.025 1930.695 2611.355 1930.710 ;
        RECT 2611.025 1884.100 2611.355 1884.105 ;
        RECT 2611.025 1884.090 2611.610 1884.100 ;
        RECT 2610.800 1883.790 2611.610 1884.090 ;
        RECT 2611.025 1883.780 2611.610 1883.790 ;
        RECT 2611.025 1883.775 2611.355 1883.780 ;
        RECT 2611.230 1850.090 2611.610 1850.100 ;
        RECT 2610.350 1849.790 2611.610 1850.090 ;
        RECT 2610.350 1848.740 2610.650 1849.790 ;
        RECT 2611.230 1849.780 2611.610 1849.790 ;
        RECT 2610.310 1848.420 2610.690 1848.740 ;
        RECT 2609.390 1786.850 2609.770 1786.860 ;
        RECT 2611.025 1786.850 2611.355 1786.865 ;
        RECT 2609.390 1786.550 2611.355 1786.850 ;
        RECT 2609.390 1786.540 2609.770 1786.550 ;
        RECT 2611.025 1786.535 2611.355 1786.550 ;
        RECT 2608.470 1752.850 2608.850 1752.860 ;
        RECT 2611.025 1752.850 2611.355 1752.865 ;
        RECT 2608.470 1752.550 2611.355 1752.850 ;
        RECT 2608.470 1752.540 2608.850 1752.550 ;
        RECT 2611.025 1752.535 2611.355 1752.550 ;
        RECT 2608.470 1738.260 2608.850 1738.580 ;
        RECT 2608.510 1737.890 2608.810 1738.260 ;
        RECT 2611.025 1737.890 2611.355 1737.905 ;
        RECT 2608.510 1737.590 2611.355 1737.890 ;
        RECT 2611.025 1737.575 2611.355 1737.590 ;
        RECT 2609.390 1690.970 2609.770 1690.980 ;
        RECT 2611.025 1690.970 2611.355 1690.985 ;
        RECT 2609.390 1690.670 2611.355 1690.970 ;
        RECT 2609.390 1690.660 2609.770 1690.670 ;
        RECT 2611.025 1690.655 2611.355 1690.670 ;
        RECT 2609.390 1656.660 2609.770 1656.980 ;
        RECT 2609.430 1655.610 2609.730 1656.660 ;
        RECT 2610.310 1655.610 2610.690 1655.620 ;
        RECT 2609.430 1655.310 2610.690 1655.610 ;
        RECT 2610.310 1655.300 2610.690 1655.310 ;
        RECT 2610.310 1642.010 2610.690 1642.020 ;
        RECT 2611.025 1642.010 2611.355 1642.025 ;
        RECT 2610.310 1641.710 2611.355 1642.010 ;
        RECT 2610.310 1641.700 2610.690 1641.710 ;
        RECT 2611.025 1641.695 2611.355 1641.710 ;
        RECT 2611.025 1595.090 2611.355 1595.105 ;
        RECT 2609.430 1594.790 2611.355 1595.090 ;
        RECT 2609.430 1594.420 2609.730 1594.790 ;
        RECT 2611.025 1594.775 2611.355 1594.790 ;
        RECT 2609.390 1594.100 2609.770 1594.420 ;
        RECT 2609.390 1560.100 2609.770 1560.420 ;
        RECT 2609.430 1559.050 2609.730 1560.100 ;
        RECT 2610.310 1559.050 2610.690 1559.060 ;
        RECT 2609.430 1558.750 2610.690 1559.050 ;
        RECT 2610.310 1558.740 2610.690 1558.750 ;
        RECT 2610.310 1545.140 2610.690 1545.460 ;
        RECT 2610.350 1544.770 2610.650 1545.140 ;
        RECT 2611.025 1544.770 2611.355 1544.785 ;
        RECT 2610.350 1544.470 2611.355 1544.770 ;
        RECT 2611.025 1544.455 2611.355 1544.470 ;
        RECT 2609.390 1510.770 2609.770 1510.780 ;
        RECT 2611.025 1510.770 2611.355 1510.785 ;
        RECT 2609.390 1510.470 2611.355 1510.770 ;
        RECT 2609.390 1510.460 2609.770 1510.470 ;
        RECT 2611.025 1510.455 2611.355 1510.470 ;
        RECT 2610.310 1448.580 2610.690 1448.900 ;
        RECT 2610.350 1448.210 2610.650 1448.580 ;
        RECT 2611.025 1448.210 2611.355 1448.225 ;
        RECT 2610.350 1447.910 2611.355 1448.210 ;
        RECT 2611.025 1447.895 2611.355 1447.910 ;
        RECT 2611.025 1401.970 2611.355 1401.985 ;
        RECT 2609.430 1401.670 2611.355 1401.970 ;
        RECT 2609.430 1401.300 2609.730 1401.670 ;
        RECT 2611.025 1401.655 2611.355 1401.670 ;
        RECT 2609.390 1400.980 2609.770 1401.300 ;
        RECT 2609.390 1366.980 2609.770 1367.300 ;
        RECT 2609.430 1365.250 2609.730 1366.980 ;
        RECT 2610.310 1365.250 2610.690 1365.260 ;
        RECT 2609.430 1364.950 2610.690 1365.250 ;
        RECT 2610.310 1364.940 2610.690 1364.950 ;
        RECT 2610.310 1352.330 2610.690 1352.340 ;
        RECT 2611.025 1352.330 2611.355 1352.345 ;
        RECT 2610.310 1352.030 2611.355 1352.330 ;
        RECT 2610.310 1352.020 2610.690 1352.030 ;
        RECT 2611.025 1352.015 2611.355 1352.030 ;
        RECT 2611.025 1305.410 2611.355 1305.425 ;
        RECT 2609.430 1305.110 2611.355 1305.410 ;
        RECT 2609.430 1304.740 2609.730 1305.110 ;
        RECT 2611.025 1305.095 2611.355 1305.110 ;
        RECT 2609.390 1304.420 2609.770 1304.740 ;
        RECT 2609.390 1269.740 2609.770 1270.060 ;
        RECT 2609.430 1268.690 2609.730 1269.740 ;
        RECT 2610.310 1268.690 2610.690 1268.700 ;
        RECT 2609.430 1268.390 2610.690 1268.690 ;
        RECT 2610.310 1268.380 2610.690 1268.390 ;
        RECT 2610.310 1255.770 2610.690 1255.780 ;
        RECT 2611.025 1255.770 2611.355 1255.785 ;
        RECT 2610.310 1255.470 2611.355 1255.770 ;
        RECT 2610.310 1255.460 2610.690 1255.470 ;
        RECT 2611.025 1255.455 2611.355 1255.470 ;
        RECT 2611.025 1208.850 2611.355 1208.865 ;
        RECT 2609.430 1208.550 2611.355 1208.850 ;
        RECT 2609.430 1208.180 2609.730 1208.550 ;
        RECT 2611.025 1208.535 2611.355 1208.550 ;
        RECT 2609.390 1207.860 2609.770 1208.180 ;
        RECT 2609.390 1173.180 2609.770 1173.500 ;
        RECT 2609.430 1172.130 2609.730 1173.180 ;
        RECT 2610.310 1172.130 2610.690 1172.140 ;
        RECT 2609.430 1171.830 2610.690 1172.130 ;
        RECT 2610.310 1171.820 2610.690 1171.830 ;
        RECT 2609.390 1110.930 2609.770 1110.940 ;
        RECT 2611.025 1110.930 2611.355 1110.945 ;
        RECT 2609.390 1110.630 2611.355 1110.930 ;
        RECT 2609.390 1110.620 2609.770 1110.630 ;
        RECT 2611.025 1110.615 2611.355 1110.630 ;
        RECT 2610.310 1063.330 2610.690 1063.340 ;
        RECT 2611.025 1063.330 2611.355 1063.345 ;
        RECT 2610.310 1063.030 2611.355 1063.330 ;
        RECT 2610.310 1063.020 2610.690 1063.030 ;
        RECT 2611.025 1063.015 2611.355 1063.030 ;
        RECT 2610.310 1062.650 2610.690 1062.660 ;
        RECT 2611.025 1062.650 2611.355 1062.665 ;
        RECT 2610.310 1062.350 2611.355 1062.650 ;
        RECT 2610.310 1062.340 2610.690 1062.350 ;
        RECT 2611.025 1062.335 2611.355 1062.350 ;
        RECT 2609.390 1031.370 2609.770 1031.380 ;
        RECT 2611.025 1031.370 2611.355 1031.385 ;
        RECT 2609.390 1031.070 2611.355 1031.370 ;
        RECT 2609.390 1031.060 2609.770 1031.070 ;
        RECT 2611.025 1031.055 2611.355 1031.070 ;
        RECT 2607.805 1000.090 2608.135 1000.105 ;
        RECT 2609.390 1000.090 2609.770 1000.100 ;
        RECT 2607.805 999.790 2609.770 1000.090 ;
        RECT 2607.805 999.775 2608.135 999.790 ;
        RECT 2609.390 999.780 2609.770 999.790 ;
        RECT 2607.805 952.490 2608.135 952.505 ;
        RECT 2608.470 952.490 2608.850 952.500 ;
        RECT 2607.805 952.190 2608.850 952.490 ;
        RECT 2607.805 952.175 2608.135 952.190 ;
        RECT 2608.470 952.180 2608.850 952.190 ;
        RECT 2609.390 883.810 2609.770 883.820 ;
        RECT 2608.510 883.510 2609.770 883.810 ;
        RECT 2608.510 882.460 2608.810 883.510 ;
        RECT 2609.390 883.500 2609.770 883.510 ;
        RECT 2608.470 882.140 2608.850 882.460 ;
        RECT 2608.470 869.530 2608.850 869.540 ;
        RECT 2611.025 869.530 2611.355 869.545 ;
        RECT 2608.470 869.230 2611.355 869.530 ;
        RECT 2608.470 869.220 2608.850 869.230 ;
        RECT 2611.025 869.215 2611.355 869.230 ;
        RECT 2609.390 821.250 2609.770 821.260 ;
        RECT 2611.025 821.250 2611.355 821.265 ;
        RECT 2609.390 820.950 2611.355 821.250 ;
        RECT 2609.390 820.940 2609.770 820.950 ;
        RECT 2611.025 820.935 2611.355 820.950 ;
        RECT 2609.390 787.250 2609.770 787.260 ;
        RECT 2608.510 786.950 2609.770 787.250 ;
        RECT 2608.510 785.900 2608.810 786.950 ;
        RECT 2609.390 786.940 2609.770 786.950 ;
        RECT 2608.470 785.580 2608.850 785.900 ;
        RECT 2608.470 738.290 2608.850 738.300 ;
        RECT 2612.150 738.290 2612.530 738.300 ;
        RECT 2608.470 737.990 2612.530 738.290 ;
        RECT 2608.470 737.980 2608.850 737.990 ;
        RECT 2612.150 737.980 2612.530 737.990 ;
        RECT 2612.150 690.690 2612.530 690.700 ;
        RECT 2611.270 690.390 2612.530 690.690 ;
        RECT 2611.270 689.340 2611.570 690.390 ;
        RECT 2612.150 690.380 2612.530 690.390 ;
        RECT 2611.230 689.020 2611.610 689.340 ;
        RECT 2611.485 675.740 2611.815 675.745 ;
        RECT 2611.230 675.730 2611.815 675.740 ;
        RECT 2611.230 675.430 2612.040 675.730 ;
        RECT 2611.230 675.420 2611.815 675.430 ;
        RECT 2611.485 675.415 2611.815 675.420 ;
        RECT 2609.390 628.130 2609.770 628.140 ;
        RECT 2611.485 628.130 2611.815 628.145 ;
        RECT 2609.390 627.830 2611.815 628.130 ;
        RECT 2609.390 627.820 2609.770 627.830 ;
        RECT 2611.485 627.815 2611.815 627.830 ;
        RECT 2609.390 593.820 2609.770 594.140 ;
        RECT 2609.430 592.770 2609.730 593.820 ;
        RECT 2610.310 592.770 2610.690 592.780 ;
        RECT 2609.430 592.470 2610.690 592.770 ;
        RECT 2610.310 592.460 2610.690 592.470 ;
        RECT 2610.310 579.170 2610.690 579.180 ;
        RECT 2611.025 579.170 2611.355 579.185 ;
        RECT 2610.310 578.870 2611.355 579.170 ;
        RECT 2610.310 578.860 2610.690 578.870 ;
        RECT 2611.025 578.855 2611.355 578.870 ;
        RECT 2609.390 531.570 2609.770 531.580 ;
        RECT 2611.025 531.570 2611.355 531.585 ;
        RECT 2609.390 531.270 2611.355 531.570 ;
        RECT 2609.390 531.260 2609.770 531.270 ;
        RECT 2611.025 531.255 2611.355 531.270 ;
        RECT 1724.605 494.170 1724.935 494.185 ;
        RECT 2609.390 494.170 2609.770 494.180 ;
        RECT 1724.605 493.870 2609.770 494.170 ;
        RECT 1724.605 493.855 1724.935 493.870 ;
        RECT 2609.390 493.860 2609.770 493.870 ;
      LAYER via3 ;
        RECT 2455.780 2999.660 2456.100 2999.980 ;
        RECT 2465.900 2999.660 2466.220 2999.980 ;
        RECT 2557.900 2990.140 2558.220 2990.460 ;
        RECT 2576.300 2990.140 2576.620 2990.460 ;
        RECT 2610.340 2960.220 2610.660 2960.540 ;
        RECT 2609.420 2958.860 2609.740 2959.180 ;
        RECT 2609.420 2911.940 2609.740 2912.260 ;
        RECT 2610.340 2910.580 2610.660 2910.900 ;
        RECT 2610.340 2897.660 2610.660 2897.980 ;
        RECT 2609.420 2850.060 2609.740 2850.380 ;
        RECT 2609.420 2815.380 2609.740 2815.700 ;
        RECT 2610.340 2814.020 2610.660 2814.340 ;
        RECT 2610.340 2801.100 2610.660 2801.420 ;
        RECT 2611.260 2753.500 2611.580 2753.820 ;
        RECT 2611.260 2719.500 2611.580 2719.820 ;
        RECT 2610.340 2718.140 2610.660 2718.460 ;
        RECT 2610.340 2704.540 2610.660 2704.860 ;
        RECT 2609.420 2656.940 2609.740 2657.260 ;
        RECT 2609.420 2622.260 2609.740 2622.580 ;
        RECT 2610.340 2620.900 2610.660 2621.220 ;
        RECT 2610.340 2607.980 2610.660 2608.300 ;
        RECT 2609.420 2560.380 2609.740 2560.700 ;
        RECT 2609.420 2525.700 2609.740 2526.020 ;
        RECT 2608.500 2524.340 2608.820 2524.660 ;
        RECT 2608.500 2511.420 2608.820 2511.740 ;
        RECT 2609.420 2463.140 2609.740 2463.460 ;
        RECT 2609.420 2429.140 2609.740 2429.460 ;
        RECT 2608.500 2427.780 2608.820 2428.100 ;
        RECT 2608.500 2380.180 2608.820 2380.500 ;
        RECT 2612.180 2380.180 2612.500 2380.500 ;
        RECT 2612.180 2332.580 2612.500 2332.900 ;
        RECT 2611.260 2331.220 2611.580 2331.540 ;
        RECT 2611.260 2317.620 2611.580 2317.940 ;
        RECT 2609.420 2270.020 2609.740 2270.340 ;
        RECT 2609.420 2236.020 2609.740 2236.340 ;
        RECT 2610.340 2234.660 2610.660 2234.980 ;
        RECT 2608.500 2187.060 2608.820 2187.380 ;
        RECT 2611.260 2187.060 2611.580 2187.380 ;
        RECT 2611.260 2139.460 2611.580 2139.780 ;
        RECT 2610.340 2138.100 2610.660 2138.420 ;
        RECT 2610.340 2124.500 2610.660 2124.820 ;
        RECT 2609.420 2076.900 2609.740 2077.220 ;
        RECT 2609.420 2042.900 2609.740 2043.220 ;
        RECT 2608.500 2041.540 2608.820 2041.860 ;
        RECT 2608.500 2027.940 2608.820 2028.260 ;
        RECT 2609.420 1980.340 2609.740 1980.660 ;
        RECT 2609.420 1946.340 2609.740 1946.660 ;
        RECT 2610.340 1944.980 2610.660 1945.300 ;
        RECT 2610.340 1931.380 2610.660 1931.700 ;
        RECT 2611.260 1883.780 2611.580 1884.100 ;
        RECT 2611.260 1849.780 2611.580 1850.100 ;
        RECT 2610.340 1848.420 2610.660 1848.740 ;
        RECT 2609.420 1786.540 2609.740 1786.860 ;
        RECT 2608.500 1752.540 2608.820 1752.860 ;
        RECT 2608.500 1738.260 2608.820 1738.580 ;
        RECT 2609.420 1690.660 2609.740 1690.980 ;
        RECT 2609.420 1656.660 2609.740 1656.980 ;
        RECT 2610.340 1655.300 2610.660 1655.620 ;
        RECT 2610.340 1641.700 2610.660 1642.020 ;
        RECT 2609.420 1594.100 2609.740 1594.420 ;
        RECT 2609.420 1560.100 2609.740 1560.420 ;
        RECT 2610.340 1558.740 2610.660 1559.060 ;
        RECT 2610.340 1545.140 2610.660 1545.460 ;
        RECT 2609.420 1510.460 2609.740 1510.780 ;
        RECT 2610.340 1448.580 2610.660 1448.900 ;
        RECT 2609.420 1400.980 2609.740 1401.300 ;
        RECT 2609.420 1366.980 2609.740 1367.300 ;
        RECT 2610.340 1364.940 2610.660 1365.260 ;
        RECT 2610.340 1352.020 2610.660 1352.340 ;
        RECT 2609.420 1304.420 2609.740 1304.740 ;
        RECT 2609.420 1269.740 2609.740 1270.060 ;
        RECT 2610.340 1268.380 2610.660 1268.700 ;
        RECT 2610.340 1255.460 2610.660 1255.780 ;
        RECT 2609.420 1207.860 2609.740 1208.180 ;
        RECT 2609.420 1173.180 2609.740 1173.500 ;
        RECT 2610.340 1171.820 2610.660 1172.140 ;
        RECT 2609.420 1110.620 2609.740 1110.940 ;
        RECT 2610.340 1063.020 2610.660 1063.340 ;
        RECT 2610.340 1062.340 2610.660 1062.660 ;
        RECT 2609.420 1031.060 2609.740 1031.380 ;
        RECT 2609.420 999.780 2609.740 1000.100 ;
        RECT 2608.500 952.180 2608.820 952.500 ;
        RECT 2609.420 883.500 2609.740 883.820 ;
        RECT 2608.500 882.140 2608.820 882.460 ;
        RECT 2608.500 869.220 2608.820 869.540 ;
        RECT 2609.420 820.940 2609.740 821.260 ;
        RECT 2609.420 786.940 2609.740 787.260 ;
        RECT 2608.500 785.580 2608.820 785.900 ;
        RECT 2608.500 737.980 2608.820 738.300 ;
        RECT 2612.180 737.980 2612.500 738.300 ;
        RECT 2612.180 690.380 2612.500 690.700 ;
        RECT 2611.260 689.020 2611.580 689.340 ;
        RECT 2611.260 675.420 2611.580 675.740 ;
        RECT 2609.420 627.820 2609.740 628.140 ;
        RECT 2609.420 593.820 2609.740 594.140 ;
        RECT 2610.340 592.460 2610.660 592.780 ;
        RECT 2610.340 578.860 2610.660 579.180 ;
        RECT 2609.420 531.260 2609.740 531.580 ;
        RECT 2609.420 493.860 2609.740 494.180 ;
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 3010.000 475.020 3538.100 ;
        RECT 652.020 3010.000 655.020 3538.100 ;
        RECT 832.020 3010.000 835.020 3538.100 ;
        RECT 1012.020 3010.000 1015.020 3538.100 ;
        RECT 1192.020 3010.000 1195.020 3538.100 ;
        RECT 1372.020 3010.000 1375.020 3538.100 ;
        RECT 1552.020 3010.000 1555.020 3538.100 ;
        RECT 1732.020 3010.000 1735.020 3538.100 ;
        RECT 1912.020 3010.000 1915.020 3538.100 ;
        RECT 2092.020 3010.000 2095.020 3538.100 ;
        RECT 2272.020 3010.000 2275.020 3538.100 ;
        RECT 2452.020 3010.000 2455.020 3538.100 ;
        RECT 2455.775 2999.655 2456.105 2999.985 ;
        RECT 2465.895 2999.655 2466.225 2999.985 ;
        RECT 2024.790 2996.510 2025.970 2997.690 ;
        RECT 2455.790 2990.890 2456.090 2999.655 ;
        RECT 2465.910 2994.290 2466.210 2999.655 ;
        RECT 2465.470 2993.110 2466.650 2994.290 ;
        RECT 2455.350 2989.710 2456.530 2990.890 ;
        RECT 2557.470 2989.710 2558.650 2990.890 ;
        RECT 2575.870 2989.710 2577.050 2990.890 ;
        RECT 2609.910 2989.710 2611.090 2990.890 ;
        RECT 2610.350 2960.545 2610.650 2989.710 ;
        RECT 2610.335 2960.215 2610.665 2960.545 ;
        RECT 2609.415 2958.855 2609.745 2959.185 ;
        RECT 2609.430 2912.265 2609.730 2958.855 ;
        RECT 2609.415 2911.935 2609.745 2912.265 ;
        RECT 2610.335 2910.575 2610.665 2910.905 ;
        RECT 2610.350 2897.985 2610.650 2910.575 ;
        RECT 2610.335 2897.655 2610.665 2897.985 ;
        RECT 2609.415 2850.055 2609.745 2850.385 ;
        RECT 2609.430 2815.705 2609.730 2850.055 ;
        RECT 2609.415 2815.375 2609.745 2815.705 ;
        RECT 2610.335 2814.015 2610.665 2814.345 ;
        RECT 2610.350 2801.425 2610.650 2814.015 ;
        RECT 2610.335 2801.095 2610.665 2801.425 ;
        RECT 2611.255 2753.495 2611.585 2753.825 ;
        RECT 2611.270 2719.825 2611.570 2753.495 ;
        RECT 2611.255 2719.495 2611.585 2719.825 ;
        RECT 2610.335 2718.135 2610.665 2718.465 ;
        RECT 2610.350 2704.865 2610.650 2718.135 ;
        RECT 2610.335 2704.535 2610.665 2704.865 ;
        RECT 2609.415 2656.935 2609.745 2657.265 ;
        RECT 2609.430 2622.585 2609.730 2656.935 ;
        RECT 2609.415 2622.255 2609.745 2622.585 ;
        RECT 2610.335 2620.895 2610.665 2621.225 ;
        RECT 2610.350 2608.305 2610.650 2620.895 ;
        RECT 2610.335 2607.975 2610.665 2608.305 ;
        RECT 2609.415 2560.375 2609.745 2560.705 ;
        RECT 2609.430 2526.025 2609.730 2560.375 ;
        RECT 2609.415 2525.695 2609.745 2526.025 ;
        RECT 2608.495 2524.335 2608.825 2524.665 ;
        RECT 2608.510 2511.745 2608.810 2524.335 ;
        RECT 2608.495 2511.415 2608.825 2511.745 ;
        RECT 2609.415 2463.135 2609.745 2463.465 ;
        RECT 2609.430 2429.465 2609.730 2463.135 ;
        RECT 2609.415 2429.135 2609.745 2429.465 ;
        RECT 2608.495 2427.775 2608.825 2428.105 ;
        RECT 2608.510 2380.505 2608.810 2427.775 ;
        RECT 2608.495 2380.175 2608.825 2380.505 ;
        RECT 2612.175 2380.175 2612.505 2380.505 ;
        RECT 2612.190 2332.905 2612.490 2380.175 ;
        RECT 2612.175 2332.575 2612.505 2332.905 ;
        RECT 2611.255 2331.215 2611.585 2331.545 ;
        RECT 2611.270 2317.945 2611.570 2331.215 ;
        RECT 2611.255 2317.615 2611.585 2317.945 ;
        RECT 2609.415 2270.015 2609.745 2270.345 ;
        RECT 2609.430 2236.345 2609.730 2270.015 ;
        RECT 2609.415 2236.015 2609.745 2236.345 ;
        RECT 2610.335 2234.655 2610.665 2234.985 ;
        RECT 2610.350 2188.050 2610.650 2234.655 ;
        RECT 2608.510 2187.750 2610.650 2188.050 ;
        RECT 2608.510 2187.385 2608.810 2187.750 ;
        RECT 2608.495 2187.055 2608.825 2187.385 ;
        RECT 2611.255 2187.055 2611.585 2187.385 ;
        RECT 2611.270 2139.785 2611.570 2187.055 ;
        RECT 2611.255 2139.455 2611.585 2139.785 ;
        RECT 2610.335 2138.095 2610.665 2138.425 ;
        RECT 2610.350 2124.825 2610.650 2138.095 ;
        RECT 2610.335 2124.495 2610.665 2124.825 ;
        RECT 2609.415 2076.895 2609.745 2077.225 ;
        RECT 2609.430 2043.225 2609.730 2076.895 ;
        RECT 2609.415 2042.895 2609.745 2043.225 ;
        RECT 2608.495 2041.535 2608.825 2041.865 ;
        RECT 2608.510 2028.265 2608.810 2041.535 ;
        RECT 2608.495 2027.935 2608.825 2028.265 ;
        RECT 2609.415 1980.335 2609.745 1980.665 ;
        RECT 2609.430 1946.665 2609.730 1980.335 ;
        RECT 2609.415 1946.335 2609.745 1946.665 ;
        RECT 2610.335 1944.975 2610.665 1945.305 ;
        RECT 2610.350 1931.705 2610.650 1944.975 ;
        RECT 2610.335 1931.375 2610.665 1931.705 ;
        RECT 2611.255 1883.775 2611.585 1884.105 ;
        RECT 2611.270 1850.105 2611.570 1883.775 ;
        RECT 2611.255 1849.775 2611.585 1850.105 ;
        RECT 2610.335 1848.415 2610.665 1848.745 ;
        RECT 2610.350 1800.450 2610.650 1848.415 ;
        RECT 2609.430 1800.150 2610.650 1800.450 ;
        RECT 2609.430 1786.865 2609.730 1800.150 ;
        RECT 2609.415 1786.535 2609.745 1786.865 ;
        RECT 2608.495 1752.535 2608.825 1752.865 ;
        RECT 2608.510 1738.585 2608.810 1752.535 ;
        RECT 2608.495 1738.255 2608.825 1738.585 ;
        RECT 2609.415 1690.655 2609.745 1690.985 ;
        RECT 2609.430 1656.985 2609.730 1690.655 ;
        RECT 2609.415 1656.655 2609.745 1656.985 ;
        RECT 2610.335 1655.295 2610.665 1655.625 ;
        RECT 2610.350 1642.025 2610.650 1655.295 ;
        RECT 2610.335 1641.695 2610.665 1642.025 ;
        RECT 2609.415 1594.095 2609.745 1594.425 ;
        RECT 2609.430 1560.425 2609.730 1594.095 ;
        RECT 2609.415 1560.095 2609.745 1560.425 ;
        RECT 2610.335 1558.735 2610.665 1559.065 ;
        RECT 2610.350 1545.465 2610.650 1558.735 ;
        RECT 2610.335 1545.135 2610.665 1545.465 ;
        RECT 2609.415 1510.455 2609.745 1510.785 ;
        RECT 2609.430 1463.850 2609.730 1510.455 ;
        RECT 2609.430 1463.550 2610.650 1463.850 ;
        RECT 2610.350 1448.905 2610.650 1463.550 ;
        RECT 2610.335 1448.575 2610.665 1448.905 ;
        RECT 2609.415 1400.975 2609.745 1401.305 ;
        RECT 2609.430 1367.305 2609.730 1400.975 ;
        RECT 2609.415 1366.975 2609.745 1367.305 ;
        RECT 2610.335 1364.935 2610.665 1365.265 ;
        RECT 2610.350 1352.345 2610.650 1364.935 ;
        RECT 2610.335 1352.015 2610.665 1352.345 ;
        RECT 2609.415 1304.415 2609.745 1304.745 ;
        RECT 2609.430 1270.065 2609.730 1304.415 ;
        RECT 2609.415 1269.735 2609.745 1270.065 ;
        RECT 2610.335 1268.375 2610.665 1268.705 ;
        RECT 2610.350 1255.785 2610.650 1268.375 ;
        RECT 2610.335 1255.455 2610.665 1255.785 ;
        RECT 2609.415 1207.855 2609.745 1208.185 ;
        RECT 2609.430 1173.505 2609.730 1207.855 ;
        RECT 2609.415 1173.175 2609.745 1173.505 ;
        RECT 2610.335 1171.815 2610.665 1172.145 ;
        RECT 2610.350 1137.450 2610.650 1171.815 ;
        RECT 2607.590 1137.150 2610.650 1137.450 ;
        RECT 2607.590 1123.850 2607.890 1137.150 ;
        RECT 2607.590 1123.550 2609.730 1123.850 ;
        RECT 2609.430 1110.945 2609.730 1123.550 ;
        RECT 2609.415 1110.615 2609.745 1110.945 ;
        RECT 2610.335 1063.015 2610.665 1063.345 ;
        RECT 2610.350 1062.665 2610.650 1063.015 ;
        RECT 2610.335 1062.335 2610.665 1062.665 ;
        RECT 2609.415 1031.055 2609.745 1031.385 ;
        RECT 2609.430 1000.105 2609.730 1031.055 ;
        RECT 2609.415 999.775 2609.745 1000.105 ;
        RECT 2608.495 952.175 2608.825 952.505 ;
        RECT 2608.510 930.050 2608.810 952.175 ;
        RECT 2608.510 929.750 2609.730 930.050 ;
        RECT 2609.430 883.825 2609.730 929.750 ;
        RECT 2609.415 883.495 2609.745 883.825 ;
        RECT 2608.495 882.135 2608.825 882.465 ;
        RECT 2608.510 869.545 2608.810 882.135 ;
        RECT 2608.495 869.215 2608.825 869.545 ;
        RECT 2609.415 820.935 2609.745 821.265 ;
        RECT 2609.430 787.265 2609.730 820.935 ;
        RECT 2609.415 786.935 2609.745 787.265 ;
        RECT 2608.495 785.575 2608.825 785.905 ;
        RECT 2608.510 738.305 2608.810 785.575 ;
        RECT 2608.495 737.975 2608.825 738.305 ;
        RECT 2612.175 737.975 2612.505 738.305 ;
        RECT 2612.190 690.705 2612.490 737.975 ;
        RECT 2612.175 690.375 2612.505 690.705 ;
        RECT 2611.255 689.015 2611.585 689.345 ;
        RECT 2611.270 675.745 2611.570 689.015 ;
        RECT 2611.255 675.415 2611.585 675.745 ;
        RECT 2609.415 627.815 2609.745 628.145 ;
        RECT 2609.430 594.145 2609.730 627.815 ;
        RECT 2609.415 593.815 2609.745 594.145 ;
        RECT 2610.335 592.455 2610.665 592.785 ;
        RECT 2610.350 579.185 2610.650 592.455 ;
        RECT 2610.335 578.855 2610.665 579.185 ;
        RECT 2609.415 531.255 2609.745 531.585 ;
        RECT 472.020 -18.420 475.020 510.000 ;
        RECT 652.020 -18.420 655.020 510.000 ;
        RECT 832.020 -18.420 835.020 510.000 ;
        RECT 1012.020 -18.420 1015.020 510.000 ;
        RECT 1192.020 -18.420 1195.020 510.000 ;
        RECT 1372.020 -18.420 1375.020 510.000 ;
        RECT 1552.020 -18.420 1555.020 510.000 ;
        RECT 1732.020 -18.420 1735.020 510.000 ;
        RECT 1912.020 -18.420 1915.020 510.000 ;
        RECT 2092.020 -18.420 2095.020 510.000 ;
        RECT 2272.020 -18.420 2275.020 510.000 ;
        RECT 2452.020 -18.420 2455.020 510.000 ;
        RECT 2609.430 494.185 2609.730 531.255 ;
        RECT 2609.415 493.855 2609.745 494.185 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 2024.580 2995.400 2026.180 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT 2023.660 2994.500 2026.180 2995.400 ;
        RECT 2023.660 2992.900 2103.460 2994.500 ;
        RECT 2101.860 2991.100 2103.460 2992.900 ;
        RECT 2122.100 2992.900 2131.060 2994.500 ;
        RECT 2465.260 2992.900 2486.180 2994.500 ;
        RECT 2101.860 2989.500 2111.740 2991.100 ;
        RECT 2110.140 2987.700 2111.740 2989.500 ;
        RECT 2122.100 2987.700 2123.700 2992.900 ;
        RECT 2129.460 2991.100 2131.060 2992.900 ;
        RECT 2484.580 2991.100 2486.180 2992.900 ;
        RECT 2129.460 2989.500 2456.740 2991.100 ;
        RECT 2484.580 2989.500 2558.860 2991.100 ;
        RECT 2575.660 2989.500 2611.300 2991.100 ;
        RECT 2110.140 2986.100 2123.700 2987.700 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.710 704.040 2523.030 704.100 ;
        RECT 2542.030 704.040 2542.350 704.100 ;
        RECT 2522.710 703.900 2542.350 704.040 ;
        RECT 2522.710 703.840 2523.030 703.900 ;
        RECT 2542.030 703.840 2542.350 703.900 ;
        RECT 1745.310 481.000 1745.630 481.060 ;
        RECT 2542.030 481.000 2542.350 481.060 ;
        RECT 1745.310 480.860 2542.350 481.000 ;
        RECT 1745.310 480.800 1745.630 480.860 ;
        RECT 2542.030 480.800 2542.350 480.860 ;
        RECT 1739.330 15.200 1739.650 15.260 ;
        RECT 1745.310 15.200 1745.630 15.260 ;
        RECT 1739.330 15.060 1745.630 15.200 ;
        RECT 1739.330 15.000 1739.650 15.060 ;
        RECT 1745.310 15.000 1745.630 15.060 ;
      LAYER via ;
        RECT 2522.740 703.840 2523.000 704.100 ;
        RECT 2542.060 703.840 2542.320 704.100 ;
        RECT 1745.340 480.800 1745.600 481.060 ;
        RECT 2542.060 480.800 2542.320 481.060 ;
        RECT 1739.360 15.000 1739.620 15.260 ;
        RECT 1745.340 15.000 1745.600 15.260 ;
      LAYER met2 ;
        RECT 2522.730 704.635 2523.010 705.005 ;
        RECT 2522.800 704.130 2522.940 704.635 ;
        RECT 2522.740 703.810 2523.000 704.130 ;
        RECT 2542.060 703.810 2542.320 704.130 ;
        RECT 2542.120 481.090 2542.260 703.810 ;
        RECT 1745.340 480.770 1745.600 481.090 ;
        RECT 2542.060 480.770 2542.320 481.090 ;
        RECT 1745.400 15.290 1745.540 480.770 ;
        RECT 1739.360 14.970 1739.620 15.290 ;
        RECT 1745.340 14.970 1745.600 15.290 ;
        RECT 1739.420 2.400 1739.560 14.970 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
      LAYER via2 ;
        RECT 2522.730 704.680 2523.010 704.960 ;
      LAYER met3 ;
        RECT 2506.000 704.970 2510.000 705.120 ;
        RECT 2522.705 704.970 2523.035 704.985 ;
        RECT 2506.000 704.670 2523.035 704.970 ;
        RECT 2506.000 704.520 2510.000 704.670 ;
        RECT 2522.705 704.655 2523.035 704.670 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.630 280.060 407.950 280.120 ;
        RECT 1753.130 280.060 1753.450 280.120 ;
        RECT 407.630 279.920 1753.450 280.060 ;
        RECT 407.630 279.860 407.950 279.920 ;
        RECT 1753.130 279.860 1753.450 279.920 ;
        RECT 1753.130 62.120 1753.450 62.180 ;
        RECT 1756.810 62.120 1757.130 62.180 ;
        RECT 1753.130 61.980 1757.130 62.120 ;
        RECT 1753.130 61.920 1753.450 61.980 ;
        RECT 1756.810 61.920 1757.130 61.980 ;
      LAYER via ;
        RECT 407.660 279.860 407.920 280.120 ;
        RECT 1753.160 279.860 1753.420 280.120 ;
        RECT 1753.160 61.920 1753.420 62.180 ;
        RECT 1756.840 61.920 1757.100 62.180 ;
      LAYER met2 ;
        RECT 407.650 2046.955 407.930 2047.325 ;
        RECT 407.720 280.150 407.860 2046.955 ;
        RECT 407.660 279.830 407.920 280.150 ;
        RECT 1753.160 279.830 1753.420 280.150 ;
        RECT 1753.220 62.210 1753.360 279.830 ;
        RECT 1753.160 61.890 1753.420 62.210 ;
        RECT 1756.840 61.890 1757.100 62.210 ;
        RECT 1756.900 2.400 1757.040 61.890 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
      LAYER via2 ;
        RECT 407.650 2047.000 407.930 2047.280 ;
      LAYER met3 ;
        RECT 407.625 2047.290 407.955 2047.305 ;
        RECT 410.000 2047.290 414.000 2047.440 ;
        RECT 407.625 2046.990 414.000 2047.290 ;
        RECT 407.625 2046.975 407.955 2046.990 ;
        RECT 410.000 2046.840 414.000 2046.990 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1950.930 3031.340 1951.250 3031.400 ;
        RECT 2602.750 3031.340 2603.070 3031.400 ;
        RECT 1950.930 3031.200 2603.070 3031.340 ;
        RECT 1950.930 3031.140 1951.250 3031.200 ;
        RECT 2602.750 3031.140 2603.070 3031.200 ;
        RECT 1779.810 486.780 1780.130 486.840 ;
        RECT 2602.750 486.780 2603.070 486.840 ;
        RECT 1779.810 486.640 2603.070 486.780 ;
        RECT 1779.810 486.580 1780.130 486.640 ;
        RECT 2602.750 486.580 2603.070 486.640 ;
        RECT 1774.750 15.880 1775.070 15.940 ;
        RECT 1779.810 15.880 1780.130 15.940 ;
        RECT 1774.750 15.740 1780.130 15.880 ;
        RECT 1774.750 15.680 1775.070 15.740 ;
        RECT 1779.810 15.680 1780.130 15.740 ;
      LAYER via ;
        RECT 1950.960 3031.140 1951.220 3031.400 ;
        RECT 2602.780 3031.140 2603.040 3031.400 ;
        RECT 1779.840 486.580 1780.100 486.840 ;
        RECT 2602.780 486.580 2603.040 486.840 ;
        RECT 1774.780 15.680 1775.040 15.940 ;
        RECT 1779.840 15.680 1780.100 15.940 ;
      LAYER met2 ;
        RECT 1950.960 3031.110 1951.220 3031.430 ;
        RECT 2602.780 3031.110 2603.040 3031.430 ;
        RECT 1951.020 3010.000 1951.160 3031.110 ;
        RECT 1951.020 3009.340 1951.370 3010.000 ;
        RECT 1951.090 3006.000 1951.370 3009.340 ;
        RECT 2602.840 486.870 2602.980 3031.110 ;
        RECT 1779.840 486.550 1780.100 486.870 ;
        RECT 2602.780 486.550 2603.040 486.870 ;
        RECT 1779.900 15.970 1780.040 486.550 ;
        RECT 1774.780 15.650 1775.040 15.970 ;
        RECT 1779.840 15.650 1780.100 15.970 ;
        RECT 1774.840 2.400 1774.980 15.650 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 356.110 911.100 356.430 911.160 ;
        RECT 393.370 911.100 393.690 911.160 ;
        RECT 356.110 910.960 393.690 911.100 ;
        RECT 356.110 910.900 356.430 910.960 ;
        RECT 393.370 910.900 393.690 910.960 ;
        RECT 356.110 44.780 356.430 44.840 ;
        RECT 1792.690 44.780 1793.010 44.840 ;
        RECT 356.110 44.640 1793.010 44.780 ;
        RECT 356.110 44.580 356.430 44.640 ;
        RECT 1792.690 44.580 1793.010 44.640 ;
      LAYER via ;
        RECT 356.140 910.900 356.400 911.160 ;
        RECT 393.400 910.900 393.660 911.160 ;
        RECT 356.140 44.580 356.400 44.840 ;
        RECT 1792.720 44.580 1792.980 44.840 ;
      LAYER met2 ;
        RECT 393.390 915.435 393.670 915.805 ;
        RECT 393.460 911.190 393.600 915.435 ;
        RECT 356.140 910.870 356.400 911.190 ;
        RECT 393.400 910.870 393.660 911.190 ;
        RECT 356.200 44.870 356.340 910.870 ;
        RECT 356.140 44.550 356.400 44.870 ;
        RECT 1792.720 44.550 1792.980 44.870 ;
        RECT 1792.780 2.400 1792.920 44.550 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
      LAYER via2 ;
        RECT 393.390 915.480 393.670 915.760 ;
      LAYER met3 ;
        RECT 393.365 915.770 393.695 915.785 ;
        RECT 410.000 915.770 414.000 915.920 ;
        RECT 393.365 915.470 414.000 915.770 ;
        RECT 393.365 915.455 393.695 915.470 ;
        RECT 410.000 915.320 414.000 915.470 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.870 16.900 1808.190 16.960 ;
        RECT 1810.630 16.900 1810.950 16.960 ;
        RECT 1807.870 16.760 1810.950 16.900 ;
        RECT 1807.870 16.700 1808.190 16.760 ;
        RECT 1810.630 16.700 1810.950 16.760 ;
      LAYER via ;
        RECT 1807.900 16.700 1808.160 16.960 ;
        RECT 1810.660 16.700 1810.920 16.960 ;
      LAYER met2 ;
        RECT 1808.490 510.410 1808.770 514.000 ;
        RECT 1807.960 510.270 1808.770 510.410 ;
        RECT 1807.960 16.990 1808.100 510.270 ;
        RECT 1808.490 510.000 1808.770 510.270 ;
        RECT 1807.900 16.670 1808.160 16.990 ;
        RECT 1810.660 16.670 1810.920 16.990 ;
        RECT 1810.720 2.400 1810.860 16.670 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.010 472.840 1835.330 472.900 ;
        RECT 2507.990 472.840 2508.310 472.900 ;
        RECT 1835.010 472.700 2508.310 472.840 ;
        RECT 1835.010 472.640 1835.330 472.700 ;
        RECT 2507.990 472.640 2508.310 472.700 ;
        RECT 1828.570 16.220 1828.890 16.280 ;
        RECT 1835.010 16.220 1835.330 16.280 ;
        RECT 1828.570 16.080 1835.330 16.220 ;
        RECT 1828.570 16.020 1828.890 16.080 ;
        RECT 1835.010 16.020 1835.330 16.080 ;
      LAYER via ;
        RECT 1835.040 472.640 1835.300 472.900 ;
        RECT 2508.020 472.640 2508.280 472.900 ;
        RECT 1828.600 16.020 1828.860 16.280 ;
        RECT 1835.040 16.020 1835.300 16.280 ;
      LAYER met2 ;
        RECT 2508.010 1541.035 2508.290 1541.405 ;
        RECT 2508.080 472.930 2508.220 1541.035 ;
        RECT 1835.040 472.610 1835.300 472.930 ;
        RECT 2508.020 472.610 2508.280 472.930 ;
        RECT 1835.100 16.310 1835.240 472.610 ;
        RECT 1828.600 15.990 1828.860 16.310 ;
        RECT 1835.040 15.990 1835.300 16.310 ;
        RECT 1828.660 2.400 1828.800 15.990 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 2508.010 1541.080 2508.290 1541.360 ;
      LAYER met3 ;
        RECT 2506.000 1543.640 2510.000 1544.240 ;
        RECT 2508.230 1541.385 2508.530 1543.640 ;
        RECT 2507.985 1541.070 2508.530 1541.385 ;
        RECT 2507.985 1541.055 2508.315 1541.070 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 2829.380 234.530 2829.440 ;
        RECT 393.370 2829.380 393.690 2829.440 ;
        RECT 234.210 2829.240 393.690 2829.380 ;
        RECT 234.210 2829.180 234.530 2829.240 ;
        RECT 393.370 2829.180 393.690 2829.240 ;
      LAYER via ;
        RECT 234.240 2829.180 234.500 2829.440 ;
        RECT 393.400 2829.180 393.660 2829.440 ;
      LAYER met2 ;
        RECT 393.390 2833.035 393.670 2833.405 ;
        RECT 393.460 2829.470 393.600 2833.035 ;
        RECT 234.240 2829.150 234.500 2829.470 ;
        RECT 393.400 2829.150 393.660 2829.470 ;
        RECT 234.300 45.405 234.440 2829.150 ;
        RECT 234.230 45.035 234.510 45.405 ;
        RECT 1846.070 45.035 1846.350 45.405 ;
        RECT 1846.140 2.400 1846.280 45.035 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 393.390 2833.080 393.670 2833.360 ;
        RECT 234.230 45.080 234.510 45.360 ;
        RECT 1846.070 45.080 1846.350 45.360 ;
      LAYER met3 ;
        RECT 393.365 2833.370 393.695 2833.385 ;
        RECT 410.000 2833.370 414.000 2833.520 ;
        RECT 393.365 2833.070 414.000 2833.370 ;
        RECT 393.365 2833.055 393.695 2833.070 ;
        RECT 410.000 2832.920 414.000 2833.070 ;
        RECT 234.205 45.370 234.535 45.385 ;
        RECT 1846.045 45.370 1846.375 45.385 ;
        RECT 234.205 45.070 1846.375 45.370 ;
        RECT 234.205 45.055 234.535 45.070 ;
        RECT 1846.045 45.055 1846.375 45.070 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 307.810 2394.520 308.130 2394.580 ;
        RECT 393.370 2394.520 393.690 2394.580 ;
        RECT 307.810 2394.380 393.690 2394.520 ;
        RECT 307.810 2394.320 308.130 2394.380 ;
        RECT 393.370 2394.320 393.690 2394.380 ;
        RECT 307.810 60.420 308.130 60.480 ;
        RECT 1863.070 60.420 1863.390 60.480 ;
        RECT 307.810 60.280 1863.390 60.420 ;
        RECT 307.810 60.220 308.130 60.280 ;
        RECT 1863.070 60.220 1863.390 60.280 ;
      LAYER via ;
        RECT 307.840 2394.320 308.100 2394.580 ;
        RECT 393.400 2394.320 393.660 2394.580 ;
        RECT 307.840 60.220 308.100 60.480 ;
        RECT 1863.100 60.220 1863.360 60.480 ;
      LAYER met2 ;
        RECT 393.390 2395.115 393.670 2395.485 ;
        RECT 393.460 2394.610 393.600 2395.115 ;
        RECT 307.840 2394.290 308.100 2394.610 ;
        RECT 393.400 2394.290 393.660 2394.610 ;
        RECT 307.900 60.510 308.040 2394.290 ;
        RECT 307.840 60.190 308.100 60.510 ;
        RECT 1863.100 60.190 1863.360 60.510 ;
        RECT 1863.160 17.410 1863.300 60.190 ;
        RECT 1863.160 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 393.390 2395.160 393.670 2395.440 ;
      LAYER met3 ;
        RECT 393.365 2395.450 393.695 2395.465 ;
        RECT 410.000 2395.450 414.000 2395.600 ;
        RECT 393.365 2395.150 414.000 2395.450 ;
        RECT 393.365 2395.135 393.695 2395.150 ;
        RECT 410.000 2395.000 414.000 2395.150 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 16.900 740.530 16.960 ;
        RECT 744.810 16.900 745.130 16.960 ;
        RECT 740.210 16.760 745.130 16.900 ;
        RECT 740.210 16.700 740.530 16.760 ;
        RECT 744.810 16.700 745.130 16.760 ;
      LAYER via ;
        RECT 740.240 16.700 740.500 16.960 ;
        RECT 744.840 16.700 745.100 16.960 ;
      LAYER met2 ;
        RECT 744.830 182.395 745.110 182.765 ;
        RECT 744.900 16.990 745.040 182.395 ;
        RECT 740.240 16.670 740.500 16.990 ;
        RECT 744.840 16.670 745.100 16.990 ;
        RECT 740.300 2.400 740.440 16.670 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 744.830 182.440 745.110 182.720 ;
      LAYER met3 ;
        RECT 2506.000 2895.930 2510.000 2896.080 ;
        RECT 2527.510 2895.930 2527.890 2895.940 ;
        RECT 2506.000 2895.630 2527.890 2895.930 ;
        RECT 2506.000 2895.480 2510.000 2895.630 ;
        RECT 2527.510 2895.620 2527.890 2895.630 ;
        RECT 744.805 182.730 745.135 182.745 ;
        RECT 2527.510 182.730 2527.890 182.740 ;
        RECT 744.805 182.430 2527.890 182.730 ;
        RECT 744.805 182.415 745.135 182.430 ;
        RECT 2527.510 182.420 2527.890 182.430 ;
      LAYER via3 ;
        RECT 2527.540 2895.620 2527.860 2895.940 ;
        RECT 2527.540 182.420 2527.860 182.740 ;
      LAYER met4 ;
        RECT 2527.535 2895.615 2527.865 2895.945 ;
        RECT 2527.550 182.745 2527.850 2895.615 ;
        RECT 2527.535 182.415 2527.865 182.745 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1716.330 3016.380 1716.650 3016.440 ;
        RECT 2560.430 3016.380 2560.750 3016.440 ;
        RECT 1716.330 3016.240 2560.750 3016.380 ;
        RECT 1716.330 3016.180 1716.650 3016.240 ;
        RECT 2560.430 3016.180 2560.750 3016.240 ;
        RECT 1881.930 45.120 1882.250 45.180 ;
        RECT 2560.430 45.120 2560.750 45.180 ;
        RECT 1881.930 44.980 2560.750 45.120 ;
        RECT 1881.930 44.920 1882.250 44.980 ;
        RECT 2560.430 44.920 2560.750 44.980 ;
      LAYER via ;
        RECT 1716.360 3016.180 1716.620 3016.440 ;
        RECT 2560.460 3016.180 2560.720 3016.440 ;
        RECT 1881.960 44.920 1882.220 45.180 ;
        RECT 2560.460 44.920 2560.720 45.180 ;
      LAYER met2 ;
        RECT 1716.360 3016.150 1716.620 3016.470 ;
        RECT 2560.460 3016.150 2560.720 3016.470 ;
        RECT 1716.420 3010.000 1716.560 3016.150 ;
        RECT 1716.420 3009.340 1716.770 3010.000 ;
        RECT 1716.490 3006.000 1716.770 3009.340 ;
        RECT 2560.520 45.210 2560.660 3016.150 ;
        RECT 1881.960 44.890 1882.220 45.210 ;
        RECT 2560.460 44.890 2560.720 45.210 ;
        RECT 1882.020 2.400 1882.160 44.890 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 286.180 1904.330 286.240 ;
        RECT 2159.770 286.180 2160.090 286.240 ;
        RECT 1904.010 286.040 2160.090 286.180 ;
        RECT 1904.010 285.980 1904.330 286.040 ;
        RECT 2159.770 285.980 2160.090 286.040 ;
        RECT 1899.870 16.900 1900.190 16.960 ;
        RECT 1904.010 16.900 1904.330 16.960 ;
        RECT 1899.870 16.760 1904.330 16.900 ;
        RECT 1899.870 16.700 1900.190 16.760 ;
        RECT 1904.010 16.700 1904.330 16.760 ;
      LAYER via ;
        RECT 1904.040 285.980 1904.300 286.240 ;
        RECT 2159.800 285.980 2160.060 286.240 ;
        RECT 1899.900 16.700 1900.160 16.960 ;
        RECT 1904.040 16.700 1904.300 16.960 ;
      LAYER met2 ;
        RECT 2166.370 510.410 2166.650 514.000 ;
        RECT 2159.860 510.270 2166.650 510.410 ;
        RECT 2159.860 286.270 2160.000 510.270 ;
        RECT 2166.370 510.000 2166.650 510.270 ;
        RECT 1904.040 285.950 1904.300 286.270 ;
        RECT 2159.800 285.950 2160.060 286.270 ;
        RECT 1904.100 16.990 1904.240 285.950 ;
        RECT 1899.900 16.670 1900.160 16.990 ;
        RECT 1904.040 16.670 1904.300 16.990 ;
        RECT 1899.960 2.400 1900.100 16.670 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 404.410 258.640 404.730 258.700 ;
        RECT 1911.370 258.640 1911.690 258.700 ;
        RECT 404.410 258.500 1911.690 258.640 ;
        RECT 404.410 258.440 404.730 258.500 ;
        RECT 1911.370 258.440 1911.690 258.500 ;
        RECT 1911.370 16.900 1911.690 16.960 ;
        RECT 1917.810 16.900 1918.130 16.960 ;
        RECT 1911.370 16.760 1918.130 16.900 ;
        RECT 1911.370 16.700 1911.690 16.760 ;
        RECT 1917.810 16.700 1918.130 16.760 ;
      LAYER via ;
        RECT 404.440 258.440 404.700 258.700 ;
        RECT 1911.400 258.440 1911.660 258.700 ;
        RECT 1911.400 16.700 1911.660 16.960 ;
        RECT 1917.840 16.700 1918.100 16.960 ;
      LAYER met2 ;
        RECT 404.430 1700.155 404.710 1700.525 ;
        RECT 404.500 258.730 404.640 1700.155 ;
        RECT 404.440 258.410 404.700 258.730 ;
        RECT 1911.400 258.410 1911.660 258.730 ;
        RECT 1911.460 16.990 1911.600 258.410 ;
        RECT 1911.400 16.670 1911.660 16.990 ;
        RECT 1917.840 16.670 1918.100 16.990 ;
        RECT 1917.900 2.400 1918.040 16.670 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
      LAYER via2 ;
        RECT 404.430 1700.200 404.710 1700.480 ;
      LAYER met3 ;
        RECT 404.405 1700.490 404.735 1700.505 ;
        RECT 410.000 1700.490 414.000 1700.640 ;
        RECT 404.405 1700.190 414.000 1700.490 ;
        RECT 404.405 1700.175 404.735 1700.190 ;
        RECT 410.000 1700.040 414.000 1700.190 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 397.050 3018.420 397.370 3018.480 ;
        RECT 542.410 3018.420 542.730 3018.480 ;
        RECT 397.050 3018.280 542.730 3018.420 ;
        RECT 397.050 3018.220 397.370 3018.280 ;
        RECT 542.410 3018.220 542.730 3018.280 ;
      LAYER via ;
        RECT 397.080 3018.220 397.340 3018.480 ;
        RECT 542.440 3018.220 542.700 3018.480 ;
      LAYER met2 ;
        RECT 397.080 3018.190 397.340 3018.510 ;
        RECT 542.440 3018.190 542.700 3018.510 ;
        RECT 397.140 938.925 397.280 3018.190 ;
        RECT 542.500 3010.000 542.640 3018.190 ;
        RECT 542.500 3009.340 542.850 3010.000 ;
        RECT 542.570 3006.000 542.850 3009.340 ;
        RECT 397.070 938.555 397.350 938.925 ;
        RECT 1932.090 58.635 1932.370 59.005 ;
        RECT 1932.160 17.410 1932.300 58.635 ;
        RECT 1932.160 17.270 1935.520 17.410 ;
        RECT 1935.380 2.400 1935.520 17.270 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 397.070 938.600 397.350 938.880 ;
        RECT 1932.090 58.680 1932.370 58.960 ;
      LAYER met3 ;
        RECT 377.470 938.890 377.850 938.900 ;
        RECT 397.045 938.890 397.375 938.905 ;
        RECT 377.470 938.590 397.375 938.890 ;
        RECT 377.470 938.580 377.850 938.590 ;
        RECT 397.045 938.575 397.375 938.590 ;
        RECT 377.470 58.970 377.850 58.980 ;
        RECT 1932.065 58.970 1932.395 58.985 ;
        RECT 377.470 58.670 1932.395 58.970 ;
        RECT 377.470 58.660 377.850 58.670 ;
        RECT 1932.065 58.655 1932.395 58.670 ;
      LAYER via3 ;
        RECT 377.500 938.580 377.820 938.900 ;
        RECT 377.500 58.660 377.820 58.980 ;
      LAYER met4 ;
        RECT 377.495 938.575 377.825 938.905 ;
        RECT 377.510 58.985 377.810 938.575 ;
        RECT 377.495 58.655 377.825 58.985 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 396.590 3025.220 396.910 3025.280 ;
        RECT 801.850 3025.220 802.170 3025.280 ;
        RECT 396.590 3025.080 802.170 3025.220 ;
        RECT 396.590 3025.020 396.910 3025.080 ;
        RECT 801.850 3025.020 802.170 3025.080 ;
        RECT 368.990 631.280 369.310 631.340 ;
        RECT 396.590 631.280 396.910 631.340 ;
        RECT 368.990 631.140 396.910 631.280 ;
        RECT 368.990 631.080 369.310 631.140 ;
        RECT 396.590 631.080 396.910 631.140 ;
        RECT 365.310 545.260 365.630 545.320 ;
        RECT 368.990 545.260 369.310 545.320 ;
        RECT 365.310 545.120 369.310 545.260 ;
        RECT 365.310 545.060 365.630 545.120 ;
        RECT 368.990 545.060 369.310 545.120 ;
      LAYER via ;
        RECT 396.620 3025.020 396.880 3025.280 ;
        RECT 801.880 3025.020 802.140 3025.280 ;
        RECT 369.020 631.080 369.280 631.340 ;
        RECT 396.620 631.080 396.880 631.340 ;
        RECT 365.340 545.060 365.600 545.320 ;
        RECT 369.020 545.060 369.280 545.320 ;
      LAYER met2 ;
        RECT 396.620 3024.990 396.880 3025.310 ;
        RECT 801.880 3024.990 802.140 3025.310 ;
        RECT 396.680 631.370 396.820 3024.990 ;
        RECT 801.940 3010.000 802.080 3024.990 ;
        RECT 801.940 3009.340 802.290 3010.000 ;
        RECT 802.010 3006.000 802.290 3009.340 ;
        RECT 369.020 631.050 369.280 631.370 ;
        RECT 396.620 631.050 396.880 631.370 ;
        RECT 369.080 545.350 369.220 631.050 ;
        RECT 365.340 545.030 365.600 545.350 ;
        RECT 369.020 545.030 369.280 545.350 ;
        RECT 365.400 46.085 365.540 545.030 ;
        RECT 365.330 45.715 365.610 46.085 ;
        RECT 1953.250 45.715 1953.530 46.085 ;
        RECT 1953.320 2.400 1953.460 45.715 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER via2 ;
        RECT 365.330 45.760 365.610 46.040 ;
        RECT 1953.250 45.760 1953.530 46.040 ;
      LAYER met3 ;
        RECT 365.305 46.050 365.635 46.065 ;
        RECT 1953.225 46.050 1953.555 46.065 ;
        RECT 365.305 45.750 1953.555 46.050 ;
        RECT 365.305 45.735 365.635 45.750 ;
        RECT 1953.225 45.735 1953.555 45.750 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1254.950 251.840 1255.270 251.900 ;
        RECT 1966.570 251.840 1966.890 251.900 ;
        RECT 1254.950 251.700 1966.890 251.840 ;
        RECT 1254.950 251.640 1255.270 251.700 ;
        RECT 1966.570 251.640 1966.890 251.700 ;
        RECT 1966.570 2.960 1966.890 3.020 ;
        RECT 1971.170 2.960 1971.490 3.020 ;
        RECT 1966.570 2.820 1971.490 2.960 ;
        RECT 1966.570 2.760 1966.890 2.820 ;
        RECT 1971.170 2.760 1971.490 2.820 ;
      LAYER via ;
        RECT 1254.980 251.640 1255.240 251.900 ;
        RECT 1966.600 251.640 1966.860 251.900 ;
        RECT 1966.600 2.760 1966.860 3.020 ;
        RECT 1971.200 2.760 1971.460 3.020 ;
      LAYER met2 ;
        RECT 1252.810 510.410 1253.090 514.000 ;
        RECT 1252.810 510.270 1255.180 510.410 ;
        RECT 1252.810 510.000 1253.090 510.270 ;
        RECT 1255.040 251.930 1255.180 510.270 ;
        RECT 1254.980 251.610 1255.240 251.930 ;
        RECT 1966.600 251.610 1966.860 251.930 ;
        RECT 1966.660 3.050 1966.800 251.610 ;
        RECT 1966.600 2.730 1966.860 3.050 ;
        RECT 1971.200 2.730 1971.460 3.050 ;
        RECT 1971.260 2.400 1971.400 2.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 481.680 1994.030 481.740 ;
        RECT 2508.910 481.680 2509.230 481.740 ;
        RECT 1993.710 481.540 2509.230 481.680 ;
        RECT 1993.710 481.480 1994.030 481.540 ;
        RECT 2508.910 481.480 2509.230 481.540 ;
        RECT 1989.110 20.300 1989.430 20.360 ;
        RECT 1993.710 20.300 1994.030 20.360 ;
        RECT 1989.110 20.160 1994.030 20.300 ;
        RECT 1989.110 20.100 1989.430 20.160 ;
        RECT 1993.710 20.100 1994.030 20.160 ;
      LAYER via ;
        RECT 1993.740 481.480 1994.000 481.740 ;
        RECT 2508.940 481.480 2509.200 481.740 ;
        RECT 1989.140 20.100 1989.400 20.360 ;
        RECT 1993.740 20.100 1994.000 20.360 ;
      LAYER met2 ;
        RECT 2508.930 1395.515 2509.210 1395.885 ;
        RECT 2509.000 481.770 2509.140 1395.515 ;
        RECT 1993.740 481.450 1994.000 481.770 ;
        RECT 2508.940 481.450 2509.200 481.770 ;
        RECT 1993.800 20.390 1993.940 481.450 ;
        RECT 1989.140 20.070 1989.400 20.390 ;
        RECT 1993.740 20.070 1994.000 20.390 ;
        RECT 1989.200 2.400 1989.340 20.070 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 2508.930 1395.560 2509.210 1395.840 ;
      LAYER met3 ;
        RECT 2506.000 1398.120 2510.000 1398.720 ;
        RECT 2509.150 1395.865 2509.450 1398.120 ;
        RECT 2508.905 1395.550 2509.450 1395.865 ;
        RECT 2508.905 1395.535 2509.235 1395.550 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2518.570 828.140 2518.890 828.200 ;
        RECT 2561.810 828.140 2562.130 828.200 ;
        RECT 2518.570 828.000 2562.130 828.140 ;
        RECT 2518.570 827.940 2518.890 828.000 ;
        RECT 2561.810 827.940 2562.130 828.000 ;
        RECT 2006.590 18.940 2006.910 19.000 ;
        RECT 2561.810 18.940 2562.130 19.000 ;
        RECT 2006.590 18.800 2562.130 18.940 ;
        RECT 2006.590 18.740 2006.910 18.800 ;
        RECT 2561.810 18.740 2562.130 18.800 ;
      LAYER via ;
        RECT 2518.600 827.940 2518.860 828.200 ;
        RECT 2561.840 827.940 2562.100 828.200 ;
        RECT 2006.620 18.740 2006.880 19.000 ;
        RECT 2561.840 18.740 2562.100 19.000 ;
      LAYER met2 ;
        RECT 2518.590 832.475 2518.870 832.845 ;
        RECT 2518.660 828.230 2518.800 832.475 ;
        RECT 2518.600 827.910 2518.860 828.230 ;
        RECT 2561.840 827.910 2562.100 828.230 ;
        RECT 2561.900 19.030 2562.040 827.910 ;
        RECT 2006.620 18.710 2006.880 19.030 ;
        RECT 2561.840 18.710 2562.100 19.030 ;
        RECT 2006.680 2.400 2006.820 18.710 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 2518.590 832.520 2518.870 832.800 ;
      LAYER met3 ;
        RECT 2506.000 832.810 2510.000 832.960 ;
        RECT 2518.565 832.810 2518.895 832.825 ;
        RECT 2506.000 832.510 2518.895 832.810 ;
        RECT 2506.000 832.360 2510.000 832.510 ;
        RECT 2518.565 832.495 2518.895 832.510 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 408.090 245.380 408.410 245.440 ;
        RECT 2021.770 245.380 2022.090 245.440 ;
        RECT 408.090 245.240 2022.090 245.380 ;
        RECT 408.090 245.180 408.410 245.240 ;
        RECT 2021.770 245.180 2022.090 245.240 ;
        RECT 2021.770 62.120 2022.090 62.180 ;
        RECT 2024.530 62.120 2024.850 62.180 ;
        RECT 2021.770 61.980 2024.850 62.120 ;
        RECT 2021.770 61.920 2022.090 61.980 ;
        RECT 2024.530 61.920 2024.850 61.980 ;
      LAYER via ;
        RECT 408.120 245.180 408.380 245.440 ;
        RECT 2021.800 245.180 2022.060 245.440 ;
        RECT 2021.800 61.920 2022.060 62.180 ;
        RECT 2024.560 61.920 2024.820 62.180 ;
      LAYER met2 ;
        RECT 408.110 1353.355 408.390 1353.725 ;
        RECT 408.180 245.470 408.320 1353.355 ;
        RECT 408.120 245.150 408.380 245.470 ;
        RECT 2021.800 245.150 2022.060 245.470 ;
        RECT 2021.860 62.210 2022.000 245.150 ;
        RECT 2021.800 61.890 2022.060 62.210 ;
        RECT 2024.560 61.890 2024.820 62.210 ;
        RECT 2024.620 2.400 2024.760 61.890 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
      LAYER via2 ;
        RECT 408.110 1353.400 408.390 1353.680 ;
      LAYER met3 ;
        RECT 408.085 1353.690 408.415 1353.705 ;
        RECT 410.000 1353.690 414.000 1353.840 ;
        RECT 408.085 1353.390 414.000 1353.690 ;
        RECT 408.085 1353.375 408.415 1353.390 ;
        RECT 410.000 1353.240 414.000 1353.390 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 155.280 2049.230 155.340 ;
        RECT 2346.070 155.280 2346.390 155.340 ;
        RECT 2048.910 155.140 2346.390 155.280 ;
        RECT 2048.910 155.080 2049.230 155.140 ;
        RECT 2346.070 155.080 2346.390 155.140 ;
        RECT 2042.470 20.300 2042.790 20.360 ;
        RECT 2048.910 20.300 2049.230 20.360 ;
        RECT 2042.470 20.160 2049.230 20.300 ;
        RECT 2042.470 20.100 2042.790 20.160 ;
        RECT 2048.910 20.100 2049.230 20.160 ;
      LAYER via ;
        RECT 2048.940 155.080 2049.200 155.340 ;
        RECT 2346.100 155.080 2346.360 155.340 ;
        RECT 2042.500 20.100 2042.760 20.360 ;
        RECT 2048.940 20.100 2049.200 20.360 ;
      LAYER met2 ;
        RECT 2352.210 510.410 2352.490 514.000 ;
        RECT 2346.160 510.270 2352.490 510.410 ;
        RECT 2346.160 155.370 2346.300 510.270 ;
        RECT 2352.210 510.000 2352.490 510.270 ;
        RECT 2048.940 155.050 2049.200 155.370 ;
        RECT 2346.100 155.050 2346.360 155.370 ;
        RECT 2049.000 20.390 2049.140 155.050 ;
        RECT 2042.500 20.070 2042.760 20.390 ;
        RECT 2048.940 20.070 2049.200 20.390 ;
        RECT 2042.560 2.400 2042.700 20.070 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1994.340 2519.810 1994.400 ;
        RECT 2604.130 1994.340 2604.450 1994.400 ;
        RECT 2519.490 1994.200 2604.450 1994.340 ;
        RECT 2519.490 1994.140 2519.810 1994.200 ;
        RECT 2604.130 1994.140 2604.450 1994.200 ;
        RECT 758.610 479.640 758.930 479.700 ;
        RECT 2604.130 479.640 2604.450 479.700 ;
        RECT 758.610 479.500 2604.450 479.640 ;
        RECT 758.610 479.440 758.930 479.500 ;
        RECT 2604.130 479.440 2604.450 479.500 ;
      LAYER via ;
        RECT 2519.520 1994.140 2519.780 1994.400 ;
        RECT 2604.160 1994.140 2604.420 1994.400 ;
        RECT 758.640 479.440 758.900 479.700 ;
        RECT 2604.160 479.440 2604.420 479.700 ;
      LAYER met2 ;
        RECT 2519.510 2000.715 2519.790 2001.085 ;
        RECT 2519.580 1994.430 2519.720 2000.715 ;
        RECT 2519.520 1994.110 2519.780 1994.430 ;
        RECT 2604.160 1994.110 2604.420 1994.430 ;
        RECT 2604.220 479.730 2604.360 1994.110 ;
        RECT 758.640 479.410 758.900 479.730 ;
        RECT 2604.160 479.410 2604.420 479.730 ;
        RECT 758.700 17.410 758.840 479.410 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2000.760 2519.790 2001.040 ;
      LAYER met3 ;
        RECT 2506.000 2001.050 2510.000 2001.200 ;
        RECT 2519.485 2001.050 2519.815 2001.065 ;
        RECT 2506.000 2000.750 2519.815 2001.050 ;
        RECT 2506.000 2000.600 2510.000 2000.750 ;
        RECT 2519.485 2000.735 2519.815 2000.750 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 79.460 2063.030 79.520 ;
        RECT 2139.070 79.460 2139.390 79.520 ;
        RECT 2062.710 79.320 2139.390 79.460 ;
        RECT 2062.710 79.260 2063.030 79.320 ;
        RECT 2139.070 79.260 2139.390 79.320 ;
        RECT 2060.410 20.300 2060.730 20.360 ;
        RECT 2062.710 20.300 2063.030 20.360 ;
        RECT 2060.410 20.160 2063.030 20.300 ;
        RECT 2060.410 20.100 2060.730 20.160 ;
        RECT 2062.710 20.100 2063.030 20.160 ;
      LAYER via ;
        RECT 2062.740 79.260 2063.000 79.520 ;
        RECT 2139.100 79.260 2139.360 79.520 ;
        RECT 2060.440 20.100 2060.700 20.360 ;
        RECT 2062.740 20.100 2063.000 20.360 ;
      LAYER met2 ;
        RECT 2141.530 510.410 2141.810 514.000 ;
        RECT 2139.160 510.270 2141.810 510.410 ;
        RECT 2139.160 79.550 2139.300 510.270 ;
        RECT 2141.530 510.000 2141.810 510.270 ;
        RECT 2062.740 79.230 2063.000 79.550 ;
        RECT 2139.100 79.230 2139.360 79.550 ;
        RECT 2062.800 20.390 2062.940 79.230 ;
        RECT 2060.440 20.070 2060.700 20.390 ;
        RECT 2062.740 20.070 2063.000 20.390 ;
        RECT 2060.500 2.400 2060.640 20.070 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2083.485 513.145 2083.655 513.995 ;
      LAYER mcon ;
        RECT 2083.485 513.825 2083.655 513.995 ;
      LAYER met1 ;
        RECT 2516.270 552.400 2516.590 552.460 ;
        RECT 2546.170 552.400 2546.490 552.460 ;
        RECT 2516.270 552.260 2546.490 552.400 ;
        RECT 2516.270 552.200 2516.590 552.260 ;
        RECT 2546.170 552.200 2546.490 552.260 ;
        RECT 2546.170 514.320 2546.490 514.380 ;
        RECT 2083.500 514.180 2546.490 514.320 ;
        RECT 2083.500 514.025 2083.640 514.180 ;
        RECT 2546.170 514.120 2546.490 514.180 ;
        RECT 2083.425 513.795 2083.715 514.025 ;
        RECT 2083.410 513.300 2083.730 513.360 ;
        RECT 2083.410 513.160 2083.925 513.300 ;
        RECT 2083.410 513.100 2083.730 513.160 ;
        RECT 2078.350 15.540 2078.670 15.600 ;
        RECT 2083.410 15.540 2083.730 15.600 ;
        RECT 2078.350 15.400 2083.730 15.540 ;
        RECT 2078.350 15.340 2078.670 15.400 ;
        RECT 2083.410 15.340 2083.730 15.400 ;
      LAYER via ;
        RECT 2516.300 552.200 2516.560 552.460 ;
        RECT 2546.200 552.200 2546.460 552.460 ;
        RECT 2546.200 514.120 2546.460 514.380 ;
        RECT 2083.440 513.100 2083.700 513.360 ;
        RECT 2078.380 15.340 2078.640 15.600 ;
        RECT 2083.440 15.340 2083.700 15.600 ;
      LAYER met2 ;
        RECT 2516.290 557.755 2516.570 558.125 ;
        RECT 2516.360 552.490 2516.500 557.755 ;
        RECT 2516.300 552.170 2516.560 552.490 ;
        RECT 2546.200 552.170 2546.460 552.490 ;
        RECT 2546.260 514.410 2546.400 552.170 ;
        RECT 2546.200 514.090 2546.460 514.410 ;
        RECT 2083.440 513.070 2083.700 513.390 ;
        RECT 2083.500 15.630 2083.640 513.070 ;
        RECT 2078.380 15.310 2078.640 15.630 ;
        RECT 2083.440 15.310 2083.700 15.630 ;
        RECT 2078.440 2.400 2078.580 15.310 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
      LAYER via2 ;
        RECT 2516.290 557.800 2516.570 558.080 ;
      LAYER met3 ;
        RECT 2506.000 558.090 2510.000 558.240 ;
        RECT 2516.265 558.090 2516.595 558.105 ;
        RECT 2506.000 557.790 2516.595 558.090 ;
        RECT 2506.000 557.640 2510.000 557.790 ;
        RECT 2516.265 557.775 2516.595 557.790 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2746.420 2519.810 2746.480 ;
        RECT 2594.930 2746.420 2595.250 2746.480 ;
        RECT 2519.490 2746.280 2595.250 2746.420 ;
        RECT 2519.490 2746.220 2519.810 2746.280 ;
        RECT 2594.930 2746.220 2595.250 2746.280 ;
        RECT 2097.210 495.960 2097.530 496.020 ;
        RECT 2594.930 495.960 2595.250 496.020 ;
        RECT 2097.210 495.820 2595.250 495.960 ;
        RECT 2097.210 495.760 2097.530 495.820 ;
        RECT 2594.930 495.760 2595.250 495.820 ;
      LAYER via ;
        RECT 2519.520 2746.220 2519.780 2746.480 ;
        RECT 2594.960 2746.220 2595.220 2746.480 ;
        RECT 2097.240 495.760 2097.500 496.020 ;
        RECT 2594.960 495.760 2595.220 496.020 ;
      LAYER met2 ;
        RECT 2519.510 2750.075 2519.790 2750.445 ;
        RECT 2519.580 2746.510 2519.720 2750.075 ;
        RECT 2519.520 2746.190 2519.780 2746.510 ;
        RECT 2594.960 2746.190 2595.220 2746.510 ;
        RECT 2595.020 496.050 2595.160 2746.190 ;
        RECT 2097.240 495.730 2097.500 496.050 ;
        RECT 2594.960 495.730 2595.220 496.050 ;
        RECT 2097.300 17.410 2097.440 495.730 ;
        RECT 2095.920 17.270 2097.440 17.410 ;
        RECT 2095.920 2.400 2096.060 17.270 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2750.120 2519.790 2750.400 ;
      LAYER met3 ;
        RECT 2506.000 2750.410 2510.000 2750.560 ;
        RECT 2519.485 2750.410 2519.815 2750.425 ;
        RECT 2506.000 2750.110 2519.815 2750.410 ;
        RECT 2506.000 2749.960 2510.000 2750.110 ;
        RECT 2519.485 2750.095 2519.815 2750.110 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1372.325 3003.305 1372.495 3006.535 ;
      LAYER mcon ;
        RECT 1372.325 3006.365 1372.495 3006.535 ;
      LAYER met1 ;
        RECT 1372.250 3006.520 1372.570 3006.580 ;
        RECT 1372.055 3006.380 1372.570 3006.520 ;
        RECT 1372.250 3006.320 1372.570 3006.380 ;
        RECT 1372.265 3003.460 1372.555 3003.505 ;
        RECT 2581.130 3003.460 2581.450 3003.520 ;
        RECT 1372.265 3003.320 2581.450 3003.460 ;
        RECT 1372.265 3003.275 1372.555 3003.320 ;
        RECT 2581.130 3003.260 2581.450 3003.320 ;
        RECT 2113.770 32.200 2114.090 32.260 ;
        RECT 2581.130 32.200 2581.450 32.260 ;
        RECT 2113.770 32.060 2581.450 32.200 ;
        RECT 2113.770 32.000 2114.090 32.060 ;
        RECT 2581.130 32.000 2581.450 32.060 ;
      LAYER via ;
        RECT 1372.280 3006.320 1372.540 3006.580 ;
        RECT 2581.160 3003.260 2581.420 3003.520 ;
        RECT 2113.800 32.000 2114.060 32.260 ;
        RECT 2581.160 32.000 2581.420 32.260 ;
      LAYER met2 ;
        RECT 1370.570 3006.690 1370.850 3010.000 ;
        RECT 1370.570 3006.610 1372.480 3006.690 ;
        RECT 1370.570 3006.550 1372.540 3006.610 ;
        RECT 1370.570 3006.000 1370.850 3006.550 ;
        RECT 1372.280 3006.290 1372.540 3006.550 ;
        RECT 2581.160 3003.230 2581.420 3003.550 ;
        RECT 2581.220 32.290 2581.360 3003.230 ;
        RECT 2113.800 31.970 2114.060 32.290 ;
        RECT 2581.160 31.970 2581.420 32.290 ;
        RECT 2113.860 2.400 2114.000 31.970 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 511.130 499.360 511.450 499.420 ;
        RECT 517.110 499.360 517.430 499.420 ;
        RECT 511.130 499.220 517.430 499.360 ;
        RECT 511.130 499.160 511.450 499.220 ;
        RECT 517.110 499.160 517.430 499.220 ;
        RECT 517.110 224.640 517.430 224.700 ;
        RECT 2125.270 224.640 2125.590 224.700 ;
        RECT 517.110 224.500 2125.590 224.640 ;
        RECT 517.110 224.440 517.430 224.500 ;
        RECT 2125.270 224.440 2125.590 224.500 ;
        RECT 2125.270 16.900 2125.590 16.960 ;
        RECT 2131.710 16.900 2132.030 16.960 ;
        RECT 2125.270 16.760 2132.030 16.900 ;
        RECT 2125.270 16.700 2125.590 16.760 ;
        RECT 2131.710 16.700 2132.030 16.760 ;
      LAYER via ;
        RECT 511.160 499.160 511.420 499.420 ;
        RECT 517.140 499.160 517.400 499.420 ;
        RECT 517.140 224.440 517.400 224.700 ;
        RECT 2125.300 224.440 2125.560 224.700 ;
        RECT 2125.300 16.700 2125.560 16.960 ;
        RECT 2131.740 16.700 2132.000 16.960 ;
      LAYER met2 ;
        RECT 511.290 510.340 511.570 514.000 ;
        RECT 511.220 510.000 511.570 510.340 ;
        RECT 511.220 499.450 511.360 510.000 ;
        RECT 511.160 499.130 511.420 499.450 ;
        RECT 517.140 499.130 517.400 499.450 ;
        RECT 517.200 224.730 517.340 499.130 ;
        RECT 517.140 224.410 517.400 224.730 ;
        RECT 2125.300 224.410 2125.560 224.730 ;
        RECT 2125.360 16.990 2125.500 224.410 ;
        RECT 2125.300 16.670 2125.560 16.990 ;
        RECT 2131.740 16.670 2132.000 16.990 ;
        RECT 2131.800 2.400 2131.940 16.670 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1672.170 496.980 1672.490 497.040 ;
        RECT 1676.310 496.980 1676.630 497.040 ;
        RECT 1672.170 496.840 1676.630 496.980 ;
        RECT 1672.170 496.780 1672.490 496.840 ;
        RECT 1676.310 496.780 1676.630 496.840 ;
        RECT 1676.310 231.440 1676.630 231.500 ;
        RECT 2145.970 231.440 2146.290 231.500 ;
        RECT 1676.310 231.300 2146.290 231.440 ;
        RECT 1676.310 231.240 1676.630 231.300 ;
        RECT 2145.970 231.240 2146.290 231.300 ;
      LAYER via ;
        RECT 1672.200 496.780 1672.460 497.040 ;
        RECT 1676.340 496.780 1676.600 497.040 ;
        RECT 1676.340 231.240 1676.600 231.500 ;
        RECT 2146.000 231.240 2146.260 231.500 ;
      LAYER met2 ;
        RECT 1672.330 510.340 1672.610 514.000 ;
        RECT 1672.260 510.000 1672.610 510.340 ;
        RECT 1672.260 497.070 1672.400 510.000 ;
        RECT 1672.200 496.750 1672.460 497.070 ;
        RECT 1676.340 496.750 1676.600 497.070 ;
        RECT 1676.400 231.530 1676.540 496.750 ;
        RECT 1676.340 231.210 1676.600 231.530 ;
        RECT 2146.000 231.210 2146.260 231.530 ;
        RECT 2146.060 16.730 2146.200 231.210 ;
        RECT 2146.060 16.590 2149.880 16.730 ;
        RECT 2149.740 2.400 2149.880 16.590 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.150 237.475 2167.430 237.845 ;
        RECT 2167.220 17.410 2167.360 237.475 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 2167.150 237.520 2167.430 237.800 ;
      LAYER met3 ;
        RECT 405.990 2668.810 406.370 2668.820 ;
        RECT 410.000 2668.810 414.000 2668.960 ;
        RECT 405.990 2668.510 414.000 2668.810 ;
        RECT 405.990 2668.500 406.370 2668.510 ;
        RECT 410.000 2668.360 414.000 2668.510 ;
        RECT 405.990 237.810 406.370 237.820 ;
        RECT 2167.125 237.810 2167.455 237.825 ;
        RECT 405.990 237.510 2167.455 237.810 ;
        RECT 405.990 237.500 406.370 237.510 ;
        RECT 2167.125 237.495 2167.455 237.510 ;
      LAYER via3 ;
        RECT 406.020 2668.500 406.340 2668.820 ;
        RECT 406.020 237.500 406.340 237.820 ;
      LAYER met4 ;
        RECT 406.015 2668.495 406.345 2668.825 ;
        RECT 406.030 237.825 406.330 2668.495 ;
        RECT 406.015 237.495 406.345 237.825 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 398.965 379.525 399.135 427.635 ;
        RECT 399.425 254.405 399.595 289.595 ;
      LAYER mcon ;
        RECT 398.965 427.465 399.135 427.635 ;
        RECT 399.425 289.425 399.595 289.595 ;
      LAYER met1 ;
        RECT 397.510 1052.200 397.830 1052.260 ;
        RECT 398.430 1052.200 398.750 1052.260 ;
        RECT 397.510 1052.060 398.750 1052.200 ;
        RECT 397.510 1052.000 397.830 1052.060 ;
        RECT 398.430 1052.000 398.750 1052.060 ;
        RECT 397.510 997.800 397.830 997.860 ;
        RECT 398.430 997.800 398.750 997.860 ;
        RECT 397.510 997.660 398.750 997.800 ;
        RECT 397.510 997.600 397.830 997.660 ;
        RECT 398.430 997.600 398.750 997.660 ;
        RECT 397.510 952.580 397.830 952.640 ;
        RECT 398.430 952.580 398.750 952.640 ;
        RECT 397.510 952.440 398.750 952.580 ;
        RECT 397.510 952.380 397.830 952.440 ;
        RECT 398.430 952.380 398.750 952.440 ;
        RECT 397.510 903.960 397.830 904.020 ;
        RECT 398.430 903.960 398.750 904.020 ;
        RECT 397.510 903.820 398.750 903.960 ;
        RECT 397.510 903.760 397.830 903.820 ;
        RECT 398.430 903.760 398.750 903.820 ;
        RECT 397.510 855.680 397.830 855.740 ;
        RECT 398.430 855.680 398.750 855.740 ;
        RECT 397.510 855.540 398.750 855.680 ;
        RECT 397.510 855.480 397.830 855.540 ;
        RECT 398.430 855.480 398.750 855.540 ;
        RECT 397.510 831.540 397.830 831.600 ;
        RECT 398.430 831.540 398.750 831.600 ;
        RECT 397.510 831.400 398.750 831.540 ;
        RECT 397.510 831.340 397.830 831.400 ;
        RECT 398.430 831.340 398.750 831.400 ;
        RECT 397.510 759.120 397.830 759.180 ;
        RECT 398.430 759.120 398.750 759.180 ;
        RECT 397.510 758.980 398.750 759.120 ;
        RECT 397.510 758.920 397.830 758.980 ;
        RECT 398.430 758.920 398.750 758.980 ;
        RECT 398.430 710.500 398.750 710.560 ;
        RECT 399.810 710.500 400.130 710.560 ;
        RECT 398.430 710.360 400.130 710.500 ;
        RECT 398.430 710.300 398.750 710.360 ;
        RECT 399.810 710.300 400.130 710.360 ;
        RECT 398.430 662.560 398.750 662.620 ;
        RECT 399.810 662.560 400.130 662.620 ;
        RECT 398.430 662.420 400.130 662.560 ;
        RECT 398.430 662.360 398.750 662.420 ;
        RECT 399.810 662.360 400.130 662.420 ;
        RECT 398.430 613.940 398.750 614.000 ;
        RECT 399.810 613.940 400.130 614.000 ;
        RECT 398.430 613.800 400.130 613.940 ;
        RECT 398.430 613.740 398.750 613.800 ;
        RECT 399.810 613.740 400.130 613.800 ;
        RECT 398.430 566.000 398.750 566.060 ;
        RECT 399.810 566.000 400.130 566.060 ;
        RECT 398.430 565.860 400.130 566.000 ;
        RECT 398.430 565.800 398.750 565.860 ;
        RECT 399.810 565.800 400.130 565.860 ;
        RECT 398.430 511.260 398.750 511.320 ;
        RECT 399.350 511.260 399.670 511.320 ;
        RECT 398.430 511.120 399.670 511.260 ;
        RECT 398.430 511.060 398.750 511.120 ;
        RECT 399.350 511.060 399.670 511.120 ;
        RECT 398.890 427.620 399.210 427.680 ;
        RECT 398.695 427.480 399.210 427.620 ;
        RECT 398.890 427.420 399.210 427.480 ;
        RECT 398.905 379.680 399.195 379.725 ;
        RECT 399.810 379.680 400.130 379.740 ;
        RECT 398.905 379.540 400.130 379.680 ;
        RECT 398.905 379.495 399.195 379.540 ;
        RECT 399.810 379.480 400.130 379.540 ;
        RECT 398.890 338.200 399.210 338.260 ;
        RECT 399.810 338.200 400.130 338.260 ;
        RECT 398.890 338.060 400.130 338.200 ;
        RECT 398.890 338.000 399.210 338.060 ;
        RECT 399.810 338.000 400.130 338.060 ;
        RECT 398.430 303.520 398.750 303.580 ;
        RECT 399.350 303.520 399.670 303.580 ;
        RECT 398.430 303.380 399.670 303.520 ;
        RECT 398.430 303.320 398.750 303.380 ;
        RECT 399.350 303.320 399.670 303.380 ;
        RECT 399.350 289.580 399.670 289.640 ;
        RECT 399.155 289.440 399.670 289.580 ;
        RECT 399.350 289.380 399.670 289.440 ;
        RECT 399.350 254.560 399.670 254.620 ;
        RECT 399.155 254.420 399.670 254.560 ;
        RECT 399.350 254.360 399.670 254.420 ;
        RECT 399.350 189.620 399.670 189.680 ;
        RECT 2180.470 189.620 2180.790 189.680 ;
        RECT 399.350 189.480 2180.790 189.620 ;
        RECT 399.350 189.420 399.670 189.480 ;
        RECT 2180.470 189.420 2180.790 189.480 ;
      LAYER via ;
        RECT 397.540 1052.000 397.800 1052.260 ;
        RECT 398.460 1052.000 398.720 1052.260 ;
        RECT 397.540 997.600 397.800 997.860 ;
        RECT 398.460 997.600 398.720 997.860 ;
        RECT 397.540 952.380 397.800 952.640 ;
        RECT 398.460 952.380 398.720 952.640 ;
        RECT 397.540 903.760 397.800 904.020 ;
        RECT 398.460 903.760 398.720 904.020 ;
        RECT 397.540 855.480 397.800 855.740 ;
        RECT 398.460 855.480 398.720 855.740 ;
        RECT 397.540 831.340 397.800 831.600 ;
        RECT 398.460 831.340 398.720 831.600 ;
        RECT 397.540 758.920 397.800 759.180 ;
        RECT 398.460 758.920 398.720 759.180 ;
        RECT 398.460 710.300 398.720 710.560 ;
        RECT 399.840 710.300 400.100 710.560 ;
        RECT 398.460 662.360 398.720 662.620 ;
        RECT 399.840 662.360 400.100 662.620 ;
        RECT 398.460 613.740 398.720 614.000 ;
        RECT 399.840 613.740 400.100 614.000 ;
        RECT 398.460 565.800 398.720 566.060 ;
        RECT 399.840 565.800 400.100 566.060 ;
        RECT 398.460 511.060 398.720 511.320 ;
        RECT 399.380 511.060 399.640 511.320 ;
        RECT 398.920 427.420 399.180 427.680 ;
        RECT 399.840 379.480 400.100 379.740 ;
        RECT 398.920 338.000 399.180 338.260 ;
        RECT 399.840 338.000 400.100 338.260 ;
        RECT 398.460 303.320 398.720 303.580 ;
        RECT 399.380 303.320 399.640 303.580 ;
        RECT 399.380 289.380 399.640 289.640 ;
        RECT 399.380 254.360 399.640 254.620 ;
        RECT 399.380 189.420 399.640 189.680 ;
        RECT 2180.500 189.420 2180.760 189.680 ;
      LAYER met2 ;
        RECT 398.450 1298.955 398.730 1299.325 ;
        RECT 398.520 1221.010 398.660 1298.955 ;
        RECT 398.060 1220.870 398.660 1221.010 ;
        RECT 398.060 1125.130 398.200 1220.870 ;
        RECT 397.600 1124.990 398.200 1125.130 ;
        RECT 397.600 1052.290 397.740 1124.990 ;
        RECT 397.540 1051.970 397.800 1052.290 ;
        RECT 398.460 1051.970 398.720 1052.290 ;
        RECT 398.520 997.890 398.660 1051.970 ;
        RECT 397.540 997.570 397.800 997.890 ;
        RECT 398.460 997.570 398.720 997.890 ;
        RECT 397.600 952.670 397.740 997.570 ;
        RECT 397.540 952.350 397.800 952.670 ;
        RECT 398.460 952.350 398.720 952.670 ;
        RECT 398.520 904.050 398.660 952.350 ;
        RECT 397.540 903.730 397.800 904.050 ;
        RECT 398.460 903.730 398.720 904.050 ;
        RECT 397.600 855.770 397.740 903.730 ;
        RECT 397.540 855.450 397.800 855.770 ;
        RECT 398.460 855.450 398.720 855.770 ;
        RECT 398.520 831.630 398.660 855.450 ;
        RECT 397.540 831.310 397.800 831.630 ;
        RECT 398.460 831.310 398.720 831.630 ;
        RECT 397.600 759.210 397.740 831.310 ;
        RECT 397.540 758.890 397.800 759.210 ;
        RECT 398.460 758.890 398.720 759.210 ;
        RECT 398.520 710.590 398.660 758.890 ;
        RECT 398.460 710.270 398.720 710.590 ;
        RECT 399.840 710.270 400.100 710.590 ;
        RECT 399.900 662.650 400.040 710.270 ;
        RECT 398.460 662.330 398.720 662.650 ;
        RECT 399.840 662.330 400.100 662.650 ;
        RECT 398.520 614.030 398.660 662.330 ;
        RECT 398.460 613.710 398.720 614.030 ;
        RECT 399.840 613.710 400.100 614.030 ;
        RECT 399.900 566.090 400.040 613.710 ;
        RECT 398.460 565.770 398.720 566.090 ;
        RECT 399.840 565.770 400.100 566.090 ;
        RECT 398.520 511.350 398.660 565.770 ;
        RECT 398.460 511.030 398.720 511.350 ;
        RECT 399.380 511.030 399.640 511.350 ;
        RECT 399.440 434.930 399.580 511.030 ;
        RECT 398.980 434.790 399.580 434.930 ;
        RECT 398.980 427.710 399.120 434.790 ;
        RECT 398.920 427.390 399.180 427.710 ;
        RECT 399.840 379.450 400.100 379.770 ;
        RECT 399.900 338.290 400.040 379.450 ;
        RECT 398.920 337.970 399.180 338.290 ;
        RECT 399.840 337.970 400.100 338.290 ;
        RECT 398.980 303.690 399.120 337.970 ;
        RECT 398.520 303.610 399.120 303.690 ;
        RECT 398.460 303.550 399.120 303.610 ;
        RECT 398.460 303.290 398.720 303.550 ;
        RECT 399.380 303.290 399.640 303.610 ;
        RECT 399.440 289.670 399.580 303.290 ;
        RECT 399.380 289.350 399.640 289.670 ;
        RECT 399.380 254.330 399.640 254.650 ;
        RECT 399.440 189.710 399.580 254.330 ;
        RECT 399.380 189.390 399.640 189.710 ;
        RECT 2180.500 189.390 2180.760 189.710 ;
        RECT 2180.560 16.730 2180.700 189.390 ;
        RECT 2180.560 16.590 2185.300 16.730 ;
        RECT 2185.160 2.400 2185.300 16.590 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
      LAYER via2 ;
        RECT 398.450 1299.000 398.730 1299.280 ;
      LAYER met3 ;
        RECT 398.425 1299.290 398.755 1299.305 ;
        RECT 410.000 1299.290 414.000 1299.440 ;
        RECT 398.425 1298.990 414.000 1299.290 ;
        RECT 398.425 1298.975 398.755 1298.990 ;
        RECT 410.000 1298.840 414.000 1298.990 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 142.020 2118.230 142.080 ;
        RECT 2201.170 142.020 2201.490 142.080 ;
        RECT 2117.910 141.880 2201.490 142.020 ;
        RECT 2117.910 141.820 2118.230 141.880 ;
        RECT 2201.170 141.820 2201.490 141.880 ;
      LAYER via ;
        RECT 2117.940 141.820 2118.200 142.080 ;
        RECT 2201.200 141.820 2201.460 142.080 ;
      LAYER met2 ;
        RECT 2117.610 510.410 2117.890 514.000 ;
        RECT 2117.080 510.270 2117.890 510.410 ;
        RECT 2117.080 483.325 2117.220 510.270 ;
        RECT 2117.610 510.000 2117.890 510.270 ;
        RECT 2117.010 482.955 2117.290 483.325 ;
        RECT 2117.930 482.955 2118.210 483.325 ;
        RECT 2118.000 142.110 2118.140 482.955 ;
        RECT 2117.940 141.790 2118.200 142.110 ;
        RECT 2201.200 141.790 2201.460 142.110 ;
        RECT 2201.260 16.730 2201.400 141.790 ;
        RECT 2201.260 16.590 2203.240 16.730 ;
        RECT 2203.100 2.400 2203.240 16.590 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
      LAYER via2 ;
        RECT 2117.010 483.000 2117.290 483.280 ;
        RECT 2117.930 483.000 2118.210 483.280 ;
      LAYER met3 ;
        RECT 2116.985 483.290 2117.315 483.305 ;
        RECT 2117.905 483.290 2118.235 483.305 ;
        RECT 2116.985 482.990 2118.235 483.290 ;
        RECT 2116.985 482.975 2117.315 482.990 ;
        RECT 2117.905 482.975 2118.235 482.990 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 915.085 3001.945 915.255 3006.535 ;
      LAYER mcon ;
        RECT 915.085 3006.365 915.255 3006.535 ;
      LAYER met1 ;
        RECT 915.010 3006.520 915.330 3006.580 ;
        RECT 914.815 3006.380 915.330 3006.520 ;
        RECT 915.010 3006.320 915.330 3006.380 ;
        RECT 915.025 3002.100 915.315 3002.145 ;
        RECT 2594.470 3002.100 2594.790 3002.160 ;
        RECT 915.025 3001.960 2594.790 3002.100 ;
        RECT 915.025 3001.915 915.315 3001.960 ;
        RECT 2594.470 3001.900 2594.790 3001.960 ;
        RECT 2220.950 45.460 2221.270 45.520 ;
        RECT 2594.470 45.460 2594.790 45.520 ;
        RECT 2220.950 45.320 2594.790 45.460 ;
        RECT 2220.950 45.260 2221.270 45.320 ;
        RECT 2594.470 45.260 2594.790 45.320 ;
      LAYER via ;
        RECT 915.040 3006.320 915.300 3006.580 ;
        RECT 2594.500 3001.900 2594.760 3002.160 ;
        RECT 2220.980 45.260 2221.240 45.520 ;
        RECT 2594.500 45.260 2594.760 45.520 ;
      LAYER met2 ;
        RECT 913.330 3006.690 913.610 3010.000 ;
        RECT 913.330 3006.610 915.240 3006.690 ;
        RECT 913.330 3006.550 915.300 3006.610 ;
        RECT 913.330 3006.000 913.610 3006.550 ;
        RECT 915.040 3006.290 915.300 3006.550 ;
        RECT 2594.500 3001.870 2594.760 3002.190 ;
        RECT 2594.560 45.550 2594.700 3001.870 ;
        RECT 2220.980 45.230 2221.240 45.550 ;
        RECT 2594.500 45.230 2594.760 45.550 ;
        RECT 2221.040 2.400 2221.180 45.230 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 231.100 779.630 231.160 ;
        RECT 2463.370 231.100 2463.690 231.160 ;
        RECT 779.310 230.960 2463.690 231.100 ;
        RECT 779.310 230.900 779.630 230.960 ;
        RECT 2463.370 230.900 2463.690 230.960 ;
        RECT 775.630 16.560 775.950 16.620 ;
        RECT 779.310 16.560 779.630 16.620 ;
        RECT 775.630 16.420 779.630 16.560 ;
        RECT 775.630 16.360 775.950 16.420 ;
        RECT 779.310 16.360 779.630 16.420 ;
      LAYER via ;
        RECT 779.340 230.900 779.600 231.160 ;
        RECT 2463.400 230.900 2463.660 231.160 ;
        RECT 775.660 16.360 775.920 16.620 ;
        RECT 779.340 16.360 779.600 16.620 ;
      LAYER met2 ;
        RECT 2463.530 510.340 2463.810 514.000 ;
        RECT 2463.460 510.000 2463.810 510.340 ;
        RECT 2463.460 231.190 2463.600 510.000 ;
        RECT 779.340 230.870 779.600 231.190 ;
        RECT 2463.400 230.870 2463.660 231.190 ;
        RECT 779.400 16.650 779.540 230.870 ;
        RECT 775.660 16.330 775.920 16.650 ;
        RECT 779.340 16.330 779.600 16.650 ;
        RECT 775.720 2.400 775.860 16.330 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 3009.580 1186.730 3009.640 ;
        RECT 2573.770 3009.580 2574.090 3009.640 ;
        RECT 1186.410 3009.440 2574.090 3009.580 ;
        RECT 1186.410 3009.380 1186.730 3009.440 ;
        RECT 2573.770 3009.380 2574.090 3009.440 ;
        RECT 2238.890 32.880 2239.210 32.940 ;
        RECT 2573.770 32.880 2574.090 32.940 ;
        RECT 2238.890 32.740 2574.090 32.880 ;
        RECT 2238.890 32.680 2239.210 32.740 ;
        RECT 2573.770 32.680 2574.090 32.740 ;
      LAYER via ;
        RECT 1186.440 3009.380 1186.700 3009.640 ;
        RECT 2573.800 3009.380 2574.060 3009.640 ;
        RECT 2238.920 32.680 2239.180 32.940 ;
        RECT 2573.800 32.680 2574.060 32.940 ;
      LAYER met2 ;
        RECT 1185.650 3009.410 1185.930 3010.000 ;
        RECT 1186.440 3009.410 1186.700 3009.670 ;
        RECT 1185.650 3009.350 1186.700 3009.410 ;
        RECT 2573.800 3009.350 2574.060 3009.670 ;
        RECT 1185.650 3009.270 1186.640 3009.350 ;
        RECT 1185.650 3006.000 1185.930 3009.270 ;
        RECT 2573.860 32.970 2574.000 3009.350 ;
        RECT 2238.920 32.650 2239.180 32.970 ;
        RECT 2573.800 32.650 2574.060 32.970 ;
        RECT 2238.980 2.400 2239.120 32.650 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2210.390 3016.635 2210.670 3017.005 ;
        RECT 2210.460 3010.000 2210.600 3016.635 ;
        RECT 2210.460 3009.340 2210.810 3010.000 ;
        RECT 2210.530 3006.000 2210.810 3009.340 ;
        RECT 2256.850 18.515 2257.130 18.885 ;
        RECT 2256.920 9.250 2257.060 18.515 ;
        RECT 2256.460 9.110 2257.060 9.250 ;
        RECT 2256.460 2.400 2256.600 9.110 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
      LAYER via2 ;
        RECT 2210.390 3016.680 2210.670 3016.960 ;
        RECT 2256.850 18.560 2257.130 18.840 ;
      LAYER met3 ;
        RECT 2210.365 3016.970 2210.695 3016.985 ;
        RECT 2429.990 3016.970 2430.370 3016.980 ;
        RECT 2210.365 3016.670 2430.370 3016.970 ;
        RECT 2210.365 3016.655 2210.695 3016.670 ;
        RECT 2429.990 3016.660 2430.370 3016.670 ;
        RECT 2256.825 18.850 2257.155 18.865 ;
        RECT 2429.990 18.850 2430.370 18.860 ;
        RECT 2256.825 18.550 2430.370 18.850 ;
        RECT 2256.825 18.535 2257.155 18.550 ;
        RECT 2429.990 18.540 2430.370 18.550 ;
      LAYER via3 ;
        RECT 2430.020 3016.660 2430.340 3016.980 ;
        RECT 2430.020 18.540 2430.340 18.860 ;
      LAYER met4 ;
        RECT 2430.015 3016.655 2430.345 3016.985 ;
        RECT 2430.030 18.865 2430.330 3016.655 ;
        RECT 2430.015 18.535 2430.345 18.865 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2270.170 62.120 2270.490 62.180 ;
        RECT 2274.310 62.120 2274.630 62.180 ;
        RECT 2270.170 61.980 2274.630 62.120 ;
        RECT 2270.170 61.920 2270.490 61.980 ;
        RECT 2274.310 61.920 2274.630 61.980 ;
      LAYER via ;
        RECT 2270.200 61.920 2270.460 62.180 ;
        RECT 2274.340 61.920 2274.600 62.180 ;
      LAYER met2 ;
        RECT 2270.190 452.355 2270.470 452.725 ;
        RECT 2270.260 62.210 2270.400 452.355 ;
        RECT 2270.200 61.890 2270.460 62.210 ;
        RECT 2274.340 61.890 2274.600 62.210 ;
        RECT 2274.400 2.400 2274.540 61.890 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
      LAYER via2 ;
        RECT 2270.190 452.400 2270.470 452.680 ;
      LAYER met3 ;
        RECT 396.790 1225.850 397.170 1225.860 ;
        RECT 410.000 1225.850 414.000 1226.000 ;
        RECT 396.790 1225.550 414.000 1225.850 ;
        RECT 396.790 1225.540 397.170 1225.550 ;
        RECT 410.000 1225.400 414.000 1225.550 ;
        RECT 396.790 452.690 397.170 452.700 ;
        RECT 2270.165 452.690 2270.495 452.705 ;
        RECT 396.790 452.390 2270.495 452.690 ;
        RECT 396.790 452.380 397.170 452.390 ;
        RECT 2270.165 452.375 2270.495 452.390 ;
      LAYER via3 ;
        RECT 396.820 1225.540 397.140 1225.860 ;
        RECT 396.820 452.380 397.140 452.700 ;
      LAYER met4 ;
        RECT 396.815 1225.535 397.145 1225.865 ;
        RECT 396.830 452.705 397.130 1225.535 ;
        RECT 396.815 452.375 397.145 452.705 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2290.890 299.355 2291.170 299.725 ;
        RECT 2290.960 16.730 2291.100 299.355 ;
        RECT 2290.960 16.590 2292.480 16.730 ;
        RECT 2292.340 2.400 2292.480 16.590 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
      LAYER via2 ;
        RECT 2290.890 299.400 2291.170 299.680 ;
      LAYER met3 ;
        RECT 408.750 1865.050 409.130 1865.060 ;
        RECT 410.000 1865.050 414.000 1865.200 ;
        RECT 408.750 1864.750 414.000 1865.050 ;
        RECT 408.750 1864.740 409.130 1864.750 ;
        RECT 410.000 1864.600 414.000 1864.750 ;
        RECT 408.750 299.690 409.130 299.700 ;
        RECT 2290.865 299.690 2291.195 299.705 ;
        RECT 408.750 299.390 2291.195 299.690 ;
        RECT 408.750 299.380 409.130 299.390 ;
        RECT 2290.865 299.375 2291.195 299.390 ;
      LAYER via3 ;
        RECT 408.780 1864.740 409.100 1865.060 ;
        RECT 408.780 299.380 409.100 299.700 ;
      LAYER met4 ;
        RECT 408.775 1864.735 409.105 1865.065 ;
        RECT 408.790 299.705 409.090 1864.735 ;
        RECT 408.775 299.375 409.105 299.705 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.570 502.420 1276.890 502.480 ;
        RECT 1283.010 502.420 1283.330 502.480 ;
        RECT 1276.570 502.280 1283.330 502.420 ;
        RECT 1276.570 502.220 1276.890 502.280 ;
        RECT 1283.010 502.220 1283.330 502.280 ;
        RECT 1283.010 162.080 1283.330 162.140 ;
        RECT 2304.670 162.080 2304.990 162.140 ;
        RECT 1283.010 161.940 2304.990 162.080 ;
        RECT 1283.010 161.880 1283.330 161.940 ;
        RECT 2304.670 161.880 2304.990 161.940 ;
      LAYER via ;
        RECT 1276.600 502.220 1276.860 502.480 ;
        RECT 1283.040 502.220 1283.300 502.480 ;
        RECT 1283.040 161.880 1283.300 162.140 ;
        RECT 2304.700 161.880 2304.960 162.140 ;
      LAYER met2 ;
        RECT 1276.730 510.340 1277.010 514.000 ;
        RECT 1276.660 510.000 1277.010 510.340 ;
        RECT 1276.660 502.510 1276.800 510.000 ;
        RECT 1276.600 502.190 1276.860 502.510 ;
        RECT 1283.040 502.190 1283.300 502.510 ;
        RECT 1283.100 162.170 1283.240 502.190 ;
        RECT 1283.040 161.850 1283.300 162.170 ;
        RECT 2304.700 161.850 2304.960 162.170 ;
        RECT 2304.760 17.410 2304.900 161.850 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.910 3023.435 790.190 3023.805 ;
        RECT 789.980 3010.000 790.120 3023.435 ;
        RECT 789.980 3009.340 790.330 3010.000 ;
        RECT 790.050 3006.000 790.330 3009.340 ;
        RECT 2481.790 227.275 2482.070 227.645 ;
        RECT 2481.860 203.845 2482.000 227.275 ;
        RECT 2481.790 203.475 2482.070 203.845 ;
        RECT 2328.150 13.755 2328.430 14.125 ;
        RECT 2328.220 2.400 2328.360 13.755 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
      LAYER via2 ;
        RECT 789.910 3023.480 790.190 3023.760 ;
        RECT 2481.790 227.320 2482.070 227.600 ;
        RECT 2481.790 203.520 2482.070 203.800 ;
        RECT 2328.150 13.800 2328.430 14.080 ;
      LAYER met3 ;
        RECT 789.885 3023.770 790.215 3023.785 ;
        RECT 2484.270 3023.770 2484.650 3023.780 ;
        RECT 789.885 3023.470 2484.650 3023.770 ;
        RECT 789.885 3023.455 790.215 3023.470 ;
        RECT 2484.270 3023.460 2484.650 3023.470 ;
        RECT 2484.270 3014.620 2484.650 3014.940 ;
        RECT 2484.310 3014.250 2484.610 3014.620 ;
        RECT 2486.110 3014.250 2486.490 3014.260 ;
        RECT 2484.310 3013.950 2486.490 3014.250 ;
        RECT 2486.110 3013.940 2486.490 3013.950 ;
        RECT 2482.430 469.380 2482.810 469.700 ;
        RECT 2482.470 468.340 2482.770 469.380 ;
        RECT 2482.430 468.020 2482.810 468.340 ;
        RECT 2482.430 428.210 2482.810 428.220 ;
        RECT 2481.550 427.910 2482.810 428.210 ;
        RECT 2481.550 426.850 2481.850 427.910 ;
        RECT 2482.430 427.900 2482.810 427.910 ;
        RECT 2482.430 426.850 2482.810 426.860 ;
        RECT 2481.550 426.550 2482.810 426.850 ;
        RECT 2482.430 426.540 2482.810 426.550 ;
        RECT 2481.765 227.610 2482.095 227.625 ;
        RECT 2482.430 227.610 2482.810 227.620 ;
        RECT 2481.765 227.310 2482.810 227.610 ;
        RECT 2481.765 227.295 2482.095 227.310 ;
        RECT 2482.430 227.300 2482.810 227.310 ;
        RECT 2481.765 203.820 2482.095 203.825 ;
        RECT 2481.510 203.810 2482.095 203.820 ;
        RECT 2481.310 203.510 2482.095 203.810 ;
        RECT 2481.510 203.500 2482.095 203.510 ;
        RECT 2481.765 203.495 2482.095 203.500 ;
        RECT 2481.510 63.050 2481.890 63.060 ;
        RECT 2480.630 62.750 2481.890 63.050 ;
        RECT 2480.630 61.700 2480.930 62.750 ;
        RECT 2481.510 62.740 2481.890 62.750 ;
        RECT 2480.590 61.380 2480.970 61.700 ;
        RECT 2328.125 14.090 2328.455 14.105 ;
        RECT 2330.630 14.090 2331.010 14.100 ;
        RECT 2328.125 13.790 2331.010 14.090 ;
        RECT 2328.125 13.775 2328.455 13.790 ;
        RECT 2330.630 13.780 2331.010 13.790 ;
      LAYER via3 ;
        RECT 2484.300 3023.460 2484.620 3023.780 ;
        RECT 2484.300 3014.620 2484.620 3014.940 ;
        RECT 2486.140 3013.940 2486.460 3014.260 ;
        RECT 2482.460 469.380 2482.780 469.700 ;
        RECT 2482.460 468.020 2482.780 468.340 ;
        RECT 2482.460 427.900 2482.780 428.220 ;
        RECT 2482.460 426.540 2482.780 426.860 ;
        RECT 2482.460 227.300 2482.780 227.620 ;
        RECT 2481.540 203.500 2481.860 203.820 ;
        RECT 2481.540 62.740 2481.860 63.060 ;
        RECT 2480.620 61.380 2480.940 61.700 ;
        RECT 2330.660 13.780 2330.980 14.100 ;
      LAYER met4 ;
        RECT 2484.295 3023.455 2484.625 3023.785 ;
        RECT 2484.310 3014.945 2484.610 3023.455 ;
        RECT 2484.295 3014.615 2484.625 3014.945 ;
        RECT 2486.135 3013.935 2486.465 3014.265 ;
        RECT 2486.150 2970.050 2486.450 3013.935 ;
        RECT 2484.310 2969.750 2486.450 2970.050 ;
        RECT 2484.310 2925.850 2484.610 2969.750 ;
        RECT 2484.310 2925.550 2485.530 2925.850 ;
        RECT 2485.230 2885.490 2485.530 2925.550 ;
        RECT 2484.790 2884.310 2485.970 2885.490 ;
        RECT 2493.070 2884.310 2494.250 2885.490 ;
        RECT 2493.510 2824.290 2493.810 2884.310 ;
        RECT 2483.870 2823.110 2485.050 2824.290 ;
        RECT 2493.070 2823.110 2494.250 2824.290 ;
        RECT 2484.310 2742.250 2484.610 2823.110 ;
        RECT 2483.390 2741.950 2484.610 2742.250 ;
        RECT 2483.390 2718.450 2483.690 2741.950 ;
        RECT 2483.390 2718.150 2485.530 2718.450 ;
        RECT 2485.230 2711.650 2485.530 2718.150 ;
        RECT 2483.390 2711.350 2485.530 2711.650 ;
        RECT 2483.390 2667.450 2483.690 2711.350 ;
        RECT 2483.390 2667.150 2485.530 2667.450 ;
        RECT 2485.230 2650.450 2485.530 2667.150 ;
        RECT 2483.390 2650.150 2485.530 2650.450 ;
        RECT 2483.390 2616.450 2483.690 2650.150 ;
        RECT 2483.390 2616.150 2485.530 2616.450 ;
        RECT 2485.230 2575.650 2485.530 2616.150 ;
        RECT 2484.310 2575.350 2485.530 2575.650 ;
        RECT 2484.310 2266.690 2484.610 2575.350 ;
        RECT 2483.870 2265.510 2485.050 2266.690 ;
        RECT 2489.390 2265.510 2490.570 2266.690 ;
        RECT 2489.830 2252.650 2490.130 2265.510 ;
        RECT 2488.910 2252.350 2490.130 2252.650 ;
        RECT 2488.910 2218.650 2489.210 2252.350 ;
        RECT 2488.910 2218.350 2490.130 2218.650 ;
        RECT 2489.830 2164.690 2490.130 2218.350 ;
        RECT 2484.790 2163.510 2485.970 2164.690 ;
        RECT 2489.390 2163.510 2490.570 2164.690 ;
        RECT 2485.230 2075.850 2485.530 2163.510 ;
        RECT 2484.310 2075.550 2485.530 2075.850 ;
        RECT 2484.310 2021.450 2484.610 2075.550 ;
        RECT 2480.630 2021.150 2484.610 2021.450 ;
        RECT 2480.630 2014.650 2480.930 2021.150 ;
        RECT 2480.630 2014.350 2481.850 2014.650 ;
        RECT 2481.550 1970.450 2481.850 2014.350 ;
        RECT 2481.550 1970.150 2483.690 1970.450 ;
        RECT 2483.390 1939.850 2483.690 1970.150 ;
        RECT 2483.390 1939.550 2485.530 1939.850 ;
        RECT 2485.230 1916.050 2485.530 1939.550 ;
        RECT 2484.310 1915.750 2485.530 1916.050 ;
        RECT 2484.310 1885.450 2484.610 1915.750 ;
        RECT 2484.310 1885.150 2485.530 1885.450 ;
        RECT 2485.230 1790.250 2485.530 1885.150 ;
        RECT 2485.230 1789.950 2488.290 1790.250 ;
        RECT 2487.990 1742.650 2488.290 1789.950 ;
        RECT 2485.230 1742.350 2488.290 1742.650 ;
        RECT 2485.230 1647.450 2485.530 1742.350 ;
        RECT 2484.310 1647.150 2485.530 1647.450 ;
        RECT 2484.310 1572.650 2484.610 1647.150 ;
        RECT 2484.310 1572.350 2485.530 1572.650 ;
        RECT 2485.230 1453.650 2485.530 1572.350 ;
        RECT 2484.310 1453.350 2485.530 1453.650 ;
        RECT 2484.310 1334.650 2484.610 1453.350 ;
        RECT 2483.390 1334.350 2484.610 1334.650 ;
        RECT 2483.390 1304.050 2483.690 1334.350 ;
        RECT 2482.470 1303.750 2483.690 1304.050 ;
        RECT 2482.470 1259.850 2482.770 1303.750 ;
        RECT 2480.630 1259.550 2482.770 1259.850 ;
        RECT 2480.630 1062.650 2480.930 1259.550 ;
        RECT 2480.630 1062.350 2481.850 1062.650 ;
        RECT 2481.550 1015.050 2481.850 1062.350 ;
        RECT 2480.630 1014.750 2481.850 1015.050 ;
        RECT 2480.630 938.890 2480.930 1014.750 ;
        RECT 2480.630 938.590 2483.690 938.890 ;
        RECT 2483.390 916.450 2483.690 938.590 ;
        RECT 2481.550 916.150 2483.690 916.450 ;
        RECT 2481.550 899.450 2481.850 916.150 ;
        RECT 2480.630 899.150 2481.850 899.450 ;
        RECT 2480.630 848.450 2480.930 899.150 ;
        RECT 2480.630 848.150 2481.850 848.450 ;
        RECT 2481.550 678.450 2481.850 848.150 ;
        RECT 2480.630 678.150 2481.850 678.450 ;
        RECT 2480.630 661.450 2480.930 678.150 ;
        RECT 2480.630 661.150 2481.850 661.450 ;
        RECT 2481.550 510.490 2481.850 661.150 ;
        RECT 2481.550 510.190 2482.770 510.490 ;
        RECT 2482.470 469.705 2482.770 510.190 ;
        RECT 2482.455 469.375 2482.785 469.705 ;
        RECT 2482.455 468.015 2482.785 468.345 ;
        RECT 2482.470 428.225 2482.770 468.015 ;
        RECT 2482.455 427.895 2482.785 428.225 ;
        RECT 2482.455 426.535 2482.785 426.865 ;
        RECT 2482.470 318.050 2482.770 426.535 ;
        RECT 2481.550 317.750 2482.770 318.050 ;
        RECT 2481.550 307.850 2481.850 317.750 ;
        RECT 2481.550 307.550 2482.770 307.850 ;
        RECT 2482.470 227.625 2482.770 307.550 ;
        RECT 2482.455 227.295 2482.785 227.625 ;
        RECT 2481.535 203.495 2481.865 203.825 ;
        RECT 2481.550 63.065 2481.850 203.495 ;
        RECT 2481.535 62.735 2481.865 63.065 ;
        RECT 2480.615 61.375 2480.945 61.705 ;
        RECT 2480.630 19.290 2480.930 61.375 ;
        RECT 2330.230 18.110 2331.410 19.290 ;
        RECT 2480.190 18.110 2481.370 19.290 ;
        RECT 2330.670 14.105 2330.970 18.110 ;
        RECT 2330.655 13.775 2330.985 14.105 ;
      LAYER met5 ;
        RECT 2484.580 2884.100 2494.460 2885.700 ;
        RECT 2483.660 2822.900 2494.460 2824.500 ;
        RECT 2483.660 2265.300 2490.780 2266.900 ;
        RECT 2484.580 2163.300 2490.780 2164.900 ;
        RECT 2330.020 17.900 2481.580 19.500 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 496.640 2345.930 496.700 ;
        RECT 2514.430 496.640 2514.750 496.700 ;
        RECT 2345.610 496.500 2514.750 496.640 ;
        RECT 2345.610 496.440 2345.930 496.500 ;
        RECT 2514.430 496.440 2514.750 496.500 ;
      LAYER via ;
        RECT 2345.640 496.440 2345.900 496.700 ;
        RECT 2514.460 496.440 2514.720 496.700 ;
      LAYER met2 ;
        RECT 2514.450 1088.155 2514.730 1088.525 ;
        RECT 2514.520 496.730 2514.660 1088.155 ;
        RECT 2345.640 496.410 2345.900 496.730 ;
        RECT 2514.460 496.410 2514.720 496.730 ;
        RECT 2345.700 2.400 2345.840 496.410 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 2514.450 1088.200 2514.730 1088.480 ;
      LAYER met3 ;
        RECT 2506.000 1088.490 2510.000 1088.640 ;
        RECT 2514.425 1088.490 2514.755 1088.505 ;
        RECT 2506.000 1088.190 2514.755 1088.490 ;
        RECT 2506.000 1088.040 2510.000 1088.190 ;
        RECT 2514.425 1088.175 2514.755 1088.190 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 308.270 2484.280 308.590 2484.340 ;
        RECT 393.370 2484.280 393.690 2484.340 ;
        RECT 308.270 2484.140 393.690 2484.280 ;
        RECT 308.270 2484.080 308.590 2484.140 ;
        RECT 393.370 2484.080 393.690 2484.140 ;
        RECT 308.270 60.080 308.590 60.140 ;
        RECT 2363.550 60.080 2363.870 60.140 ;
        RECT 308.270 59.940 2363.870 60.080 ;
        RECT 308.270 59.880 308.590 59.940 ;
        RECT 2363.550 59.880 2363.870 59.940 ;
      LAYER via ;
        RECT 308.300 2484.080 308.560 2484.340 ;
        RECT 393.400 2484.080 393.660 2484.340 ;
        RECT 308.300 59.880 308.560 60.140 ;
        RECT 2363.580 59.880 2363.840 60.140 ;
      LAYER met2 ;
        RECT 393.390 2486.235 393.670 2486.605 ;
        RECT 393.460 2484.370 393.600 2486.235 ;
        RECT 308.300 2484.050 308.560 2484.370 ;
        RECT 393.400 2484.050 393.660 2484.370 ;
        RECT 308.360 60.170 308.500 2484.050 ;
        RECT 308.300 59.850 308.560 60.170 ;
        RECT 2363.580 59.850 2363.840 60.170 ;
        RECT 2363.640 2.400 2363.780 59.850 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 393.390 2486.280 393.670 2486.560 ;
      LAYER met3 ;
        RECT 393.365 2486.570 393.695 2486.585 ;
        RECT 410.000 2486.570 414.000 2486.720 ;
        RECT 393.365 2486.270 414.000 2486.570 ;
        RECT 393.365 2486.255 393.695 2486.270 ;
        RECT 410.000 2486.120 414.000 2486.270 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1919.650 496.980 1919.970 497.040 ;
        RECT 1924.710 496.980 1925.030 497.040 ;
        RECT 1919.650 496.840 1925.030 496.980 ;
        RECT 1919.650 496.780 1919.970 496.840 ;
        RECT 1924.710 496.780 1925.030 496.840 ;
        RECT 1924.710 258.640 1925.030 258.700 ;
        RECT 2380.570 258.640 2380.890 258.700 ;
        RECT 1924.710 258.500 2380.890 258.640 ;
        RECT 1924.710 258.440 1925.030 258.500 ;
        RECT 2380.570 258.440 2380.890 258.500 ;
      LAYER via ;
        RECT 1919.680 496.780 1919.940 497.040 ;
        RECT 1924.740 496.780 1925.000 497.040 ;
        RECT 1924.740 258.440 1925.000 258.700 ;
        RECT 2380.600 258.440 2380.860 258.700 ;
      LAYER met2 ;
        RECT 1919.810 510.340 1920.090 514.000 ;
        RECT 1919.740 510.000 1920.090 510.340 ;
        RECT 1919.740 497.070 1919.880 510.000 ;
        RECT 1919.680 496.750 1919.940 497.070 ;
        RECT 1924.740 496.750 1925.000 497.070 ;
        RECT 1924.800 258.730 1924.940 496.750 ;
        RECT 1924.740 258.410 1925.000 258.730 ;
        RECT 2380.600 258.410 2380.860 258.730 ;
        RECT 2380.660 17.410 2380.800 258.410 ;
        RECT 2380.660 17.270 2381.720 17.410 ;
        RECT 2381.580 2.400 2381.720 17.270 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2400.350 509.220 2400.670 509.280 ;
        RECT 2512.590 509.220 2512.910 509.280 ;
        RECT 2400.350 509.080 2512.910 509.220 ;
        RECT 2400.350 509.020 2400.670 509.080 ;
        RECT 2512.590 509.020 2512.910 509.080 ;
      LAYER via ;
        RECT 2400.380 509.020 2400.640 509.280 ;
        RECT 2512.620 509.020 2512.880 509.280 ;
      LAYER met2 ;
        RECT 2512.610 2055.115 2512.890 2055.485 ;
        RECT 2512.680 509.310 2512.820 2055.115 ;
        RECT 2400.380 508.990 2400.640 509.310 ;
        RECT 2512.620 508.990 2512.880 509.310 ;
        RECT 2400.440 481.850 2400.580 508.990 ;
        RECT 2400.440 481.710 2401.040 481.850 ;
        RECT 2400.900 17.410 2401.040 481.710 ;
        RECT 2399.520 17.270 2401.040 17.410 ;
        RECT 2399.520 2.400 2399.660 17.270 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 2512.610 2055.160 2512.890 2055.440 ;
      LAYER met3 ;
        RECT 2506.000 2055.450 2510.000 2055.600 ;
        RECT 2512.585 2055.450 2512.915 2055.465 ;
        RECT 2506.000 2055.150 2512.915 2055.450 ;
        RECT 2506.000 2055.000 2510.000 2055.150 ;
        RECT 2512.585 2055.135 2512.915 2055.150 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 469.345 16.065 469.515 20.315 ;
        RECT 517.185 16.065 517.355 20.315 ;
        RECT 565.945 16.405 566.115 20.315 ;
        RECT 613.785 16.405 613.955 20.315 ;
        RECT 662.545 16.405 662.715 20.315 ;
        RECT 734.765 16.405 734.935 20.315 ;
        RECT 786.745 16.745 786.915 20.315 ;
      LAYER mcon ;
        RECT 469.345 20.145 469.515 20.315 ;
        RECT 517.185 20.145 517.355 20.315 ;
        RECT 565.945 20.145 566.115 20.315 ;
        RECT 613.785 20.145 613.955 20.315 ;
        RECT 662.545 20.145 662.715 20.315 ;
        RECT 734.765 20.145 734.935 20.315 ;
        RECT 786.745 20.145 786.915 20.315 ;
      LAYER met1 ;
        RECT 399.350 511.940 399.670 512.000 ;
        RECT 424.190 511.940 424.510 512.000 ;
        RECT 399.350 511.800 424.510 511.940 ;
        RECT 399.350 511.740 399.670 511.800 ;
        RECT 424.190 511.740 424.510 511.800 ;
        RECT 424.190 20.300 424.510 20.360 ;
        RECT 469.285 20.300 469.575 20.345 ;
        RECT 424.190 20.160 469.575 20.300 ;
        RECT 424.190 20.100 424.510 20.160 ;
        RECT 469.285 20.115 469.575 20.160 ;
        RECT 517.125 20.300 517.415 20.345 ;
        RECT 565.885 20.300 566.175 20.345 ;
        RECT 517.125 20.160 566.175 20.300 ;
        RECT 517.125 20.115 517.415 20.160 ;
        RECT 565.885 20.115 566.175 20.160 ;
        RECT 613.725 20.300 614.015 20.345 ;
        RECT 662.485 20.300 662.775 20.345 ;
        RECT 613.725 20.160 662.775 20.300 ;
        RECT 613.725 20.115 614.015 20.160 ;
        RECT 662.485 20.115 662.775 20.160 ;
        RECT 734.705 20.300 734.995 20.345 ;
        RECT 786.685 20.300 786.975 20.345 ;
        RECT 734.705 20.160 786.975 20.300 ;
        RECT 734.705 20.115 734.995 20.160 ;
        RECT 786.685 20.115 786.975 20.160 ;
        RECT 786.685 16.900 786.975 16.945 ;
        RECT 793.570 16.900 793.890 16.960 ;
        RECT 786.685 16.760 793.890 16.900 ;
        RECT 786.685 16.715 786.975 16.760 ;
        RECT 793.570 16.700 793.890 16.760 ;
        RECT 565.885 16.560 566.175 16.605 ;
        RECT 613.725 16.560 614.015 16.605 ;
        RECT 565.885 16.420 614.015 16.560 ;
        RECT 565.885 16.375 566.175 16.420 ;
        RECT 613.725 16.375 614.015 16.420 ;
        RECT 662.485 16.560 662.775 16.605 ;
        RECT 734.705 16.560 734.995 16.605 ;
        RECT 662.485 16.420 734.995 16.560 ;
        RECT 662.485 16.375 662.775 16.420 ;
        RECT 734.705 16.375 734.995 16.420 ;
        RECT 469.285 16.220 469.575 16.265 ;
        RECT 517.125 16.220 517.415 16.265 ;
        RECT 469.285 16.080 517.415 16.220 ;
        RECT 469.285 16.035 469.575 16.080 ;
        RECT 517.125 16.035 517.415 16.080 ;
      LAYER via ;
        RECT 399.380 511.740 399.640 512.000 ;
        RECT 424.220 511.740 424.480 512.000 ;
        RECT 424.220 20.100 424.480 20.360 ;
        RECT 793.600 16.700 793.860 16.960 ;
      LAYER met2 ;
        RECT 399.370 1955.835 399.650 1956.205 ;
        RECT 399.440 512.030 399.580 1955.835 ;
        RECT 399.380 511.710 399.640 512.030 ;
        RECT 424.220 511.710 424.480 512.030 ;
        RECT 424.280 20.390 424.420 511.710 ;
        RECT 424.220 20.070 424.480 20.390 ;
        RECT 793.600 16.670 793.860 16.990 ;
        RECT 793.660 2.400 793.800 16.670 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 399.370 1955.880 399.650 1956.160 ;
      LAYER met3 ;
        RECT 399.345 1956.170 399.675 1956.185 ;
        RECT 410.000 1956.170 414.000 1956.320 ;
        RECT 399.345 1955.870 414.000 1956.170 ;
        RECT 399.345 1955.855 399.675 1955.870 ;
        RECT 410.000 1955.720 414.000 1955.870 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 342.280 641.630 342.340 ;
        RECT 1449.070 342.280 1449.390 342.340 ;
        RECT 641.310 342.140 1449.390 342.280 ;
        RECT 641.310 342.080 641.630 342.140 ;
        RECT 1449.070 342.080 1449.390 342.140 ;
        RECT 639.010 16.900 639.330 16.960 ;
        RECT 641.310 16.900 641.630 16.960 ;
        RECT 639.010 16.760 641.630 16.900 ;
        RECT 639.010 16.700 639.330 16.760 ;
        RECT 641.310 16.700 641.630 16.760 ;
      LAYER via ;
        RECT 641.340 342.080 641.600 342.340 ;
        RECT 1449.100 342.080 1449.360 342.340 ;
        RECT 639.040 16.700 639.300 16.960 ;
        RECT 641.340 16.700 641.600 16.960 ;
      LAYER met2 ;
        RECT 1449.690 510.410 1449.970 514.000 ;
        RECT 1449.160 510.270 1449.970 510.410 ;
        RECT 1449.160 342.370 1449.300 510.270 ;
        RECT 1449.690 510.000 1449.970 510.270 ;
        RECT 641.340 342.050 641.600 342.370 ;
        RECT 1449.100 342.050 1449.360 342.370 ;
        RECT 641.400 16.990 641.540 342.050 ;
        RECT 639.040 16.670 639.300 16.990 ;
        RECT 641.340 16.670 641.600 16.990 ;
        RECT 639.100 2.400 639.240 16.670 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2388.850 499.700 2389.170 499.760 ;
        RECT 2393.450 499.700 2393.770 499.760 ;
        RECT 2388.850 499.560 2393.770 499.700 ;
        RECT 2388.850 499.500 2389.170 499.560 ;
        RECT 2393.450 499.500 2393.770 499.560 ;
        RECT 2393.450 107.000 2393.770 107.060 ;
        RECT 2421.970 107.000 2422.290 107.060 ;
        RECT 2393.450 106.860 2422.290 107.000 ;
        RECT 2393.450 106.800 2393.770 106.860 ;
        RECT 2421.970 106.800 2422.290 106.860 ;
      LAYER via ;
        RECT 2388.880 499.500 2389.140 499.760 ;
        RECT 2393.480 499.500 2393.740 499.760 ;
        RECT 2393.480 106.800 2393.740 107.060 ;
        RECT 2422.000 106.800 2422.260 107.060 ;
      LAYER met2 ;
        RECT 2389.010 510.340 2389.290 514.000 ;
        RECT 2388.940 510.000 2389.290 510.340 ;
        RECT 2388.940 499.790 2389.080 510.000 ;
        RECT 2388.880 499.470 2389.140 499.790 ;
        RECT 2393.480 499.470 2393.740 499.790 ;
        RECT 2393.540 107.090 2393.680 499.470 ;
        RECT 2393.480 106.770 2393.740 107.090 ;
        RECT 2422.000 106.770 2422.260 107.090 ;
        RECT 2422.060 16.730 2422.200 106.770 ;
        RECT 2422.060 16.590 2423.120 16.730 ;
        RECT 2422.980 2.400 2423.120 16.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2440.905 48.365 2441.075 62.475 ;
      LAYER mcon ;
        RECT 2440.905 62.305 2441.075 62.475 ;
      LAYER met1 ;
        RECT 2515.350 665.280 2515.670 665.340 ;
        RECT 2542.490 665.280 2542.810 665.340 ;
        RECT 2515.350 665.140 2542.810 665.280 ;
        RECT 2515.350 665.080 2515.670 665.140 ;
        RECT 2542.490 665.080 2542.810 665.140 ;
        RECT 2442.210 509.560 2442.530 509.620 ;
        RECT 2542.490 509.560 2542.810 509.620 ;
        RECT 2442.210 509.420 2542.810 509.560 ;
        RECT 2442.210 509.360 2442.530 509.420 ;
        RECT 2542.490 509.360 2542.810 509.420 ;
        RECT 2440.845 62.460 2441.135 62.505 ;
        RECT 2442.210 62.460 2442.530 62.520 ;
        RECT 2440.845 62.320 2442.530 62.460 ;
        RECT 2440.845 62.275 2441.135 62.320 ;
        RECT 2442.210 62.260 2442.530 62.320 ;
        RECT 2440.830 48.520 2441.150 48.580 ;
        RECT 2440.635 48.380 2441.150 48.520 ;
        RECT 2440.830 48.320 2441.150 48.380 ;
      LAYER via ;
        RECT 2515.380 665.080 2515.640 665.340 ;
        RECT 2542.520 665.080 2542.780 665.340 ;
        RECT 2442.240 509.360 2442.500 509.620 ;
        RECT 2542.520 509.360 2542.780 509.620 ;
        RECT 2442.240 62.260 2442.500 62.520 ;
        RECT 2440.860 48.320 2441.120 48.580 ;
      LAYER met2 ;
        RECT 2515.370 667.915 2515.650 668.285 ;
        RECT 2515.440 665.370 2515.580 667.915 ;
        RECT 2515.380 665.050 2515.640 665.370 ;
        RECT 2542.520 665.050 2542.780 665.370 ;
        RECT 2542.580 509.650 2542.720 665.050 ;
        RECT 2442.240 509.330 2442.500 509.650 ;
        RECT 2542.520 509.330 2542.780 509.650 ;
        RECT 2442.300 62.550 2442.440 509.330 ;
        RECT 2442.240 62.230 2442.500 62.550 ;
        RECT 2440.860 48.290 2441.120 48.610 ;
        RECT 2440.920 2.400 2441.060 48.290 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
      LAYER via2 ;
        RECT 2515.370 667.960 2515.650 668.240 ;
      LAYER met3 ;
        RECT 2506.000 668.250 2510.000 668.400 ;
        RECT 2515.345 668.250 2515.675 668.265 ;
        RECT 2506.000 667.950 2515.675 668.250 ;
        RECT 2506.000 667.800 2510.000 667.950 ;
        RECT 2515.345 667.935 2515.675 667.950 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 684.090 501.400 684.410 501.460 ;
        RECT 689.610 501.400 689.930 501.460 ;
        RECT 684.090 501.260 689.930 501.400 ;
        RECT 684.090 501.200 684.410 501.260 ;
        RECT 689.610 501.200 689.930 501.260 ;
        RECT 689.610 141.680 689.930 141.740 ;
        RECT 2456.470 141.680 2456.790 141.740 ;
        RECT 689.610 141.540 2456.790 141.680 ;
        RECT 689.610 141.480 689.930 141.540 ;
        RECT 2456.470 141.480 2456.790 141.540 ;
      LAYER via ;
        RECT 684.120 501.200 684.380 501.460 ;
        RECT 689.640 501.200 689.900 501.460 ;
        RECT 689.640 141.480 689.900 141.740 ;
        RECT 2456.500 141.480 2456.760 141.740 ;
      LAYER met2 ;
        RECT 684.250 510.340 684.530 514.000 ;
        RECT 684.180 510.000 684.530 510.340 ;
        RECT 684.180 501.490 684.320 510.000 ;
        RECT 684.120 501.170 684.380 501.490 ;
        RECT 689.640 501.170 689.900 501.490 ;
        RECT 689.700 141.770 689.840 501.170 ;
        RECT 689.640 141.450 689.900 141.770 ;
        RECT 2456.500 141.450 2456.760 141.770 ;
        RECT 2456.560 3.130 2456.700 141.450 ;
        RECT 2456.560 2.990 2459.000 3.130 ;
        RECT 2458.860 2.400 2459.000 2.990 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 203.560 524.330 203.620 ;
        RECT 2470.270 203.560 2470.590 203.620 ;
        RECT 524.010 203.420 2470.590 203.560 ;
        RECT 524.010 203.360 524.330 203.420 ;
        RECT 2470.270 203.360 2470.590 203.420 ;
        RECT 2470.270 37.980 2470.590 38.040 ;
        RECT 2476.710 37.980 2477.030 38.040 ;
        RECT 2470.270 37.840 2477.030 37.980 ;
        RECT 2470.270 37.780 2470.590 37.840 ;
        RECT 2476.710 37.780 2477.030 37.840 ;
      LAYER via ;
        RECT 524.040 203.360 524.300 203.620 ;
        RECT 2470.300 203.360 2470.560 203.620 ;
        RECT 2470.300 37.780 2470.560 38.040 ;
        RECT 2476.740 37.780 2477.000 38.040 ;
      LAYER met2 ;
        RECT 523.250 510.410 523.530 514.000 ;
        RECT 523.250 510.270 524.240 510.410 ;
        RECT 523.250 510.000 523.530 510.270 ;
        RECT 524.100 203.650 524.240 510.270 ;
        RECT 524.040 203.330 524.300 203.650 ;
        RECT 2470.300 203.330 2470.560 203.650 ;
        RECT 2470.360 38.070 2470.500 203.330 ;
        RECT 2470.300 37.750 2470.560 38.070 ;
        RECT 2476.740 37.750 2477.000 38.070 ;
        RECT 2476.800 2.400 2476.940 37.750 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1725.400 2520.730 1725.460 ;
        RECT 2569.170 1725.400 2569.490 1725.460 ;
        RECT 2520.410 1725.260 2569.490 1725.400 ;
        RECT 2520.410 1725.200 2520.730 1725.260 ;
        RECT 2569.170 1725.200 2569.490 1725.260 ;
        RECT 2497.410 509.900 2497.730 509.960 ;
        RECT 2569.170 509.900 2569.490 509.960 ;
        RECT 2497.410 509.760 2569.490 509.900 ;
        RECT 2497.410 509.700 2497.730 509.760 ;
        RECT 2569.170 509.700 2569.490 509.760 ;
        RECT 2494.650 20.300 2494.970 20.360 ;
        RECT 2497.410 20.300 2497.730 20.360 ;
        RECT 2494.650 20.160 2497.730 20.300 ;
        RECT 2494.650 20.100 2494.970 20.160 ;
        RECT 2497.410 20.100 2497.730 20.160 ;
      LAYER via ;
        RECT 2520.440 1725.200 2520.700 1725.460 ;
        RECT 2569.200 1725.200 2569.460 1725.460 ;
        RECT 2497.440 509.700 2497.700 509.960 ;
        RECT 2569.200 509.700 2569.460 509.960 ;
        RECT 2494.680 20.100 2494.940 20.360 ;
        RECT 2497.440 20.100 2497.700 20.360 ;
      LAYER met2 ;
        RECT 2520.430 1727.355 2520.710 1727.725 ;
        RECT 2520.500 1725.490 2520.640 1727.355 ;
        RECT 2520.440 1725.170 2520.700 1725.490 ;
        RECT 2569.200 1725.170 2569.460 1725.490 ;
        RECT 2569.260 509.990 2569.400 1725.170 ;
        RECT 2497.440 509.670 2497.700 509.990 ;
        RECT 2569.200 509.670 2569.460 509.990 ;
        RECT 2497.500 20.390 2497.640 509.670 ;
        RECT 2494.680 20.070 2494.940 20.390 ;
        RECT 2497.440 20.070 2497.700 20.390 ;
        RECT 2494.740 2.400 2494.880 20.070 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1727.400 2520.710 1727.680 ;
      LAYER met3 ;
        RECT 2506.000 1727.690 2510.000 1727.840 ;
        RECT 2520.405 1727.690 2520.735 1727.705 ;
        RECT 2506.000 1727.390 2520.735 1727.690 ;
        RECT 2506.000 1727.240 2510.000 1727.390 ;
        RECT 2520.405 1727.375 2520.735 1727.390 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2512.205 2.805 2512.375 48.195 ;
      LAYER mcon ;
        RECT 2512.205 48.025 2512.375 48.195 ;
      LAYER met1 ;
        RECT 403.950 93.400 404.270 93.460 ;
        RECT 2511.670 93.400 2511.990 93.460 ;
        RECT 403.950 93.260 2511.990 93.400 ;
        RECT 403.950 93.200 404.270 93.260 ;
        RECT 2511.670 93.200 2511.990 93.260 ;
        RECT 2511.670 62.120 2511.990 62.180 ;
        RECT 2512.590 62.120 2512.910 62.180 ;
        RECT 2511.670 61.980 2512.910 62.120 ;
        RECT 2511.670 61.920 2511.990 61.980 ;
        RECT 2512.590 61.920 2512.910 61.980 ;
        RECT 2512.145 48.180 2512.435 48.225 ;
        RECT 2512.590 48.180 2512.910 48.240 ;
        RECT 2512.145 48.040 2512.910 48.180 ;
        RECT 2512.145 47.995 2512.435 48.040 ;
        RECT 2512.590 47.980 2512.910 48.040 ;
        RECT 2512.130 2.960 2512.450 3.020 ;
        RECT 2511.935 2.820 2512.450 2.960 ;
        RECT 2512.130 2.760 2512.450 2.820 ;
      LAYER via ;
        RECT 403.980 93.200 404.240 93.460 ;
        RECT 2511.700 93.200 2511.960 93.460 ;
        RECT 2511.700 61.920 2511.960 62.180 ;
        RECT 2512.620 61.920 2512.880 62.180 ;
        RECT 2512.620 47.980 2512.880 48.240 ;
        RECT 2512.160 2.760 2512.420 3.020 ;
      LAYER met2 ;
        RECT 403.970 1006.555 404.250 1006.925 ;
        RECT 404.040 93.490 404.180 1006.555 ;
        RECT 403.980 93.170 404.240 93.490 ;
        RECT 2511.700 93.170 2511.960 93.490 ;
        RECT 2511.760 62.210 2511.900 93.170 ;
        RECT 2511.700 61.890 2511.960 62.210 ;
        RECT 2512.620 61.890 2512.880 62.210 ;
        RECT 2512.680 48.270 2512.820 61.890 ;
        RECT 2512.620 47.950 2512.880 48.270 ;
        RECT 2512.160 2.730 2512.420 3.050 ;
        RECT 2512.220 2.400 2512.360 2.730 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 403.970 1006.600 404.250 1006.880 ;
      LAYER met3 ;
        RECT 403.945 1006.890 404.275 1006.905 ;
        RECT 410.000 1006.890 414.000 1007.040 ;
        RECT 403.945 1006.590 414.000 1006.890 ;
        RECT 403.945 1006.575 404.275 1006.590 ;
        RECT 410.000 1006.440 414.000 1006.590 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.150 279.720 1103.470 279.780 ;
        RECT 2525.470 279.720 2525.790 279.780 ;
        RECT 1103.150 279.580 2525.790 279.720 ;
        RECT 1103.150 279.520 1103.470 279.580 ;
        RECT 2525.470 279.520 2525.790 279.580 ;
        RECT 2525.470 2.960 2525.790 3.020 ;
        RECT 2530.070 2.960 2530.390 3.020 ;
        RECT 2525.470 2.820 2530.390 2.960 ;
        RECT 2525.470 2.760 2525.790 2.820 ;
        RECT 2530.070 2.760 2530.390 2.820 ;
      LAYER via ;
        RECT 1103.180 279.520 1103.440 279.780 ;
        RECT 2525.500 279.520 2525.760 279.780 ;
        RECT 2525.500 2.760 2525.760 3.020 ;
        RECT 2530.100 2.760 2530.360 3.020 ;
      LAYER met2 ;
        RECT 1103.770 510.410 1104.050 514.000 ;
        RECT 1103.240 510.270 1104.050 510.410 ;
        RECT 1103.240 279.810 1103.380 510.270 ;
        RECT 1103.770 510.000 1104.050 510.270 ;
        RECT 1103.180 279.490 1103.440 279.810 ;
        RECT 2525.500 279.490 2525.760 279.810 ;
        RECT 2525.560 3.050 2525.700 279.490 ;
        RECT 2525.500 2.730 2525.760 3.050 ;
        RECT 2530.100 2.730 2530.360 3.050 ;
        RECT 2530.160 2.400 2530.300 2.730 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2546.190 347.635 2546.470 348.005 ;
        RECT 2546.260 3.130 2546.400 347.635 ;
        RECT 2546.260 2.990 2548.240 3.130 ;
        RECT 2548.100 2.400 2548.240 2.990 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
      LAYER via2 ;
        RECT 2546.190 347.680 2546.470 347.960 ;
      LAYER met3 ;
        RECT 381.150 2686.490 381.530 2686.500 ;
        RECT 410.000 2686.490 414.000 2686.640 ;
        RECT 381.150 2686.190 414.000 2686.490 ;
        RECT 381.150 2686.180 381.530 2686.190 ;
        RECT 410.000 2686.040 414.000 2686.190 ;
        RECT 381.150 347.970 381.530 347.980 ;
        RECT 2546.165 347.970 2546.495 347.985 ;
        RECT 381.150 347.670 2546.495 347.970 ;
        RECT 381.150 347.660 381.530 347.670 ;
        RECT 2546.165 347.655 2546.495 347.670 ;
      LAYER via3 ;
        RECT 381.180 2686.180 381.500 2686.500 ;
        RECT 381.180 347.660 381.500 347.980 ;
      LAYER met4 ;
        RECT 381.175 2686.175 381.505 2686.505 ;
        RECT 381.190 347.985 381.490 2686.175 ;
        RECT 381.175 347.655 381.505 347.985 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2557.210 20.640 2557.530 20.700 ;
        RECT 2565.950 20.640 2566.270 20.700 ;
        RECT 2557.210 20.500 2566.270 20.640 ;
        RECT 2557.210 20.440 2557.530 20.500 ;
        RECT 2565.950 20.440 2566.270 20.500 ;
      LAYER via ;
        RECT 2557.240 20.440 2557.500 20.700 ;
        RECT 2565.980 20.440 2566.240 20.700 ;
      LAYER met2 ;
        RECT 2557.230 437.395 2557.510 437.765 ;
        RECT 2557.300 20.730 2557.440 437.395 ;
        RECT 2557.240 20.410 2557.500 20.730 ;
        RECT 2565.980 20.410 2566.240 20.730 ;
        RECT 2566.040 2.400 2566.180 20.410 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
      LAYER via2 ;
        RECT 2557.230 437.440 2557.510 437.720 ;
      LAYER met3 ;
        RECT 398.630 2614.410 399.010 2614.420 ;
        RECT 410.000 2614.410 414.000 2614.560 ;
        RECT 398.630 2614.110 414.000 2614.410 ;
        RECT 398.630 2614.100 399.010 2614.110 ;
        RECT 410.000 2613.960 414.000 2614.110 ;
        RECT 398.630 437.730 399.010 437.740 ;
        RECT 2557.205 437.730 2557.535 437.745 ;
        RECT 398.630 437.430 2557.535 437.730 ;
        RECT 398.630 437.420 399.010 437.430 ;
        RECT 2557.205 437.415 2557.535 437.430 ;
      LAYER via3 ;
        RECT 398.660 2614.100 398.980 2614.420 ;
        RECT 398.660 437.420 398.980 437.740 ;
      LAYER met4 ;
        RECT 398.655 2614.095 398.985 2614.425 ;
        RECT 398.670 437.745 398.970 2614.095 ;
        RECT 398.655 437.415 398.985 437.745 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 322.530 2539.360 322.850 2539.420 ;
        RECT 393.370 2539.360 393.690 2539.420 ;
        RECT 322.530 2539.220 393.690 2539.360 ;
        RECT 322.530 2539.160 322.850 2539.220 ;
        RECT 393.370 2539.160 393.690 2539.220 ;
        RECT 322.530 59.060 322.850 59.120 ;
        RECT 2581.590 59.060 2581.910 59.120 ;
        RECT 322.530 58.920 2581.910 59.060 ;
        RECT 322.530 58.860 322.850 58.920 ;
        RECT 2581.590 58.860 2581.910 58.920 ;
      LAYER via ;
        RECT 322.560 2539.160 322.820 2539.420 ;
        RECT 393.400 2539.160 393.660 2539.420 ;
        RECT 322.560 58.860 322.820 59.120 ;
        RECT 2581.620 58.860 2581.880 59.120 ;
      LAYER met2 ;
        RECT 393.390 2540.635 393.670 2541.005 ;
        RECT 393.460 2539.450 393.600 2540.635 ;
        RECT 322.560 2539.130 322.820 2539.450 ;
        RECT 393.400 2539.130 393.660 2539.450 ;
        RECT 322.620 59.150 322.760 2539.130 ;
        RECT 322.560 58.830 322.820 59.150 ;
        RECT 2581.620 58.830 2581.880 59.150 ;
        RECT 2581.680 15.370 2581.820 58.830 ;
        RECT 2581.680 15.230 2583.660 15.370 ;
        RECT 2583.520 3.130 2583.660 15.230 ;
        RECT 2583.520 2.990 2584.120 3.130 ;
        RECT 2583.980 2.400 2584.120 2.990 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
      LAYER via2 ;
        RECT 393.390 2540.680 393.670 2540.960 ;
      LAYER met3 ;
        RECT 393.365 2540.970 393.695 2540.985 ;
        RECT 410.000 2540.970 414.000 2541.120 ;
        RECT 393.365 2540.670 414.000 2540.970 ;
        RECT 393.365 2540.655 393.695 2540.670 ;
        RECT 410.000 2540.520 414.000 2540.670 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2358.490 3031.680 2358.810 3031.740 ;
        RECT 2574.690 3031.680 2575.010 3031.740 ;
        RECT 2358.490 3031.540 2575.010 3031.680 ;
        RECT 2358.490 3031.480 2358.810 3031.540 ;
        RECT 2574.690 3031.480 2575.010 3031.540 ;
        RECT 817.490 15.200 817.810 15.260 ;
        RECT 820.710 15.200 821.030 15.260 ;
        RECT 817.490 15.060 821.030 15.200 ;
        RECT 817.490 15.000 817.810 15.060 ;
        RECT 820.710 15.000 821.030 15.060 ;
      LAYER via ;
        RECT 2358.520 3031.480 2358.780 3031.740 ;
        RECT 2574.720 3031.480 2574.980 3031.740 ;
        RECT 817.520 15.000 817.780 15.260 ;
        RECT 820.740 15.000 821.000 15.260 ;
      LAYER met2 ;
        RECT 2358.520 3031.450 2358.780 3031.770 ;
        RECT 2574.720 3031.450 2574.980 3031.770 ;
        RECT 2358.580 3010.000 2358.720 3031.450 ;
        RECT 2358.580 3009.340 2358.930 3010.000 ;
        RECT 2358.650 3006.000 2358.930 3009.340 ;
        RECT 2574.780 479.245 2574.920 3031.450 ;
        RECT 820.730 478.875 821.010 479.245 ;
        RECT 2574.710 478.875 2574.990 479.245 ;
        RECT 820.800 15.290 820.940 478.875 ;
        RECT 817.520 14.970 817.780 15.290 ;
        RECT 820.740 14.970 821.000 15.290 ;
        RECT 817.580 2.400 817.720 14.970 ;
        RECT 817.370 -4.800 817.930 2.400 ;
      LAYER via2 ;
        RECT 820.730 478.920 821.010 479.200 ;
        RECT 2574.710 478.920 2574.990 479.200 ;
      LAYER met3 ;
        RECT 820.705 479.210 821.035 479.225 ;
        RECT 2574.685 479.210 2575.015 479.225 ;
        RECT 820.705 478.910 2575.015 479.210 ;
        RECT 820.705 478.895 821.035 478.910 ;
        RECT 2574.685 478.895 2575.015 478.910 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1537.850 196.760 1538.170 196.820 ;
        RECT 2602.290 196.760 2602.610 196.820 ;
        RECT 1537.850 196.620 2602.610 196.760 ;
        RECT 1537.850 196.560 1538.170 196.620 ;
        RECT 2602.290 196.560 2602.610 196.620 ;
      LAYER via ;
        RECT 1537.880 196.560 1538.140 196.820 ;
        RECT 2602.320 196.560 2602.580 196.820 ;
      LAYER met2 ;
        RECT 1536.170 510.410 1536.450 514.000 ;
        RECT 1536.170 510.270 1538.080 510.410 ;
        RECT 1536.170 510.000 1536.450 510.270 ;
        RECT 1537.940 196.850 1538.080 510.270 ;
        RECT 1537.880 196.530 1538.140 196.850 ;
        RECT 2602.320 196.530 2602.580 196.850 ;
        RECT 2602.380 17.410 2602.520 196.530 ;
        RECT 2601.460 17.270 2602.520 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 432.010 3029.640 432.330 3029.700 ;
        RECT 2615.170 3029.640 2615.490 3029.700 ;
        RECT 432.010 3029.500 2615.490 3029.640 ;
        RECT 432.010 3029.440 432.330 3029.500 ;
        RECT 2615.170 3029.440 2615.490 3029.500 ;
      LAYER via ;
        RECT 432.040 3029.440 432.300 3029.700 ;
        RECT 2615.200 3029.440 2615.460 3029.700 ;
      LAYER met2 ;
        RECT 432.040 3029.410 432.300 3029.730 ;
        RECT 2615.200 3029.410 2615.460 3029.730 ;
        RECT 432.100 3010.000 432.240 3029.410 ;
        RECT 432.100 3009.340 432.450 3010.000 ;
        RECT 432.170 3006.000 432.450 3009.340 ;
        RECT 2615.260 16.730 2615.400 3029.410 ;
        RECT 2615.260 16.590 2619.540 16.730 ;
        RECT 2619.400 2.400 2619.540 16.590 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.150 286.520 1724.470 286.580 ;
        RECT 2635.870 286.520 2636.190 286.580 ;
        RECT 1724.150 286.380 2636.190 286.520 ;
        RECT 1724.150 286.320 1724.470 286.380 ;
        RECT 2635.870 286.320 2636.190 286.380 ;
      LAYER via ;
        RECT 1724.180 286.320 1724.440 286.580 ;
        RECT 2635.900 286.320 2636.160 286.580 ;
      LAYER met2 ;
        RECT 1722.010 510.410 1722.290 514.000 ;
        RECT 1722.010 510.270 1724.380 510.410 ;
        RECT 1722.010 510.000 1722.290 510.270 ;
        RECT 1724.240 286.610 1724.380 510.270 ;
        RECT 1724.180 286.290 1724.440 286.610 ;
        RECT 2635.900 286.290 2636.160 286.610 ;
        RECT 2635.960 16.730 2636.100 286.290 ;
        RECT 2635.960 16.590 2637.480 16.730 ;
        RECT 2637.340 2.400 2637.480 16.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 329.430 2063.360 329.750 2063.420 ;
        RECT 393.370 2063.360 393.690 2063.420 ;
        RECT 329.430 2063.220 393.690 2063.360 ;
        RECT 329.430 2063.160 329.750 2063.220 ;
        RECT 393.370 2063.160 393.690 2063.220 ;
        RECT 329.430 58.720 329.750 58.780 ;
        RECT 2649.670 58.720 2649.990 58.780 ;
        RECT 329.430 58.580 2649.990 58.720 ;
        RECT 329.430 58.520 329.750 58.580 ;
        RECT 2649.670 58.520 2649.990 58.580 ;
      LAYER via ;
        RECT 329.460 2063.160 329.720 2063.420 ;
        RECT 393.400 2063.160 393.660 2063.420 ;
        RECT 329.460 58.520 329.720 58.780 ;
        RECT 2649.700 58.520 2649.960 58.780 ;
      LAYER met2 ;
        RECT 393.390 2065.995 393.670 2066.365 ;
        RECT 393.460 2063.450 393.600 2065.995 ;
        RECT 329.460 2063.130 329.720 2063.450 ;
        RECT 393.400 2063.130 393.660 2063.450 ;
        RECT 329.520 58.810 329.660 2063.130 ;
        RECT 329.460 58.490 329.720 58.810 ;
        RECT 2649.700 58.490 2649.960 58.810 ;
        RECT 2649.760 17.410 2649.900 58.490 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 393.390 2066.040 393.670 2066.320 ;
      LAYER met3 ;
        RECT 393.365 2066.330 393.695 2066.345 ;
        RECT 410.000 2066.330 414.000 2066.480 ;
        RECT 393.365 2066.030 414.000 2066.330 ;
        RECT 393.365 2066.015 393.695 2066.030 ;
        RECT 410.000 2065.880 414.000 2066.030 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2260.050 3019.100 2260.370 3019.160 ;
        RECT 2510.290 3019.100 2510.610 3019.160 ;
        RECT 2260.050 3018.960 2510.610 3019.100 ;
        RECT 2260.050 3018.900 2260.370 3018.960 ;
        RECT 2510.290 3018.900 2510.610 3018.960 ;
        RECT 2510.290 2991.220 2510.610 2991.280 ;
        RECT 2670.370 2991.220 2670.690 2991.280 ;
        RECT 2510.290 2991.080 2670.690 2991.220 ;
        RECT 2510.290 2991.020 2510.610 2991.080 ;
        RECT 2670.370 2991.020 2670.690 2991.080 ;
      LAYER via ;
        RECT 2260.080 3018.900 2260.340 3019.160 ;
        RECT 2510.320 3018.900 2510.580 3019.160 ;
        RECT 2510.320 2991.020 2510.580 2991.280 ;
        RECT 2670.400 2991.020 2670.660 2991.280 ;
      LAYER met2 ;
        RECT 2260.080 3018.870 2260.340 3019.190 ;
        RECT 2510.320 3018.870 2510.580 3019.190 ;
        RECT 2260.140 3010.000 2260.280 3018.870 ;
        RECT 2260.140 3009.340 2260.490 3010.000 ;
        RECT 2260.210 3006.000 2260.490 3009.340 ;
        RECT 2510.380 2991.310 2510.520 3018.870 ;
        RECT 2510.320 2990.990 2510.580 2991.310 ;
        RECT 2670.400 2990.990 2670.660 2991.310 ;
        RECT 2670.460 17.410 2670.600 2990.990 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.250 2735.880 2522.570 2735.940 ;
        RECT 2684.170 2735.880 2684.490 2735.940 ;
        RECT 2522.250 2735.740 2684.490 2735.880 ;
        RECT 2522.250 2735.680 2522.570 2735.740 ;
        RECT 2684.170 2735.680 2684.490 2735.740 ;
        RECT 2684.170 11.800 2684.490 11.860 ;
        RECT 2690.610 11.800 2690.930 11.860 ;
        RECT 2684.170 11.660 2690.930 11.800 ;
        RECT 2684.170 11.600 2684.490 11.660 ;
        RECT 2690.610 11.600 2690.930 11.660 ;
      LAYER via ;
        RECT 2522.280 2735.680 2522.540 2735.940 ;
        RECT 2684.200 2735.680 2684.460 2735.940 ;
        RECT 2684.200 11.600 2684.460 11.860 ;
        RECT 2690.640 11.600 2690.900 11.860 ;
      LAYER met2 ;
        RECT 2522.270 2877.915 2522.550 2878.285 ;
        RECT 2522.340 2735.970 2522.480 2877.915 ;
        RECT 2522.280 2735.650 2522.540 2735.970 ;
        RECT 2684.200 2735.650 2684.460 2735.970 ;
        RECT 2684.260 11.890 2684.400 2735.650 ;
        RECT 2684.200 11.570 2684.460 11.890 ;
        RECT 2690.640 11.570 2690.900 11.890 ;
        RECT 2690.700 2.400 2690.840 11.570 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 2522.270 2877.960 2522.550 2878.240 ;
      LAYER met3 ;
        RECT 2506.000 2878.250 2510.000 2878.400 ;
        RECT 2522.245 2878.250 2522.575 2878.265 ;
        RECT 2506.000 2877.950 2522.575 2878.250 ;
        RECT 2506.000 2877.800 2510.000 2877.950 ;
        RECT 2522.245 2877.935 2522.575 2877.950 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1906.770 496.980 1907.090 497.040 ;
        RECT 1910.910 496.980 1911.230 497.040 ;
        RECT 1906.770 496.840 1911.230 496.980 ;
        RECT 1906.770 496.780 1907.090 496.840 ;
        RECT 1910.910 496.780 1911.230 496.840 ;
        RECT 1910.910 245.720 1911.230 245.780 ;
        RECT 2704.870 245.720 2705.190 245.780 ;
        RECT 1910.910 245.580 2705.190 245.720 ;
        RECT 1910.910 245.520 1911.230 245.580 ;
        RECT 2704.870 245.520 2705.190 245.580 ;
      LAYER via ;
        RECT 1906.800 496.780 1907.060 497.040 ;
        RECT 1910.940 496.780 1911.200 497.040 ;
        RECT 1910.940 245.520 1911.200 245.780 ;
        RECT 2704.900 245.520 2705.160 245.780 ;
      LAYER met2 ;
        RECT 1906.930 510.340 1907.210 514.000 ;
        RECT 1906.860 510.000 1907.210 510.340 ;
        RECT 1906.860 497.070 1907.000 510.000 ;
        RECT 1906.800 496.750 1907.060 497.070 ;
        RECT 1910.940 496.750 1911.200 497.070 ;
        RECT 1911.000 245.810 1911.140 496.750 ;
        RECT 1910.940 245.490 1911.200 245.810 ;
        RECT 2704.900 245.490 2705.160 245.810 ;
        RECT 2704.960 17.410 2705.100 245.490 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1414.640 2520.730 1414.700 ;
        RECT 2725.570 1414.640 2725.890 1414.700 ;
        RECT 2520.410 1414.500 2725.890 1414.640 ;
        RECT 2520.410 1414.440 2520.730 1414.500 ;
        RECT 2725.570 1414.440 2725.890 1414.500 ;
      LAYER via ;
        RECT 2520.440 1414.440 2520.700 1414.700 ;
        RECT 2725.600 1414.440 2725.860 1414.700 ;
      LAYER met2 ;
        RECT 2520.430 1415.915 2520.710 1416.285 ;
        RECT 2520.500 1414.730 2520.640 1415.915 ;
        RECT 2520.440 1414.410 2520.700 1414.730 ;
        RECT 2725.600 1414.410 2725.860 1414.730 ;
        RECT 2725.660 17.410 2725.800 1414.410 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1415.960 2520.710 1416.240 ;
      LAYER met3 ;
        RECT 2506.000 1416.250 2510.000 1416.400 ;
        RECT 2520.405 1416.250 2520.735 1416.265 ;
        RECT 2506.000 1415.950 2520.735 1416.250 ;
        RECT 2506.000 1415.800 2510.000 1415.950 ;
        RECT 2520.405 1415.935 2520.735 1415.950 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1704.660 2520.730 1704.720 ;
        RECT 2639.090 1704.660 2639.410 1704.720 ;
        RECT 2520.410 1704.520 2639.410 1704.660 ;
        RECT 2520.410 1704.460 2520.730 1704.520 ;
        RECT 2639.090 1704.460 2639.410 1704.520 ;
        RECT 2639.090 24.040 2639.410 24.100 ;
        RECT 2744.430 24.040 2744.750 24.100 ;
        RECT 2639.090 23.900 2744.750 24.040 ;
        RECT 2639.090 23.840 2639.410 23.900 ;
        RECT 2744.430 23.840 2744.750 23.900 ;
      LAYER via ;
        RECT 2520.440 1704.460 2520.700 1704.720 ;
        RECT 2639.120 1704.460 2639.380 1704.720 ;
        RECT 2639.120 23.840 2639.380 24.100 ;
        RECT 2744.460 23.840 2744.720 24.100 ;
      LAYER met2 ;
        RECT 2520.430 1708.315 2520.710 1708.685 ;
        RECT 2520.500 1704.750 2520.640 1708.315 ;
        RECT 2520.440 1704.430 2520.700 1704.750 ;
        RECT 2639.120 1704.430 2639.380 1704.750 ;
        RECT 2639.180 24.130 2639.320 1704.430 ;
        RECT 2639.120 23.810 2639.380 24.130 ;
        RECT 2744.460 23.810 2744.720 24.130 ;
        RECT 2744.520 2.400 2744.660 23.810 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1708.360 2520.710 1708.640 ;
      LAYER met3 ;
        RECT 2506.000 1708.650 2510.000 1708.800 ;
        RECT 2520.405 1708.650 2520.735 1708.665 ;
        RECT 2506.000 1708.350 2520.735 1708.650 ;
        RECT 2506.000 1708.200 2510.000 1708.350 ;
        RECT 2520.405 1708.335 2520.735 1708.350 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 409.010 113.800 409.330 113.860 ;
        RECT 2760.070 113.800 2760.390 113.860 ;
        RECT 409.010 113.660 2760.390 113.800 ;
        RECT 409.010 113.600 409.330 113.660 ;
        RECT 2760.070 113.600 2760.390 113.660 ;
      LAYER via ;
        RECT 409.040 113.600 409.300 113.860 ;
        RECT 2760.100 113.600 2760.360 113.860 ;
      LAYER met2 ;
        RECT 409.030 841.995 409.310 842.365 ;
        RECT 409.100 113.890 409.240 841.995 ;
        RECT 409.040 113.570 409.300 113.890 ;
        RECT 2760.100 113.570 2760.360 113.890 ;
        RECT 2760.160 17.410 2760.300 113.570 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
      LAYER via2 ;
        RECT 409.030 842.040 409.310 842.320 ;
      LAYER met3 ;
        RECT 409.005 842.330 409.335 842.345 ;
        RECT 410.000 842.330 414.000 842.480 ;
        RECT 409.005 842.030 414.000 842.330 ;
        RECT 409.005 842.015 409.335 842.030 ;
        RECT 410.000 841.880 414.000 842.030 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 301.830 2228.940 302.150 2229.000 ;
        RECT 393.370 2228.940 393.690 2229.000 ;
        RECT 301.830 2228.800 393.690 2228.940 ;
        RECT 301.830 2228.740 302.150 2228.800 ;
        RECT 393.370 2228.740 393.690 2228.800 ;
        RECT 301.830 18.940 302.150 19.000 ;
        RECT 835.430 18.940 835.750 19.000 ;
        RECT 301.830 18.800 835.750 18.940 ;
        RECT 301.830 18.740 302.150 18.800 ;
        RECT 835.430 18.740 835.750 18.800 ;
      LAYER via ;
        RECT 301.860 2228.740 302.120 2229.000 ;
        RECT 393.400 2228.740 393.660 2229.000 ;
        RECT 301.860 18.740 302.120 19.000 ;
        RECT 835.460 18.740 835.720 19.000 ;
      LAYER met2 ;
        RECT 393.390 2230.555 393.670 2230.925 ;
        RECT 393.460 2229.030 393.600 2230.555 ;
        RECT 301.860 2228.710 302.120 2229.030 ;
        RECT 393.400 2228.710 393.660 2229.030 ;
        RECT 301.920 19.030 302.060 2228.710 ;
        RECT 301.860 18.710 302.120 19.030 ;
        RECT 835.460 18.710 835.720 19.030 ;
        RECT 835.520 2.400 835.660 18.710 ;
        RECT 835.310 -4.800 835.870 2.400 ;
      LAYER via2 ;
        RECT 393.390 2230.600 393.670 2230.880 ;
      LAYER met3 ;
        RECT 393.365 2230.890 393.695 2230.905 ;
        RECT 410.000 2230.890 414.000 2231.040 ;
        RECT 393.365 2230.590 414.000 2230.890 ;
        RECT 393.365 2230.575 393.695 2230.590 ;
        RECT 410.000 2230.440 414.000 2230.590 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.330 3023.180 1210.650 3023.240 ;
        RECT 2773.870 3023.180 2774.190 3023.240 ;
        RECT 1210.330 3023.040 2774.190 3023.180 ;
        RECT 1210.330 3022.980 1210.650 3023.040 ;
        RECT 2773.870 3022.980 2774.190 3023.040 ;
        RECT 2773.870 17.580 2774.190 17.640 ;
        RECT 2779.850 17.580 2780.170 17.640 ;
        RECT 2773.870 17.440 2780.170 17.580 ;
        RECT 2773.870 17.380 2774.190 17.440 ;
        RECT 2779.850 17.380 2780.170 17.440 ;
      LAYER via ;
        RECT 1210.360 3022.980 1210.620 3023.240 ;
        RECT 2773.900 3022.980 2774.160 3023.240 ;
        RECT 2773.900 17.380 2774.160 17.640 ;
        RECT 2779.880 17.380 2780.140 17.640 ;
      LAYER met2 ;
        RECT 1210.360 3022.950 1210.620 3023.270 ;
        RECT 2773.900 3022.950 2774.160 3023.270 ;
        RECT 1210.420 3010.000 1210.560 3022.950 ;
        RECT 1210.420 3009.340 1210.770 3010.000 ;
        RECT 1210.490 3006.000 1210.770 3009.340 ;
        RECT 2773.960 17.670 2774.100 3022.950 ;
        RECT 2773.900 17.350 2774.160 17.670 ;
        RECT 2779.880 17.350 2780.140 17.670 ;
        RECT 2779.940 2.400 2780.080 17.350 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 691.470 3022.755 691.750 3023.125 ;
        RECT 2794.590 3022.755 2794.870 3023.125 ;
        RECT 691.540 3010.000 691.680 3022.755 ;
        RECT 691.540 3009.340 691.890 3010.000 ;
        RECT 691.610 3006.000 691.890 3009.340 ;
        RECT 2794.660 17.410 2794.800 3022.755 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
      LAYER via2 ;
        RECT 691.470 3022.800 691.750 3023.080 ;
        RECT 2794.590 3022.800 2794.870 3023.080 ;
      LAYER met3 ;
        RECT 691.445 3023.090 691.775 3023.105 ;
        RECT 2794.565 3023.090 2794.895 3023.105 ;
        RECT 691.445 3022.790 2794.895 3023.090 ;
        RECT 691.445 3022.775 691.775 3022.790 ;
        RECT 2794.565 3022.775 2794.895 3022.790 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.290 465.275 2815.570 465.645 ;
        RECT 2815.360 17.410 2815.500 465.275 ;
        RECT 2815.360 17.270 2815.960 17.410 ;
        RECT 2815.820 2.400 2815.960 17.270 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 2815.290 465.320 2815.570 465.600 ;
      LAYER met3 ;
        RECT 405.070 1280.250 405.450 1280.260 ;
        RECT 410.000 1280.250 414.000 1280.400 ;
        RECT 405.070 1279.950 414.000 1280.250 ;
        RECT 405.070 1279.940 405.450 1279.950 ;
        RECT 410.000 1279.800 414.000 1279.950 ;
        RECT 405.070 465.610 405.450 465.620 ;
        RECT 2815.265 465.610 2815.595 465.625 ;
        RECT 405.070 465.310 2815.595 465.610 ;
        RECT 405.070 465.300 405.450 465.310 ;
        RECT 2815.265 465.295 2815.595 465.310 ;
      LAYER via3 ;
        RECT 405.100 1279.940 405.420 1280.260 ;
        RECT 405.100 465.300 405.420 465.620 ;
      LAYER met4 ;
        RECT 405.095 1279.935 405.425 1280.265 ;
        RECT 405.110 465.625 405.410 1279.935 ;
        RECT 405.095 465.295 405.425 465.625 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1117.410 224.300 1117.730 224.360 ;
        RECT 2829.070 224.300 2829.390 224.360 ;
        RECT 1117.410 224.160 2829.390 224.300 ;
        RECT 1117.410 224.100 1117.730 224.160 ;
        RECT 2829.070 224.100 2829.390 224.160 ;
      LAYER via ;
        RECT 1117.440 224.100 1117.700 224.360 ;
        RECT 2829.100 224.100 2829.360 224.360 ;
      LAYER met2 ;
        RECT 1116.650 510.410 1116.930 514.000 ;
        RECT 1116.650 510.270 1117.640 510.410 ;
        RECT 1116.650 510.000 1116.930 510.270 ;
        RECT 1117.500 224.390 1117.640 510.270 ;
        RECT 1117.440 224.070 1117.700 224.390 ;
        RECT 2829.100 224.070 2829.360 224.390 ;
        RECT 2829.160 17.410 2829.300 224.070 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1852.490 3010.600 1852.810 3010.660 ;
        RECT 2849.770 3010.600 2850.090 3010.660 ;
        RECT 1852.490 3010.460 2850.090 3010.600 ;
        RECT 1852.490 3010.400 1852.810 3010.460 ;
        RECT 2849.770 3010.400 2850.090 3010.460 ;
      LAYER via ;
        RECT 1852.520 3010.400 1852.780 3010.660 ;
        RECT 2849.800 3010.400 2850.060 3010.660 ;
      LAYER met2 ;
        RECT 1852.520 3010.370 1852.780 3010.690 ;
        RECT 2849.800 3010.370 2850.060 3010.690 ;
        RECT 1852.580 3010.000 1852.720 3010.370 ;
        RECT 1852.580 3009.340 1852.930 3010.000 ;
        RECT 1852.650 3006.000 1852.930 3009.340 ;
        RECT 2849.860 16.730 2850.000 3010.370 ;
        RECT 2849.860 16.590 2851.380 16.730 ;
        RECT 2851.240 2.400 2851.380 16.590 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1062.740 2520.730 1062.800 ;
        RECT 2701.190 1062.740 2701.510 1062.800 ;
        RECT 2520.410 1062.600 2701.510 1062.740 ;
        RECT 2520.410 1062.540 2520.730 1062.600 ;
        RECT 2701.190 1062.540 2701.510 1062.600 ;
        RECT 2701.190 44.780 2701.510 44.840 ;
        RECT 2869.090 44.780 2869.410 44.840 ;
        RECT 2701.190 44.640 2869.410 44.780 ;
        RECT 2701.190 44.580 2701.510 44.640 ;
        RECT 2869.090 44.580 2869.410 44.640 ;
      LAYER via ;
        RECT 2520.440 1062.540 2520.700 1062.800 ;
        RECT 2701.220 1062.540 2701.480 1062.800 ;
        RECT 2701.220 44.580 2701.480 44.840 ;
        RECT 2869.120 44.580 2869.380 44.840 ;
      LAYER met2 ;
        RECT 2520.430 1069.115 2520.710 1069.485 ;
        RECT 2520.500 1062.830 2520.640 1069.115 ;
        RECT 2520.440 1062.510 2520.700 1062.830 ;
        RECT 2701.220 1062.510 2701.480 1062.830 ;
        RECT 2701.280 44.870 2701.420 1062.510 ;
        RECT 2701.220 44.550 2701.480 44.870 ;
        RECT 2869.120 44.550 2869.380 44.870 ;
        RECT 2869.180 2.400 2869.320 44.550 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1069.160 2520.710 1069.440 ;
      LAYER met3 ;
        RECT 2506.000 1069.450 2510.000 1069.600 ;
        RECT 2520.405 1069.450 2520.735 1069.465 ;
        RECT 2506.000 1069.150 2520.735 1069.450 ;
        RECT 2506.000 1069.000 2510.000 1069.150 ;
        RECT 2520.405 1069.135 2520.735 1069.150 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1489.550 107.340 1489.870 107.400 ;
        RECT 2884.270 107.340 2884.590 107.400 ;
        RECT 1489.550 107.200 2884.590 107.340 ;
        RECT 1489.550 107.140 1489.870 107.200 ;
        RECT 2884.270 107.140 2884.590 107.200 ;
        RECT 2884.270 2.960 2884.590 3.020 ;
        RECT 2887.030 2.960 2887.350 3.020 ;
        RECT 2884.270 2.820 2887.350 2.960 ;
        RECT 2884.270 2.760 2884.590 2.820 ;
        RECT 2887.030 2.760 2887.350 2.820 ;
      LAYER via ;
        RECT 1489.580 107.140 1489.840 107.400 ;
        RECT 2884.300 107.140 2884.560 107.400 ;
        RECT 2884.300 2.760 2884.560 3.020 ;
        RECT 2887.060 2.760 2887.320 3.020 ;
      LAYER met2 ;
        RECT 1487.410 510.410 1487.690 514.000 ;
        RECT 1487.410 510.270 1489.780 510.410 ;
        RECT 1487.410 510.000 1487.690 510.270 ;
        RECT 1489.640 107.430 1489.780 510.270 ;
        RECT 1489.580 107.110 1489.840 107.430 ;
        RECT 2884.300 107.110 2884.560 107.430 ;
        RECT 2884.360 3.050 2884.500 107.110 ;
        RECT 2884.300 2.730 2884.560 3.050 ;
        RECT 2887.060 2.730 2887.320 3.050 ;
        RECT 2887.120 2.400 2887.260 2.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2255.910 169.220 2256.230 169.280 ;
        RECT 2873.690 169.220 2874.010 169.280 ;
        RECT 2255.910 169.080 2874.010 169.220 ;
        RECT 2255.910 169.020 2256.230 169.080 ;
        RECT 2873.690 169.020 2874.010 169.080 ;
        RECT 2873.690 17.720 2874.010 17.980 ;
        RECT 2873.780 17.580 2873.920 17.720 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2873.780 17.440 2905.290 17.580 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
      LAYER via ;
        RECT 2255.940 169.020 2256.200 169.280 ;
        RECT 2873.720 169.020 2873.980 169.280 ;
        RECT 2873.720 17.720 2873.980 17.980 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
      LAYER met2 ;
        RECT 2252.850 510.410 2253.130 514.000 ;
        RECT 2252.850 510.270 2256.140 510.410 ;
        RECT 2252.850 510.000 2253.130 510.270 ;
        RECT 2256.000 169.310 2256.140 510.270 ;
        RECT 2255.940 168.990 2256.200 169.310 ;
        RECT 2873.720 168.990 2873.980 169.310 ;
        RECT 2873.780 18.010 2873.920 168.990 ;
        RECT 2873.720 17.690 2873.980 18.010 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2905.060 2.400 2905.200 17.350 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.570 498.680 609.890 498.740 ;
        RECT 613.710 498.680 614.030 498.740 ;
        RECT 609.570 498.540 614.030 498.680 ;
        RECT 609.570 498.480 609.890 498.540 ;
        RECT 613.710 498.480 614.030 498.540 ;
        RECT 613.710 99.860 614.030 99.920 ;
        RECT 848.770 99.860 849.090 99.920 ;
        RECT 613.710 99.720 849.090 99.860 ;
        RECT 613.710 99.660 614.030 99.720 ;
        RECT 848.770 99.660 849.090 99.720 ;
        RECT 848.770 62.120 849.090 62.180 ;
        RECT 852.910 62.120 853.230 62.180 ;
        RECT 848.770 61.980 853.230 62.120 ;
        RECT 848.770 61.920 849.090 61.980 ;
        RECT 852.910 61.920 853.230 61.980 ;
      LAYER via ;
        RECT 609.600 498.480 609.860 498.740 ;
        RECT 613.740 498.480 614.000 498.740 ;
        RECT 613.740 99.660 614.000 99.920 ;
        RECT 848.800 99.660 849.060 99.920 ;
        RECT 848.800 61.920 849.060 62.180 ;
        RECT 852.940 61.920 853.200 62.180 ;
      LAYER met2 ;
        RECT 609.730 510.340 610.010 514.000 ;
        RECT 609.660 510.000 610.010 510.340 ;
        RECT 609.660 498.770 609.800 510.000 ;
        RECT 609.600 498.450 609.860 498.770 ;
        RECT 613.740 498.450 614.000 498.770 ;
        RECT 613.800 99.950 613.940 498.450 ;
        RECT 613.740 99.630 614.000 99.950 ;
        RECT 848.800 99.630 849.060 99.950 ;
        RECT 848.860 62.210 849.000 99.630 ;
        RECT 848.800 61.890 849.060 62.210 ;
        RECT 852.940 61.890 853.200 62.210 ;
        RECT 853.000 2.400 853.140 61.890 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 371.290 3031.340 371.610 3031.400 ;
        RECT 1617.890 3031.340 1618.210 3031.400 ;
        RECT 371.290 3031.200 1618.210 3031.340 ;
        RECT 371.290 3031.140 371.610 3031.200 ;
        RECT 1617.890 3031.140 1618.210 3031.200 ;
        RECT 370.830 512.960 371.150 513.020 ;
        RECT 869.930 512.960 870.250 513.020 ;
        RECT 370.830 512.820 870.250 512.960 ;
        RECT 370.830 512.760 371.150 512.820 ;
        RECT 869.930 512.760 870.250 512.820 ;
      LAYER via ;
        RECT 371.320 3031.140 371.580 3031.400 ;
        RECT 1617.920 3031.140 1618.180 3031.400 ;
        RECT 370.860 512.760 371.120 513.020 ;
        RECT 869.960 512.760 870.220 513.020 ;
      LAYER met2 ;
        RECT 371.320 3031.110 371.580 3031.430 ;
        RECT 1617.920 3031.110 1618.180 3031.430 ;
        RECT 371.380 538.970 371.520 3031.110 ;
        RECT 1617.980 3010.000 1618.120 3031.110 ;
        RECT 1617.980 3009.340 1618.330 3010.000 ;
        RECT 1618.050 3006.000 1618.330 3009.340 ;
        RECT 370.920 538.830 371.520 538.970 ;
        RECT 370.920 513.050 371.060 538.830 ;
        RECT 370.860 512.730 371.120 513.050 ;
        RECT 869.960 512.730 870.220 513.050 ;
        RECT 870.020 3.130 870.160 512.730 ;
        RECT 870.020 2.990 871.080 3.130 ;
        RECT 870.940 2.400 871.080 2.990 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 883.805 448.205 883.975 482.375 ;
        RECT 883.805 338.045 883.975 385.815 ;
        RECT 883.805 241.485 883.975 289.595 ;
        RECT 883.805 158.525 883.975 193.035 ;
        RECT 884.265 48.365 884.435 96.475 ;
      LAYER mcon ;
        RECT 883.805 482.205 883.975 482.375 ;
        RECT 883.805 385.645 883.975 385.815 ;
        RECT 883.805 289.425 883.975 289.595 ;
        RECT 883.805 192.865 883.975 193.035 ;
        RECT 884.265 96.305 884.435 96.475 ;
      LAYER met1 ;
        RECT 411.310 3025.900 411.630 3025.960 ;
        RECT 1802.810 3025.900 1803.130 3025.960 ;
        RECT 411.310 3025.760 1803.130 3025.900 ;
        RECT 411.310 3025.700 411.630 3025.760 ;
        RECT 1802.810 3025.700 1803.130 3025.760 ;
        RECT 375.890 890.700 376.210 890.760 ;
        RECT 411.310 890.700 411.630 890.760 ;
        RECT 375.890 890.560 411.630 890.700 ;
        RECT 375.890 890.500 376.210 890.560 ;
        RECT 411.310 890.500 411.630 890.560 ;
        RECT 627.510 512.620 627.830 512.680 ;
        RECT 668.450 512.620 668.770 512.680 ;
        RECT 627.510 512.480 668.770 512.620 ;
        RECT 627.510 512.420 627.830 512.480 ;
        RECT 668.450 512.420 668.770 512.480 ;
        RECT 883.730 482.840 884.050 483.100 ;
        RECT 883.820 482.405 883.960 482.840 ;
        RECT 883.745 482.175 884.035 482.405 ;
        RECT 883.730 448.360 884.050 448.420 ;
        RECT 883.535 448.220 884.050 448.360 ;
        RECT 883.730 448.160 884.050 448.220 ;
        RECT 883.270 434.760 883.590 434.820 ;
        RECT 883.730 434.760 884.050 434.820 ;
        RECT 883.270 434.620 884.050 434.760 ;
        RECT 883.270 434.560 883.590 434.620 ;
        RECT 883.730 434.560 884.050 434.620 ;
        RECT 883.745 385.800 884.035 385.845 ;
        RECT 884.190 385.800 884.510 385.860 ;
        RECT 883.745 385.660 884.510 385.800 ;
        RECT 883.745 385.615 884.035 385.660 ;
        RECT 884.190 385.600 884.510 385.660 ;
        RECT 883.730 338.200 884.050 338.260 ;
        RECT 883.535 338.060 884.050 338.200 ;
        RECT 883.730 338.000 884.050 338.060 ;
        RECT 883.745 289.580 884.035 289.625 ;
        RECT 884.190 289.580 884.510 289.640 ;
        RECT 883.745 289.440 884.510 289.580 ;
        RECT 883.745 289.395 884.035 289.440 ;
        RECT 884.190 289.380 884.510 289.440 ;
        RECT 883.730 241.640 884.050 241.700 ;
        RECT 883.535 241.500 884.050 241.640 ;
        RECT 883.730 241.440 884.050 241.500 ;
        RECT 883.745 193.020 884.035 193.065 ;
        RECT 884.190 193.020 884.510 193.080 ;
        RECT 883.745 192.880 884.510 193.020 ;
        RECT 883.745 192.835 884.035 192.880 ;
        RECT 884.190 192.820 884.510 192.880 ;
        RECT 883.730 158.680 884.050 158.740 ;
        RECT 883.535 158.540 884.050 158.680 ;
        RECT 883.730 158.480 884.050 158.540 ;
        RECT 884.190 96.460 884.510 96.520 ;
        RECT 883.995 96.320 884.510 96.460 ;
        RECT 884.190 96.260 884.510 96.320 ;
        RECT 884.205 48.520 884.495 48.565 ;
        RECT 884.650 48.520 884.970 48.580 ;
        RECT 884.205 48.380 884.970 48.520 ;
        RECT 884.205 48.335 884.495 48.380 ;
        RECT 884.650 48.320 884.970 48.380 ;
        RECT 884.650 20.300 884.970 20.360 ;
        RECT 888.790 20.300 889.110 20.360 ;
        RECT 884.650 20.160 889.110 20.300 ;
        RECT 884.650 20.100 884.970 20.160 ;
        RECT 888.790 20.100 889.110 20.160 ;
      LAYER via ;
        RECT 411.340 3025.700 411.600 3025.960 ;
        RECT 1802.840 3025.700 1803.100 3025.960 ;
        RECT 375.920 890.500 376.180 890.760 ;
        RECT 411.340 890.500 411.600 890.760 ;
        RECT 627.540 512.420 627.800 512.680 ;
        RECT 668.480 512.420 668.740 512.680 ;
        RECT 883.760 482.840 884.020 483.100 ;
        RECT 883.760 448.160 884.020 448.420 ;
        RECT 883.300 434.560 883.560 434.820 ;
        RECT 883.760 434.560 884.020 434.820 ;
        RECT 884.220 385.600 884.480 385.860 ;
        RECT 883.760 338.000 884.020 338.260 ;
        RECT 884.220 289.380 884.480 289.640 ;
        RECT 883.760 241.440 884.020 241.700 ;
        RECT 884.220 192.820 884.480 193.080 ;
        RECT 883.760 158.480 884.020 158.740 ;
        RECT 884.220 96.260 884.480 96.520 ;
        RECT 884.680 48.320 884.940 48.580 ;
        RECT 884.680 20.100 884.940 20.360 ;
        RECT 888.820 20.100 889.080 20.360 ;
      LAYER met2 ;
        RECT 411.340 3025.670 411.600 3025.990 ;
        RECT 1802.840 3025.670 1803.100 3025.990 ;
        RECT 411.400 890.790 411.540 3025.670 ;
        RECT 1802.900 3010.000 1803.040 3025.670 ;
        RECT 1802.900 3009.340 1803.250 3010.000 ;
        RECT 1802.970 3006.000 1803.250 3009.340 ;
        RECT 375.920 890.470 376.180 890.790 ;
        RECT 411.340 890.470 411.600 890.790 ;
        RECT 375.980 513.925 376.120 890.470 ;
        RECT 375.910 513.555 376.190 513.925 ;
        RECT 669.460 513.670 670.060 513.810 ;
        RECT 669.460 513.245 669.600 513.670 ;
        RECT 544.730 513.130 545.010 513.245 ;
        RECT 545.650 513.130 545.930 513.245 ;
        RECT 544.730 512.990 545.930 513.130 ;
        RECT 544.730 512.875 545.010 512.990 ;
        RECT 545.650 512.875 545.930 512.990 ;
        RECT 592.110 513.130 592.390 513.245 ;
        RECT 593.030 513.130 593.310 513.245 ;
        RECT 592.110 512.990 593.310 513.130 ;
        RECT 592.110 512.875 592.390 512.990 ;
        RECT 593.030 512.875 593.310 512.990 ;
        RECT 627.530 512.875 627.810 513.245 ;
        RECT 668.470 512.875 668.750 513.245 ;
        RECT 669.390 512.875 669.670 513.245 ;
        RECT 627.600 512.710 627.740 512.875 ;
        RECT 668.540 512.710 668.680 512.875 ;
        RECT 627.540 512.390 627.800 512.710 ;
        RECT 668.480 512.390 668.740 512.710 ;
        RECT 669.920 512.565 670.060 513.670 ;
        RECT 883.750 513.130 884.030 513.245 ;
        RECT 883.360 512.990 884.030 513.130 ;
        RECT 669.850 512.195 670.130 512.565 ;
        RECT 883.360 496.810 883.500 512.990 ;
        RECT 883.750 512.875 884.030 512.990 ;
        RECT 883.360 496.670 883.960 496.810 ;
        RECT 883.820 483.130 883.960 496.670 ;
        RECT 883.760 482.810 884.020 483.130 ;
        RECT 883.760 448.130 884.020 448.450 ;
        RECT 883.820 434.930 883.960 448.130 ;
        RECT 883.360 434.850 883.960 434.930 ;
        RECT 883.300 434.790 884.020 434.850 ;
        RECT 883.300 434.530 883.560 434.790 ;
        RECT 883.760 434.530 884.020 434.790 ;
        RECT 883.820 399.570 883.960 434.530 ;
        RECT 883.820 399.430 884.420 399.570 ;
        RECT 884.280 385.890 884.420 399.430 ;
        RECT 884.220 385.570 884.480 385.890 ;
        RECT 883.760 337.970 884.020 338.290 ;
        RECT 883.820 303.690 883.960 337.970 ;
        RECT 883.820 303.550 884.420 303.690 ;
        RECT 884.280 289.670 884.420 303.550 ;
        RECT 884.220 289.350 884.480 289.670 ;
        RECT 883.760 241.410 884.020 241.730 ;
        RECT 883.820 207.130 883.960 241.410 ;
        RECT 883.820 206.990 884.420 207.130 ;
        RECT 884.280 193.110 884.420 206.990 ;
        RECT 884.220 192.790 884.480 193.110 ;
        RECT 883.760 158.450 884.020 158.770 ;
        RECT 883.820 110.570 883.960 158.450 ;
        RECT 883.820 110.430 884.420 110.570 ;
        RECT 884.280 96.550 884.420 110.430 ;
        RECT 884.220 96.230 884.480 96.550 ;
        RECT 884.680 48.290 884.940 48.610 ;
        RECT 884.740 20.390 884.880 48.290 ;
        RECT 884.680 20.070 884.940 20.390 ;
        RECT 888.820 20.070 889.080 20.390 ;
        RECT 888.880 2.400 889.020 20.070 ;
        RECT 888.670 -4.800 889.230 2.400 ;
      LAYER via2 ;
        RECT 375.910 513.600 376.190 513.880 ;
        RECT 544.730 512.920 545.010 513.200 ;
        RECT 545.650 512.920 545.930 513.200 ;
        RECT 592.110 512.920 592.390 513.200 ;
        RECT 593.030 512.920 593.310 513.200 ;
        RECT 627.530 512.920 627.810 513.200 ;
        RECT 668.470 512.920 668.750 513.200 ;
        RECT 669.390 512.920 669.670 513.200 ;
        RECT 669.850 512.240 670.130 512.520 ;
        RECT 883.750 512.920 884.030 513.200 ;
      LAYER met3 ;
        RECT 375.885 513.890 376.215 513.905 ;
        RECT 375.885 513.590 541.570 513.890 ;
        RECT 375.885 513.575 376.215 513.590 ;
        RECT 541.270 513.210 541.570 513.590 ;
        RECT 593.710 513.590 621.610 513.890 ;
        RECT 544.705 513.210 545.035 513.225 ;
        RECT 541.270 512.910 545.035 513.210 ;
        RECT 544.705 512.895 545.035 512.910 ;
        RECT 545.625 513.210 545.955 513.225 ;
        RECT 592.085 513.210 592.415 513.225 ;
        RECT 545.625 512.910 592.415 513.210 ;
        RECT 545.625 512.895 545.955 512.910 ;
        RECT 592.085 512.895 592.415 512.910 ;
        RECT 593.005 513.210 593.335 513.225 ;
        RECT 593.710 513.210 594.010 513.590 ;
        RECT 593.005 512.910 594.010 513.210 ;
        RECT 621.310 513.210 621.610 513.590 ;
        RECT 693.070 513.590 724.650 513.890 ;
        RECT 627.505 513.210 627.835 513.225 ;
        RECT 621.310 512.910 627.835 513.210 ;
        RECT 593.005 512.895 593.335 512.910 ;
        RECT 627.505 512.895 627.835 512.910 ;
        RECT 668.445 513.210 668.775 513.225 ;
        RECT 669.365 513.210 669.695 513.225 ;
        RECT 668.445 512.910 669.695 513.210 ;
        RECT 668.445 512.895 668.775 512.910 ;
        RECT 669.365 512.895 669.695 512.910 ;
        RECT 669.825 512.530 670.155 512.545 ;
        RECT 693.070 512.530 693.370 513.590 ;
        RECT 724.350 513.220 724.650 513.590 ;
        RECT 773.110 513.590 834.130 513.890 ;
        RECT 724.310 512.900 724.690 513.220 ;
        RECT 773.110 513.210 773.410 513.590 ;
        RECT 772.190 512.910 773.410 513.210 ;
        RECT 833.830 513.040 834.130 513.590 ;
        RECT 883.725 513.210 884.055 513.225 ;
        RECT 835.670 513.040 884.055 513.210 ;
        RECT 833.830 512.910 884.055 513.040 ;
        RECT 669.825 512.230 693.370 512.530 ;
        RECT 669.825 512.215 670.155 512.230 ;
        RECT 724.310 511.850 724.690 511.860 ;
        RECT 772.190 511.850 772.490 512.910 ;
        RECT 833.830 512.740 835.970 512.910 ;
        RECT 883.725 512.895 884.055 512.910 ;
        RECT 724.310 511.550 772.490 511.850 ;
        RECT 724.310 511.540 724.690 511.550 ;
      LAYER via3 ;
        RECT 724.340 512.900 724.660 513.220 ;
        RECT 724.340 511.540 724.660 511.860 ;
      LAYER met4 ;
        RECT 724.335 512.895 724.665 513.225 ;
        RECT 724.350 511.865 724.650 512.895 ;
        RECT 724.335 511.535 724.665 511.865 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.410 162.760 910.730 162.820 ;
        RECT 1262.770 162.760 1263.090 162.820 ;
        RECT 910.410 162.620 1263.090 162.760 ;
        RECT 910.410 162.560 910.730 162.620 ;
        RECT 1262.770 162.560 1263.090 162.620 ;
        RECT 906.730 14.860 907.050 14.920 ;
        RECT 910.410 14.860 910.730 14.920 ;
        RECT 906.730 14.720 910.730 14.860 ;
        RECT 906.730 14.660 907.050 14.720 ;
        RECT 910.410 14.660 910.730 14.720 ;
      LAYER via ;
        RECT 910.440 162.560 910.700 162.820 ;
        RECT 1262.800 162.560 1263.060 162.820 ;
        RECT 906.760 14.660 907.020 14.920 ;
        RECT 910.440 14.660 910.700 14.920 ;
      LAYER met2 ;
        RECT 1264.770 510.410 1265.050 514.000 ;
        RECT 1262.860 510.270 1265.050 510.410 ;
        RECT 1262.860 162.850 1263.000 510.270 ;
        RECT 1264.770 510.000 1265.050 510.270 ;
        RECT 910.440 162.530 910.700 162.850 ;
        RECT 1262.800 162.530 1263.060 162.850 ;
        RECT 910.500 14.950 910.640 162.530 ;
        RECT 906.760 14.630 907.020 14.950 ;
        RECT 910.440 14.630 910.700 14.950 ;
        RECT 906.820 2.400 906.960 14.630 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 148.480 924.530 148.540 ;
        RECT 2421.970 148.480 2422.290 148.540 ;
        RECT 924.210 148.340 2422.290 148.480 ;
        RECT 924.210 148.280 924.530 148.340 ;
        RECT 2421.970 148.280 2422.290 148.340 ;
      LAYER via ;
        RECT 924.240 148.280 924.500 148.540 ;
        RECT 2422.000 148.280 2422.260 148.540 ;
      LAYER met2 ;
        RECT 2425.810 510.410 2426.090 514.000 ;
        RECT 2422.060 510.270 2426.090 510.410 ;
        RECT 2422.060 148.570 2422.200 510.270 ;
        RECT 2425.810 510.000 2426.090 510.270 ;
        RECT 924.240 148.250 924.500 148.570 ;
        RECT 2422.000 148.250 2422.260 148.570 ;
        RECT 924.300 2.400 924.440 148.250 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 917.845 509.065 918.015 512.975 ;
      LAYER mcon ;
        RECT 917.845 512.805 918.015 512.975 ;
      LAYER met1 ;
        RECT 364.850 3026.240 365.170 3026.300 ;
        RECT 962.850 3026.240 963.170 3026.300 ;
        RECT 364.850 3026.100 963.170 3026.240 ;
        RECT 364.850 3026.040 365.170 3026.100 ;
        RECT 962.850 3026.040 963.170 3026.100 ;
        RECT 364.850 513.300 365.170 513.360 ;
        RECT 364.850 513.160 918.000 513.300 ;
        RECT 364.850 513.100 365.170 513.160 ;
        RECT 917.860 513.005 918.000 513.160 ;
        RECT 917.785 512.775 918.075 513.005 ;
        RECT 917.785 509.220 918.075 509.265 ;
        RECT 938.930 509.220 939.250 509.280 ;
        RECT 917.785 509.080 939.250 509.220 ;
        RECT 917.785 509.035 918.075 509.080 ;
        RECT 938.930 509.020 939.250 509.080 ;
        RECT 938.930 16.900 939.250 16.960 ;
        RECT 942.150 16.900 942.470 16.960 ;
        RECT 938.930 16.760 942.470 16.900 ;
        RECT 938.930 16.700 939.250 16.760 ;
        RECT 942.150 16.700 942.470 16.760 ;
      LAYER via ;
        RECT 364.880 3026.040 365.140 3026.300 ;
        RECT 962.880 3026.040 963.140 3026.300 ;
        RECT 364.880 513.100 365.140 513.360 ;
        RECT 938.960 509.020 939.220 509.280 ;
        RECT 938.960 16.700 939.220 16.960 ;
        RECT 942.180 16.700 942.440 16.960 ;
      LAYER met2 ;
        RECT 364.880 3026.010 365.140 3026.330 ;
        RECT 962.880 3026.010 963.140 3026.330 ;
        RECT 364.940 513.390 365.080 3026.010 ;
        RECT 962.940 3010.000 963.080 3026.010 ;
        RECT 962.940 3009.340 963.290 3010.000 ;
        RECT 963.010 3006.000 963.290 3009.340 ;
        RECT 364.880 513.070 365.140 513.390 ;
        RECT 938.960 508.990 939.220 509.310 ;
        RECT 939.020 16.990 939.160 508.990 ;
        RECT 938.960 16.670 939.220 16.990 ;
        RECT 942.180 16.670 942.440 16.990 ;
        RECT 942.240 2.400 942.380 16.670 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 965.610 80.140 965.930 80.200 ;
        RECT 1987.270 80.140 1987.590 80.200 ;
        RECT 965.610 80.000 1987.590 80.140 ;
        RECT 965.610 79.940 965.930 80.000 ;
        RECT 1987.270 79.940 1987.590 80.000 ;
        RECT 960.090 16.900 960.410 16.960 ;
        RECT 965.610 16.900 965.930 16.960 ;
        RECT 960.090 16.760 965.930 16.900 ;
        RECT 960.090 16.700 960.410 16.760 ;
        RECT 965.610 16.700 965.930 16.760 ;
      LAYER via ;
        RECT 965.640 79.940 965.900 80.200 ;
        RECT 1987.300 79.940 1987.560 80.200 ;
        RECT 960.120 16.700 960.380 16.960 ;
        RECT 965.640 16.700 965.900 16.960 ;
      LAYER met2 ;
        RECT 1993.410 510.410 1993.690 514.000 ;
        RECT 1987.360 510.270 1993.690 510.410 ;
        RECT 1987.360 80.230 1987.500 510.270 ;
        RECT 1993.410 510.000 1993.690 510.270 ;
        RECT 965.640 79.910 965.900 80.230 ;
        RECT 1987.300 79.910 1987.560 80.230 ;
        RECT 965.700 16.990 965.840 79.910 ;
        RECT 960.120 16.670 960.380 16.990 ;
        RECT 965.640 16.670 965.900 16.990 ;
        RECT 960.180 2.400 960.320 16.670 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2380.580 2519.810 2380.640 ;
        RECT 2582.510 2380.580 2582.830 2380.640 ;
        RECT 2519.490 2380.440 2582.830 2380.580 ;
        RECT 2519.490 2380.380 2519.810 2380.440 ;
        RECT 2582.510 2380.380 2582.830 2380.440 ;
        RECT 979.410 479.980 979.730 480.040 ;
        RECT 2582.510 479.980 2582.830 480.040 ;
        RECT 979.410 479.840 2582.830 479.980 ;
        RECT 979.410 479.780 979.730 479.840 ;
        RECT 2582.510 479.780 2582.830 479.840 ;
      LAYER via ;
        RECT 2519.520 2380.380 2519.780 2380.640 ;
        RECT 2582.540 2380.380 2582.800 2380.640 ;
        RECT 979.440 479.780 979.700 480.040 ;
        RECT 2582.540 479.780 2582.800 480.040 ;
      LAYER met2 ;
        RECT 2519.510 2384.235 2519.790 2384.605 ;
        RECT 2519.580 2380.670 2519.720 2384.235 ;
        RECT 2519.520 2380.350 2519.780 2380.670 ;
        RECT 2582.540 2380.350 2582.800 2380.670 ;
        RECT 2582.600 480.070 2582.740 2380.350 ;
        RECT 979.440 479.750 979.700 480.070 ;
        RECT 2582.540 479.750 2582.800 480.070 ;
        RECT 979.500 17.410 979.640 479.750 ;
        RECT 978.120 17.270 979.640 17.410 ;
        RECT 978.120 2.400 978.260 17.270 ;
        RECT 977.910 -4.800 978.470 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2384.280 2519.790 2384.560 ;
      LAYER met3 ;
        RECT 2506.000 2384.570 2510.000 2384.720 ;
        RECT 2519.485 2384.570 2519.815 2384.585 ;
        RECT 2506.000 2384.270 2519.815 2384.570 ;
        RECT 2506.000 2384.120 2510.000 2384.270 ;
        RECT 2519.485 2384.255 2519.815 2384.270 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1455.970 3006.320 1456.290 3006.580 ;
        RECT 364.390 3003.800 364.710 3003.860 ;
        RECT 1456.060 3003.800 1456.200 3006.320 ;
        RECT 364.390 3003.660 1456.200 3003.800 ;
        RECT 364.390 3003.600 364.710 3003.660 ;
      LAYER via ;
        RECT 1456.000 3006.320 1456.260 3006.580 ;
        RECT 364.420 3003.600 364.680 3003.860 ;
      LAYER met2 ;
        RECT 1457.050 3006.690 1457.330 3010.000 ;
        RECT 1456.060 3006.610 1457.330 3006.690 ;
        RECT 1456.000 3006.550 1457.330 3006.610 ;
        RECT 1456.000 3006.290 1456.260 3006.550 ;
        RECT 1457.050 3006.000 1457.330 3006.550 ;
        RECT 364.420 3003.570 364.680 3003.890 ;
        RECT 364.480 507.125 364.620 3003.570 ;
        RECT 364.410 506.755 364.690 507.125 ;
        RECT 656.050 506.755 656.330 507.125 ;
        RECT 656.120 17.410 656.260 506.755 ;
        RECT 656.120 17.270 657.180 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 364.410 506.800 364.690 507.080 ;
        RECT 656.050 506.800 656.330 507.080 ;
      LAYER met3 ;
        RECT 364.385 507.090 364.715 507.105 ;
        RECT 656.025 507.090 656.355 507.105 ;
        RECT 364.385 506.790 656.355 507.090 ;
        RECT 364.385 506.775 364.715 506.790 ;
        RECT 656.025 506.775 656.355 506.790 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2601.580 2519.810 2601.640 ;
        RECT 2603.670 2601.580 2603.990 2601.640 ;
        RECT 2519.490 2601.440 2603.990 2601.580 ;
        RECT 2519.490 2601.380 2519.810 2601.440 ;
        RECT 2603.670 2601.380 2603.990 2601.440 ;
        RECT 1000.110 466.720 1000.430 466.780 ;
        RECT 2603.670 466.720 2603.990 466.780 ;
        RECT 1000.110 466.580 2603.990 466.720 ;
        RECT 1000.110 466.520 1000.430 466.580 ;
        RECT 2603.670 466.520 2603.990 466.580 ;
        RECT 995.970 20.300 996.290 20.360 ;
        RECT 1000.110 20.300 1000.430 20.360 ;
        RECT 995.970 20.160 1000.430 20.300 ;
        RECT 995.970 20.100 996.290 20.160 ;
        RECT 1000.110 20.100 1000.430 20.160 ;
      LAYER via ;
        RECT 2519.520 2601.380 2519.780 2601.640 ;
        RECT 2603.700 2601.380 2603.960 2601.640 ;
        RECT 1000.140 466.520 1000.400 466.780 ;
        RECT 2603.700 466.520 2603.960 466.780 ;
        RECT 996.000 20.100 996.260 20.360 ;
        RECT 1000.140 20.100 1000.400 20.360 ;
      LAYER met2 ;
        RECT 2519.510 2603.195 2519.790 2603.565 ;
        RECT 2519.580 2601.670 2519.720 2603.195 ;
        RECT 2519.520 2601.350 2519.780 2601.670 ;
        RECT 2603.700 2601.350 2603.960 2601.670 ;
        RECT 2603.760 466.810 2603.900 2601.350 ;
        RECT 1000.140 466.490 1000.400 466.810 ;
        RECT 2603.700 466.490 2603.960 466.810 ;
        RECT 1000.200 20.390 1000.340 466.490 ;
        RECT 996.000 20.070 996.260 20.390 ;
        RECT 1000.140 20.070 1000.400 20.390 ;
        RECT 996.060 2.400 996.200 20.070 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2603.240 2519.790 2603.520 ;
      LAYER met3 ;
        RECT 2506.000 2603.530 2510.000 2603.680 ;
        RECT 2519.485 2603.530 2519.815 2603.545 ;
        RECT 2506.000 2603.230 2519.815 2603.530 ;
        RECT 2506.000 2603.080 2510.000 2603.230 ;
        RECT 2519.485 2603.215 2519.815 2603.230 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 489.585 3004.665 489.755 3006.535 ;
        RECT 917.845 513.315 918.015 513.655 ;
        RECT 917.845 513.145 918.475 513.315 ;
      LAYER mcon ;
        RECT 489.585 3006.365 489.755 3006.535 ;
        RECT 917.845 513.485 918.015 513.655 ;
        RECT 918.305 513.145 918.475 513.315 ;
      LAYER met1 ;
        RECT 489.510 3017.400 489.830 3017.460 ;
        RECT 987.690 3017.400 988.010 3017.460 ;
        RECT 489.510 3017.260 988.010 3017.400 ;
        RECT 489.510 3017.200 489.830 3017.260 ;
        RECT 987.690 3017.200 988.010 3017.260 ;
        RECT 489.510 3006.520 489.830 3006.580 ;
        RECT 489.315 3006.380 489.830 3006.520 ;
        RECT 489.510 3006.320 489.830 3006.380 ;
        RECT 405.330 3004.820 405.650 3004.880 ;
        RECT 489.525 3004.820 489.815 3004.865 ;
        RECT 405.330 3004.680 489.815 3004.820 ;
        RECT 405.330 3004.620 405.650 3004.680 ;
        RECT 489.525 3004.635 489.815 3004.680 ;
        RECT 405.330 896.820 405.650 896.880 ;
        RECT 409.470 896.820 409.790 896.880 ;
        RECT 405.330 896.680 409.790 896.820 ;
        RECT 405.330 896.620 405.650 896.680 ;
        RECT 409.470 896.620 409.790 896.680 ;
        RECT 405.330 600.340 405.650 600.400 ;
        RECT 409.470 600.340 409.790 600.400 ;
        RECT 405.330 600.200 409.790 600.340 ;
        RECT 405.330 600.140 405.650 600.200 ;
        RECT 409.470 600.140 409.790 600.200 ;
        RECT 405.330 513.640 405.650 513.700 ;
        RECT 917.785 513.640 918.075 513.685 ;
        RECT 1007.470 513.640 1007.790 513.700 ;
        RECT 405.330 513.500 918.075 513.640 ;
        RECT 405.330 513.440 405.650 513.500 ;
        RECT 917.785 513.455 918.075 513.500 ;
        RECT 919.240 513.500 1007.790 513.640 ;
        RECT 918.245 513.300 918.535 513.345 ;
        RECT 919.240 513.300 919.380 513.500 ;
        RECT 1007.470 513.440 1007.790 513.500 ;
        RECT 918.245 513.160 919.380 513.300 ;
        RECT 918.245 513.115 918.535 513.160 ;
        RECT 1007.470 37.640 1007.790 37.700 ;
        RECT 1013.450 37.640 1013.770 37.700 ;
        RECT 1007.470 37.500 1013.770 37.640 ;
        RECT 1007.470 37.440 1007.790 37.500 ;
        RECT 1013.450 37.440 1013.770 37.500 ;
      LAYER via ;
        RECT 489.540 3017.200 489.800 3017.460 ;
        RECT 987.720 3017.200 987.980 3017.460 ;
        RECT 489.540 3006.320 489.800 3006.580 ;
        RECT 405.360 3004.620 405.620 3004.880 ;
        RECT 405.360 896.620 405.620 896.880 ;
        RECT 409.500 896.620 409.760 896.880 ;
        RECT 405.360 600.140 405.620 600.400 ;
        RECT 409.500 600.140 409.760 600.400 ;
        RECT 405.360 513.440 405.620 513.700 ;
        RECT 1007.500 513.440 1007.760 513.700 ;
        RECT 1007.500 37.440 1007.760 37.700 ;
        RECT 1013.480 37.440 1013.740 37.700 ;
      LAYER met2 ;
        RECT 489.540 3017.170 489.800 3017.490 ;
        RECT 987.720 3017.170 987.980 3017.490 ;
        RECT 489.600 3006.610 489.740 3017.170 ;
        RECT 987.780 3010.000 987.920 3017.170 ;
        RECT 987.780 3009.340 988.130 3010.000 ;
        RECT 489.540 3006.290 489.800 3006.610 ;
        RECT 987.850 3006.000 988.130 3009.340 ;
        RECT 405.360 3004.590 405.620 3004.910 ;
        RECT 405.420 896.910 405.560 3004.590 ;
        RECT 405.360 896.590 405.620 896.910 ;
        RECT 409.500 896.590 409.760 896.910 ;
        RECT 409.560 600.430 409.700 896.590 ;
        RECT 405.360 600.110 405.620 600.430 ;
        RECT 409.500 600.110 409.760 600.430 ;
        RECT 405.420 513.730 405.560 600.110 ;
        RECT 405.360 513.410 405.620 513.730 ;
        RECT 1007.500 513.410 1007.760 513.730 ;
        RECT 1007.560 37.730 1007.700 513.410 ;
        RECT 1007.500 37.410 1007.760 37.730 ;
        RECT 1013.480 37.410 1013.740 37.730 ;
        RECT 1013.540 2.400 1013.680 37.410 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.390 2153.120 295.710 2153.180 ;
        RECT 393.370 2153.120 393.690 2153.180 ;
        RECT 295.390 2152.980 393.690 2153.120 ;
        RECT 295.390 2152.920 295.710 2152.980 ;
        RECT 393.370 2152.920 393.690 2152.980 ;
        RECT 295.390 47.500 295.710 47.560 ;
        RECT 1031.390 47.500 1031.710 47.560 ;
        RECT 295.390 47.360 1031.710 47.500 ;
        RECT 295.390 47.300 295.710 47.360 ;
        RECT 1031.390 47.300 1031.710 47.360 ;
      LAYER via ;
        RECT 295.420 2152.920 295.680 2153.180 ;
        RECT 393.400 2152.920 393.660 2153.180 ;
        RECT 295.420 47.300 295.680 47.560 ;
        RECT 1031.420 47.300 1031.680 47.560 ;
      LAYER met2 ;
        RECT 393.390 2157.115 393.670 2157.485 ;
        RECT 393.460 2153.210 393.600 2157.115 ;
        RECT 295.420 2152.890 295.680 2153.210 ;
        RECT 393.400 2152.890 393.660 2153.210 ;
        RECT 295.480 47.590 295.620 2152.890 ;
        RECT 295.420 47.270 295.680 47.590 ;
        RECT 1031.420 47.270 1031.680 47.590 ;
        RECT 1031.480 2.400 1031.620 47.270 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 393.390 2157.160 393.670 2157.440 ;
      LAYER met3 ;
        RECT 393.365 2157.450 393.695 2157.465 ;
        RECT 410.000 2157.450 414.000 2157.600 ;
        RECT 393.365 2157.150 414.000 2157.450 ;
        RECT 393.365 2157.135 393.695 2157.150 ;
        RECT 410.000 2157.000 414.000 2157.150 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1054.390 417.760 1054.710 417.820 ;
        RECT 2513.510 417.760 2513.830 417.820 ;
        RECT 1054.390 417.620 2513.830 417.760 ;
        RECT 1054.390 417.560 1054.710 417.620 ;
        RECT 2513.510 417.560 2513.830 417.620 ;
        RECT 1049.330 20.300 1049.650 20.360 ;
        RECT 1054.390 20.300 1054.710 20.360 ;
        RECT 1049.330 20.160 1054.710 20.300 ;
        RECT 1049.330 20.100 1049.650 20.160 ;
        RECT 1054.390 20.100 1054.710 20.160 ;
      LAYER via ;
        RECT 1054.420 417.560 1054.680 417.820 ;
        RECT 2513.540 417.560 2513.800 417.820 ;
        RECT 1049.360 20.100 1049.620 20.360 ;
        RECT 1054.420 20.100 1054.680 20.360 ;
      LAYER met2 ;
        RECT 2513.530 1324.795 2513.810 1325.165 ;
        RECT 2513.600 417.850 2513.740 1324.795 ;
        RECT 1054.420 417.530 1054.680 417.850 ;
        RECT 2513.540 417.530 2513.800 417.850 ;
        RECT 1054.480 20.390 1054.620 417.530 ;
        RECT 1049.360 20.070 1049.620 20.390 ;
        RECT 1054.420 20.070 1054.680 20.390 ;
        RECT 1049.420 2.400 1049.560 20.070 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 2513.530 1324.840 2513.810 1325.120 ;
      LAYER met3 ;
        RECT 2506.000 1325.130 2510.000 1325.280 ;
        RECT 2513.505 1325.130 2513.835 1325.145 ;
        RECT 2506.000 1324.830 2513.835 1325.130 ;
        RECT 2506.000 1324.680 2510.000 1324.830 ;
        RECT 2513.505 1324.815 2513.835 1324.830 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 398.890 486.440 399.210 486.500 ;
        RECT 1062.670 486.440 1062.990 486.500 ;
        RECT 398.890 486.300 1062.990 486.440 ;
        RECT 398.890 486.240 399.210 486.300 ;
        RECT 1062.670 486.240 1062.990 486.300 ;
        RECT 1062.670 62.120 1062.990 62.180 ;
        RECT 1067.270 62.120 1067.590 62.180 ;
        RECT 1062.670 61.980 1067.590 62.120 ;
        RECT 1062.670 61.920 1062.990 61.980 ;
        RECT 1067.270 61.920 1067.590 61.980 ;
      LAYER via ;
        RECT 398.920 486.240 399.180 486.500 ;
        RECT 1062.700 486.240 1062.960 486.500 ;
        RECT 1062.700 61.920 1062.960 62.180 ;
        RECT 1067.300 61.920 1067.560 62.180 ;
      LAYER met2 ;
        RECT 398.910 1719.195 399.190 1719.565 ;
        RECT 398.980 486.530 399.120 1719.195 ;
        RECT 398.920 486.210 399.180 486.530 ;
        RECT 1062.700 486.210 1062.960 486.530 ;
        RECT 1062.760 62.210 1062.900 486.210 ;
        RECT 1062.700 61.890 1062.960 62.210 ;
        RECT 1067.300 61.890 1067.560 62.210 ;
        RECT 1067.360 2.400 1067.500 61.890 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 398.910 1719.240 399.190 1719.520 ;
      LAYER met3 ;
        RECT 398.885 1719.530 399.215 1719.545 ;
        RECT 410.000 1719.530 414.000 1719.680 ;
        RECT 398.885 1719.230 414.000 1719.530 ;
        RECT 398.885 1719.215 399.215 1719.230 ;
        RECT 410.000 1719.080 414.000 1719.230 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2691.340 2519.810 2691.400 ;
        RECT 2609.650 2691.340 2609.970 2691.400 ;
        RECT 2519.490 2691.200 2609.970 2691.340 ;
        RECT 2519.490 2691.140 2519.810 2691.200 ;
        RECT 2609.650 2691.140 2609.970 2691.200 ;
        RECT 1089.810 467.060 1090.130 467.120 ;
        RECT 2609.650 467.060 2609.970 467.120 ;
        RECT 1089.810 466.920 2609.970 467.060 ;
        RECT 1089.810 466.860 1090.130 466.920 ;
        RECT 2609.650 466.860 2609.970 466.920 ;
        RECT 1085.210 20.300 1085.530 20.360 ;
        RECT 1089.810 20.300 1090.130 20.360 ;
        RECT 1085.210 20.160 1090.130 20.300 ;
        RECT 1085.210 20.100 1085.530 20.160 ;
        RECT 1089.810 20.100 1090.130 20.160 ;
      LAYER via ;
        RECT 2519.520 2691.140 2519.780 2691.400 ;
        RECT 2609.680 2691.140 2609.940 2691.400 ;
        RECT 1089.840 466.860 1090.100 467.120 ;
        RECT 2609.680 466.860 2609.940 467.120 ;
        RECT 1085.240 20.100 1085.500 20.360 ;
        RECT 1089.840 20.100 1090.100 20.360 ;
      LAYER met2 ;
        RECT 2519.510 2694.315 2519.790 2694.685 ;
        RECT 2519.580 2691.430 2519.720 2694.315 ;
        RECT 2519.520 2691.110 2519.780 2691.430 ;
        RECT 2609.680 2691.110 2609.940 2691.430 ;
        RECT 2609.740 467.150 2609.880 2691.110 ;
        RECT 1089.840 466.830 1090.100 467.150 ;
        RECT 2609.680 466.830 2609.940 467.150 ;
        RECT 1089.900 20.390 1090.040 466.830 ;
        RECT 1085.240 20.070 1085.500 20.390 ;
        RECT 1089.840 20.070 1090.100 20.390 ;
        RECT 1085.300 2.400 1085.440 20.070 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2694.360 2519.790 2694.640 ;
      LAYER met3 ;
        RECT 2506.000 2694.650 2510.000 2694.800 ;
        RECT 2519.485 2694.650 2519.815 2694.665 ;
        RECT 2506.000 2694.350 2519.815 2694.650 ;
        RECT 2506.000 2694.200 2510.000 2694.350 ;
        RECT 2519.485 2694.335 2519.815 2694.350 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 467.400 1103.930 467.460 ;
        RECT 2525.930 467.400 2526.250 467.460 ;
        RECT 1103.610 467.260 2526.250 467.400 ;
        RECT 1103.610 467.200 1103.930 467.260 ;
        RECT 2525.930 467.200 2526.250 467.260 ;
        RECT 1102.690 2.960 1103.010 3.020 ;
        RECT 1103.610 2.960 1103.930 3.020 ;
        RECT 1102.690 2.820 1103.930 2.960 ;
        RECT 1102.690 2.760 1103.010 2.820 ;
        RECT 1103.610 2.760 1103.930 2.820 ;
      LAYER via ;
        RECT 1103.640 467.200 1103.900 467.460 ;
        RECT 2525.960 467.200 2526.220 467.460 ;
        RECT 1102.720 2.760 1102.980 3.020 ;
        RECT 1103.640 2.760 1103.900 3.020 ;
      LAYER met2 ;
        RECT 2525.950 1963.995 2526.230 1964.365 ;
        RECT 2526.020 467.490 2526.160 1963.995 ;
        RECT 1103.640 467.170 1103.900 467.490 ;
        RECT 2525.960 467.170 2526.220 467.490 ;
        RECT 1103.700 3.050 1103.840 467.170 ;
        RECT 1102.720 2.730 1102.980 3.050 ;
        RECT 1103.640 2.730 1103.900 3.050 ;
        RECT 1102.780 2.400 1102.920 2.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 2525.950 1964.040 2526.230 1964.320 ;
      LAYER met3 ;
        RECT 2506.000 1964.330 2510.000 1964.480 ;
        RECT 2525.925 1964.330 2526.255 1964.345 ;
        RECT 2506.000 1964.030 2526.255 1964.330 ;
        RECT 2506.000 1963.880 2510.000 1964.030 ;
        RECT 2525.925 1964.015 2526.255 1964.030 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 392.910 162.080 393.230 162.140 ;
        RECT 1117.870 162.080 1118.190 162.140 ;
        RECT 392.910 161.940 1118.190 162.080 ;
        RECT 392.910 161.880 393.230 161.940 ;
        RECT 1117.870 161.880 1118.190 161.940 ;
        RECT 1117.870 2.960 1118.190 3.020 ;
        RECT 1120.630 2.960 1120.950 3.020 ;
        RECT 1117.870 2.820 1120.950 2.960 ;
        RECT 1117.870 2.760 1118.190 2.820 ;
        RECT 1120.630 2.760 1120.950 2.820 ;
      LAYER via ;
        RECT 392.940 161.880 393.200 162.140 ;
        RECT 1117.900 161.880 1118.160 162.140 ;
        RECT 1117.900 2.760 1118.160 3.020 ;
        RECT 1120.660 2.760 1120.920 3.020 ;
      LAYER met2 ;
        RECT 392.930 2174.795 393.210 2175.165 ;
        RECT 393.000 162.170 393.140 2174.795 ;
        RECT 392.940 161.850 393.200 162.170 ;
        RECT 1117.900 161.850 1118.160 162.170 ;
        RECT 1117.960 3.050 1118.100 161.850 ;
        RECT 1117.900 2.730 1118.160 3.050 ;
        RECT 1120.660 2.730 1120.920 3.050 ;
        RECT 1120.720 2.400 1120.860 2.730 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 392.930 2174.840 393.210 2175.120 ;
      LAYER met3 ;
        RECT 392.905 2175.130 393.235 2175.145 ;
        RECT 410.000 2175.130 414.000 2175.280 ;
        RECT 392.905 2174.830 414.000 2175.130 ;
        RECT 392.905 2174.815 393.235 2174.830 ;
        RECT 410.000 2174.680 414.000 2174.830 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1144.550 403.480 1144.870 403.540 ;
        RECT 2527.310 403.480 2527.630 403.540 ;
        RECT 1144.550 403.340 2527.630 403.480 ;
        RECT 1144.550 403.280 1144.870 403.340 ;
        RECT 2527.310 403.280 2527.630 403.340 ;
        RECT 1138.570 18.260 1138.890 18.320 ;
        RECT 1144.550 18.260 1144.870 18.320 ;
        RECT 1138.570 18.120 1144.870 18.260 ;
        RECT 1138.570 18.060 1138.890 18.120 ;
        RECT 1144.550 18.060 1144.870 18.120 ;
      LAYER via ;
        RECT 1144.580 403.280 1144.840 403.540 ;
        RECT 2527.340 403.280 2527.600 403.540 ;
        RECT 1138.600 18.060 1138.860 18.320 ;
        RECT 1144.580 18.060 1144.840 18.320 ;
      LAYER met2 ;
        RECT 2527.330 1507.035 2527.610 1507.405 ;
        RECT 2527.400 403.570 2527.540 1507.035 ;
        RECT 1144.580 403.250 1144.840 403.570 ;
        RECT 2527.340 403.250 2527.600 403.570 ;
        RECT 1144.640 18.350 1144.780 403.250 ;
        RECT 1138.600 18.030 1138.860 18.350 ;
        RECT 1144.580 18.030 1144.840 18.350 ;
        RECT 1138.660 2.400 1138.800 18.030 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
      LAYER via2 ;
        RECT 2527.330 1507.080 2527.610 1507.360 ;
      LAYER met3 ;
        RECT 2506.000 1507.370 2510.000 1507.520 ;
        RECT 2527.305 1507.370 2527.635 1507.385 ;
        RECT 2506.000 1507.070 2527.635 1507.370 ;
        RECT 2506.000 1506.920 2510.000 1507.070 ;
        RECT 2527.305 1507.055 2527.635 1507.070 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 390.220 786.530 390.280 ;
        RECT 1152.370 390.220 1152.690 390.280 ;
        RECT 786.210 390.080 1152.690 390.220 ;
        RECT 786.210 390.020 786.530 390.080 ;
        RECT 1152.370 390.020 1152.690 390.080 ;
      LAYER via ;
        RECT 786.240 390.020 786.500 390.280 ;
        RECT 1152.400 390.020 1152.660 390.280 ;
      LAYER met2 ;
        RECT 782.690 510.410 782.970 514.000 ;
        RECT 782.690 510.270 786.440 510.410 ;
        RECT 782.690 510.000 782.970 510.270 ;
        RECT 786.300 390.310 786.440 510.270 ;
        RECT 786.240 389.990 786.500 390.310 ;
        RECT 1152.400 389.990 1152.660 390.310 ;
        RECT 1152.460 17.410 1152.600 389.990 ;
        RECT 1152.460 17.270 1156.740 17.410 ;
        RECT 1156.600 2.400 1156.740 17.270 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2520.890 1416.595 2521.170 1416.965 ;
        RECT 2520.960 1402.005 2521.100 1416.595 ;
        RECT 2520.890 1401.635 2521.170 1402.005 ;
        RECT 2518.130 1271.755 2518.410 1272.125 ;
        RECT 2518.200 1269.405 2518.340 1271.755 ;
        RECT 2518.130 1269.035 2518.410 1269.405 ;
        RECT 2521.350 971.875 2521.630 972.245 ;
        RECT 2521.420 932.010 2521.560 971.875 ;
        RECT 2520.960 931.870 2521.560 932.010 ;
        RECT 2520.960 926.005 2521.100 931.870 ;
        RECT 2520.890 925.635 2521.170 926.005 ;
        RECT 2521.810 875.315 2522.090 875.685 ;
        RECT 2521.880 829.445 2522.020 875.315 ;
        RECT 2521.810 829.075 2522.090 829.445 ;
        RECT 675.830 396.595 676.110 396.965 ;
        RECT 675.900 16.900 676.040 396.595 ;
        RECT 674.520 16.760 676.040 16.900 ;
        RECT 674.520 2.400 674.660 16.760 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 2520.890 1416.640 2521.170 1416.920 ;
        RECT 2520.890 1401.680 2521.170 1401.960 ;
        RECT 2518.130 1271.800 2518.410 1272.080 ;
        RECT 2518.130 1269.080 2518.410 1269.360 ;
        RECT 2521.350 971.920 2521.630 972.200 ;
        RECT 2520.890 925.680 2521.170 925.960 ;
        RECT 2521.810 875.360 2522.090 875.640 ;
        RECT 2521.810 829.120 2522.090 829.400 ;
        RECT 675.830 396.640 676.110 396.920 ;
      LAYER met3 ;
        RECT 2506.000 1489.690 2510.000 1489.840 ;
        RECT 2520.150 1489.690 2520.530 1489.700 ;
        RECT 2506.000 1489.390 2520.530 1489.690 ;
        RECT 2506.000 1489.240 2510.000 1489.390 ;
        RECT 2520.150 1489.380 2520.530 1489.390 ;
        RECT 2520.150 1416.930 2520.530 1416.940 ;
        RECT 2520.865 1416.930 2521.195 1416.945 ;
        RECT 2520.150 1416.630 2521.195 1416.930 ;
        RECT 2520.150 1416.620 2520.530 1416.630 ;
        RECT 2520.865 1416.615 2521.195 1416.630 ;
        RECT 2520.865 1401.970 2521.195 1401.985 ;
        RECT 2520.190 1401.670 2521.195 1401.970 ;
        RECT 2520.190 1401.300 2520.490 1401.670 ;
        RECT 2520.865 1401.655 2521.195 1401.670 ;
        RECT 2520.150 1400.980 2520.530 1401.300 ;
        RECT 2518.105 1272.090 2518.435 1272.105 ;
        RECT 2520.150 1272.090 2520.530 1272.100 ;
        RECT 2518.105 1271.790 2520.530 1272.090 ;
        RECT 2518.105 1271.775 2518.435 1271.790 ;
        RECT 2520.150 1271.780 2520.530 1271.790 ;
        RECT 2518.105 1269.380 2518.435 1269.385 ;
        RECT 2518.105 1269.370 2518.690 1269.380 ;
        RECT 2518.105 1269.070 2518.890 1269.370 ;
        RECT 2518.105 1269.060 2518.690 1269.070 ;
        RECT 2518.105 1269.055 2518.435 1269.060 ;
        RECT 2518.310 1161.250 2518.690 1161.260 ;
        RECT 2518.310 1160.950 2521.410 1161.250 ;
        RECT 2518.310 1160.940 2518.690 1160.950 ;
        RECT 2519.230 1159.380 2519.610 1159.390 ;
        RECT 2521.110 1159.380 2521.410 1160.950 ;
        RECT 2519.230 1159.080 2521.410 1159.380 ;
        RECT 2519.230 1159.070 2519.610 1159.080 ;
        RECT 2519.230 972.580 2519.610 972.900 ;
        RECT 2519.270 972.210 2519.570 972.580 ;
        RECT 2521.325 972.210 2521.655 972.225 ;
        RECT 2519.270 971.910 2521.655 972.210 ;
        RECT 2521.325 971.895 2521.655 971.910 ;
        RECT 2520.865 925.970 2521.195 925.985 ;
        RECT 2519.270 925.670 2521.195 925.970 ;
        RECT 2519.270 925.300 2519.570 925.670 ;
        RECT 2520.865 925.655 2521.195 925.670 ;
        RECT 2519.230 924.980 2519.610 925.300 ;
        RECT 2519.230 876.020 2519.610 876.340 ;
        RECT 2519.270 875.650 2519.570 876.020 ;
        RECT 2521.785 875.650 2522.115 875.665 ;
        RECT 2519.270 875.350 2522.115 875.650 ;
        RECT 2521.785 875.335 2522.115 875.350 ;
        RECT 2521.785 829.410 2522.115 829.425 ;
        RECT 2518.580 829.110 2522.115 829.410 ;
        RECT 2518.580 828.220 2518.880 829.110 ;
        RECT 2521.785 829.095 2522.115 829.110 ;
        RECT 2519.230 828.220 2519.610 828.230 ;
        RECT 2518.580 827.920 2519.610 828.220 ;
        RECT 2519.230 827.910 2519.610 827.920 ;
        RECT 675.805 396.930 676.135 396.945 ;
        RECT 2519.230 396.930 2519.610 396.940 ;
        RECT 675.805 396.630 2519.610 396.930 ;
        RECT 675.805 396.615 676.135 396.630 ;
        RECT 2519.230 396.620 2519.610 396.630 ;
      LAYER via3 ;
        RECT 2520.180 1489.380 2520.500 1489.700 ;
        RECT 2520.180 1416.620 2520.500 1416.940 ;
        RECT 2520.180 1400.980 2520.500 1401.300 ;
        RECT 2520.180 1271.780 2520.500 1272.100 ;
        RECT 2518.340 1269.060 2518.660 1269.380 ;
        RECT 2518.340 1160.940 2518.660 1161.260 ;
        RECT 2519.260 1159.070 2519.580 1159.390 ;
        RECT 2519.260 972.580 2519.580 972.900 ;
        RECT 2519.260 924.980 2519.580 925.300 ;
        RECT 2519.260 876.020 2519.580 876.340 ;
        RECT 2519.260 827.910 2519.580 828.230 ;
        RECT 2519.260 396.620 2519.580 396.940 ;
      LAYER met4 ;
        RECT 2520.175 1489.375 2520.505 1489.705 ;
        RECT 2520.190 1416.945 2520.490 1489.375 ;
        RECT 2520.175 1416.615 2520.505 1416.945 ;
        RECT 2520.175 1400.975 2520.505 1401.305 ;
        RECT 2520.190 1272.105 2520.490 1400.975 ;
        RECT 2520.175 1271.775 2520.505 1272.105 ;
        RECT 2518.335 1269.055 2518.665 1269.385 ;
        RECT 2518.350 1161.265 2518.650 1269.055 ;
        RECT 2518.335 1160.935 2518.665 1161.265 ;
        RECT 2519.255 1159.065 2519.585 1159.395 ;
        RECT 2519.270 972.905 2519.570 1159.065 ;
        RECT 2519.255 972.575 2519.585 972.905 ;
        RECT 2519.255 924.975 2519.585 925.305 ;
        RECT 2519.270 876.345 2519.570 924.975 ;
        RECT 2519.255 876.015 2519.585 876.345 ;
        RECT 2519.255 827.905 2519.585 828.235 ;
        RECT 2519.270 824.650 2519.570 827.905 ;
        RECT 2518.350 824.350 2519.570 824.650 ;
        RECT 2518.350 729.450 2518.650 824.350 ;
        RECT 2518.350 729.150 2519.570 729.450 ;
        RECT 2519.270 630.850 2519.570 729.150 ;
        RECT 2518.350 630.550 2519.570 630.850 ;
        RECT 2518.350 437.050 2518.650 630.550 ;
        RECT 2518.350 436.750 2519.570 437.050 ;
        RECT 2519.270 396.945 2519.570 436.750 ;
        RECT 2519.255 396.615 2519.585 396.945 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 392.450 251.840 392.770 251.900 ;
        RECT 1173.070 251.840 1173.390 251.900 ;
        RECT 392.450 251.700 1173.390 251.840 ;
        RECT 392.450 251.640 392.770 251.700 ;
        RECT 1173.070 251.640 1173.390 251.700 ;
      LAYER via ;
        RECT 392.480 251.640 392.740 251.900 ;
        RECT 1173.100 251.640 1173.360 251.900 ;
      LAYER met2 ;
        RECT 392.470 2193.835 392.750 2194.205 ;
        RECT 392.540 251.930 392.680 2193.835 ;
        RECT 392.480 251.610 392.740 251.930 ;
        RECT 1173.100 251.610 1173.360 251.930 ;
        RECT 1173.160 16.730 1173.300 251.610 ;
        RECT 1173.160 16.590 1174.220 16.730 ;
        RECT 1174.080 2.400 1174.220 16.590 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 392.470 2193.880 392.750 2194.160 ;
      LAYER met3 ;
        RECT 392.445 2194.170 392.775 2194.185 ;
        RECT 410.000 2194.170 414.000 2194.320 ;
        RECT 392.445 2193.870 414.000 2194.170 ;
        RECT 392.445 2193.855 392.775 2193.870 ;
        RECT 410.000 2193.720 414.000 2193.870 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.605 593.385 414.775 620.415 ;
        RECT 414.605 511.445 414.775 576.215 ;
        RECT 416.445 446.845 416.615 479.655 ;
        RECT 416.905 289.085 417.075 331.075 ;
      LAYER mcon ;
        RECT 414.605 620.245 414.775 620.415 ;
        RECT 414.605 576.045 414.775 576.215 ;
        RECT 416.445 479.485 416.615 479.655 ;
        RECT 416.905 330.905 417.075 331.075 ;
      LAYER met1 ;
        RECT 413.150 673.780 413.470 673.840 ;
        RECT 414.530 673.780 414.850 673.840 ;
        RECT 413.150 673.640 414.850 673.780 ;
        RECT 413.150 673.580 413.470 673.640 ;
        RECT 414.530 673.580 414.850 673.640 ;
        RECT 414.530 620.400 414.850 620.460 ;
        RECT 414.335 620.260 414.850 620.400 ;
        RECT 414.530 620.200 414.850 620.260 ;
        RECT 414.530 593.540 414.850 593.600 ;
        RECT 414.335 593.400 414.850 593.540 ;
        RECT 414.530 593.340 414.850 593.400 ;
        RECT 414.530 576.200 414.850 576.260 ;
        RECT 414.335 576.060 414.850 576.200 ;
        RECT 414.530 576.000 414.850 576.060 ;
        RECT 414.545 511.600 414.835 511.645 ;
        RECT 416.830 511.600 417.150 511.660 ;
        RECT 414.545 511.460 417.150 511.600 ;
        RECT 414.545 511.415 414.835 511.460 ;
        RECT 416.830 511.400 417.150 511.460 ;
        RECT 416.385 479.640 416.675 479.685 ;
        RECT 416.830 479.640 417.150 479.700 ;
        RECT 416.385 479.500 417.150 479.640 ;
        RECT 416.385 479.455 416.675 479.500 ;
        RECT 416.830 479.440 417.150 479.500 ;
        RECT 416.370 447.000 416.690 447.060 ;
        RECT 416.175 446.860 416.690 447.000 ;
        RECT 416.370 446.800 416.690 446.860 ;
        RECT 416.830 331.060 417.150 331.120 ;
        RECT 416.635 330.920 417.150 331.060 ;
        RECT 416.830 330.860 417.150 330.920 ;
        RECT 416.845 289.240 417.135 289.285 ;
        RECT 417.750 289.240 418.070 289.300 ;
        RECT 416.845 289.100 418.070 289.240 ;
        RECT 416.845 289.055 417.135 289.100 ;
        RECT 417.750 289.040 418.070 289.100 ;
        RECT 416.830 231.440 417.150 231.500 ;
        RECT 1187.330 231.440 1187.650 231.500 ;
        RECT 416.830 231.300 1187.650 231.440 ;
        RECT 416.830 231.240 417.150 231.300 ;
        RECT 1187.330 231.240 1187.650 231.300 ;
      LAYER via ;
        RECT 413.180 673.580 413.440 673.840 ;
        RECT 414.560 673.580 414.820 673.840 ;
        RECT 414.560 620.200 414.820 620.460 ;
        RECT 414.560 593.340 414.820 593.600 ;
        RECT 414.560 576.000 414.820 576.260 ;
        RECT 416.860 511.400 417.120 511.660 ;
        RECT 416.860 479.440 417.120 479.700 ;
        RECT 416.400 446.800 416.660 447.060 ;
        RECT 416.860 330.860 417.120 331.120 ;
        RECT 417.780 289.040 418.040 289.300 ;
        RECT 416.860 231.240 417.120 231.500 ;
        RECT 1187.360 231.240 1187.620 231.500 ;
      LAYER met2 ;
        RECT 413.170 674.715 413.450 675.085 ;
        RECT 413.240 673.870 413.380 674.715 ;
        RECT 413.180 673.550 413.440 673.870 ;
        RECT 414.560 673.610 414.820 673.870 ;
        RECT 414.560 673.550 417.060 673.610 ;
        RECT 414.620 673.470 417.060 673.550 ;
        RECT 416.920 662.560 417.060 673.470 ;
        RECT 416.920 662.420 417.520 662.560 ;
        RECT 417.380 643.010 417.520 662.420 ;
        RECT 417.380 642.870 417.980 643.010 ;
        RECT 414.620 620.490 416.600 620.570 ;
        RECT 414.560 620.430 416.600 620.490 ;
        RECT 414.560 620.170 414.820 620.430 ;
        RECT 416.460 619.890 416.600 620.430 ;
        RECT 417.840 619.890 417.980 642.870 ;
        RECT 416.460 619.750 417.980 619.890 ;
        RECT 414.560 593.310 414.820 593.630 ;
        RECT 414.620 576.290 414.760 593.310 ;
        RECT 414.560 575.970 414.820 576.290 ;
        RECT 416.860 511.370 417.120 511.690 ;
        RECT 416.920 479.730 417.060 511.370 ;
        RECT 416.860 479.410 417.120 479.730 ;
        RECT 416.400 446.770 416.660 447.090 ;
        RECT 416.460 424.730 416.600 446.770 ;
        RECT 416.460 424.590 417.980 424.730 ;
        RECT 417.840 386.650 417.980 424.590 ;
        RECT 417.380 386.510 417.980 386.650 ;
        RECT 417.380 338.370 417.520 386.510 ;
        RECT 416.920 338.230 417.520 338.370 ;
        RECT 416.920 331.150 417.060 338.230 ;
        RECT 416.860 330.830 417.120 331.150 ;
        RECT 417.780 289.010 418.040 289.330 ;
        RECT 417.840 255.410 417.980 289.010 ;
        RECT 416.920 255.270 417.980 255.410 ;
        RECT 416.920 231.530 417.060 255.270 ;
        RECT 416.860 231.210 417.120 231.530 ;
        RECT 1187.360 231.210 1187.620 231.530 ;
        RECT 1187.420 17.410 1187.560 231.210 ;
        RECT 1187.420 17.270 1192.160 17.410 ;
        RECT 1192.020 2.400 1192.160 17.270 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 413.170 674.760 413.450 675.040 ;
      LAYER met3 ;
        RECT 410.000 677.320 414.000 677.920 ;
        RECT 413.390 675.065 413.690 677.320 ;
        RECT 413.145 674.750 413.690 675.065 ;
        RECT 413.145 674.735 413.475 674.750 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1209.870 16.560 1210.190 16.620 ;
        RECT 1214.010 16.560 1214.330 16.620 ;
        RECT 1209.870 16.420 1214.330 16.560 ;
        RECT 1209.870 16.360 1210.190 16.420 ;
        RECT 1214.010 16.360 1214.330 16.420 ;
      LAYER via ;
        RECT 1209.900 16.360 1210.160 16.620 ;
        RECT 1214.040 16.360 1214.300 16.620 ;
      LAYER met2 ;
        RECT 1988.670 3032.275 1988.950 3032.645 ;
        RECT 1988.740 3010.000 1988.880 3032.275 ;
        RECT 1988.740 3009.340 1989.090 3010.000 ;
        RECT 1988.810 3006.000 1989.090 3009.340 ;
        RECT 2508.930 2631.755 2509.210 2632.125 ;
        RECT 2509.000 2614.445 2509.140 2631.755 ;
        RECT 2508.930 2614.075 2509.210 2614.445 ;
        RECT 2509.390 919.515 2509.670 919.885 ;
        RECT 2509.460 613.885 2509.600 919.515 ;
        RECT 2509.390 613.515 2509.670 613.885 ;
        RECT 1214.030 485.675 1214.310 486.045 ;
        RECT 1214.100 16.650 1214.240 485.675 ;
        RECT 1209.900 16.330 1210.160 16.650 ;
        RECT 1214.040 16.330 1214.300 16.650 ;
        RECT 1209.960 2.400 1210.100 16.330 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1988.670 3032.320 1988.950 3032.600 ;
        RECT 2508.930 2631.800 2509.210 2632.080 ;
        RECT 2508.930 2614.120 2509.210 2614.400 ;
        RECT 2509.390 919.560 2509.670 919.840 ;
        RECT 2509.390 613.560 2509.670 613.840 ;
        RECT 1214.030 485.720 1214.310 486.000 ;
      LAYER met3 ;
        RECT 1988.645 3032.610 1988.975 3032.625 ;
        RECT 2504.510 3032.610 2504.890 3032.620 ;
        RECT 1988.645 3032.310 2504.890 3032.610 ;
        RECT 1988.645 3032.295 1988.975 3032.310 ;
        RECT 2504.510 3032.300 2504.890 3032.310 ;
        RECT 2506.350 2632.090 2506.730 2632.100 ;
        RECT 2508.905 2632.090 2509.235 2632.105 ;
        RECT 2506.350 2631.790 2509.235 2632.090 ;
        RECT 2506.350 2631.780 2506.730 2631.790 ;
        RECT 2508.905 2631.775 2509.235 2631.790 ;
        RECT 2506.350 2614.410 2506.730 2614.420 ;
        RECT 2508.905 2614.410 2509.235 2614.425 ;
        RECT 2506.350 2614.110 2509.235 2614.410 ;
        RECT 2506.350 2614.100 2506.730 2614.110 ;
        RECT 2508.905 2614.095 2509.235 2614.110 ;
        RECT 2507.270 919.850 2507.650 919.860 ;
        RECT 2509.365 919.850 2509.695 919.865 ;
        RECT 2507.270 919.550 2509.695 919.850 ;
        RECT 2507.270 919.540 2507.650 919.550 ;
        RECT 2509.365 919.535 2509.695 919.550 ;
        RECT 2509.365 613.850 2509.695 613.865 ;
        RECT 2510.030 613.850 2510.410 613.860 ;
        RECT 2509.365 613.550 2510.410 613.850 ;
        RECT 2509.365 613.535 2509.695 613.550 ;
        RECT 2510.030 613.540 2510.410 613.550 ;
        RECT 1214.005 486.010 1214.335 486.025 ;
        RECT 2498.990 486.010 2499.370 486.020 ;
        RECT 1214.005 485.710 2499.370 486.010 ;
        RECT 1214.005 485.695 1214.335 485.710 ;
        RECT 2498.990 485.700 2499.370 485.710 ;
      LAYER via3 ;
        RECT 2504.540 3032.300 2504.860 3032.620 ;
        RECT 2506.380 2631.780 2506.700 2632.100 ;
        RECT 2506.380 2614.100 2506.700 2614.420 ;
        RECT 2507.300 919.540 2507.620 919.860 ;
        RECT 2510.060 613.540 2510.380 613.860 ;
        RECT 2499.020 485.700 2499.340 486.020 ;
      LAYER met4 ;
        RECT 2504.535 3032.295 2504.865 3032.625 ;
        RECT 2504.550 2963.250 2504.850 3032.295 ;
        RECT 2504.550 2962.950 2505.770 2963.250 ;
        RECT 2505.470 2939.450 2505.770 2962.950 ;
        RECT 2505.470 2939.150 2506.690 2939.450 ;
        RECT 2506.390 2895.250 2506.690 2939.150 ;
        RECT 2503.630 2894.950 2506.690 2895.250 ;
        RECT 2503.630 2847.650 2503.930 2894.950 ;
        RECT 2503.630 2847.350 2506.690 2847.650 ;
        RECT 2506.390 2632.105 2506.690 2847.350 ;
        RECT 2506.375 2631.775 2506.705 2632.105 ;
        RECT 2506.375 2614.095 2506.705 2614.425 ;
        RECT 2506.390 2599.450 2506.690 2614.095 ;
        RECT 2504.550 2599.150 2506.690 2599.450 ;
        RECT 2504.550 2572.250 2504.850 2599.150 ;
        RECT 2504.550 2571.950 2508.530 2572.250 ;
        RECT 2508.230 2511.050 2508.530 2571.950 ;
        RECT 2504.550 2510.750 2508.530 2511.050 ;
        RECT 2504.550 2507.650 2504.850 2510.750 ;
        RECT 2502.710 2507.350 2504.850 2507.650 ;
        RECT 2502.710 2426.050 2503.010 2507.350 ;
        RECT 2501.790 2425.750 2503.010 2426.050 ;
        RECT 2501.790 2307.050 2502.090 2425.750 ;
        RECT 2501.790 2306.750 2503.930 2307.050 ;
        RECT 2503.630 2283.250 2503.930 2306.750 ;
        RECT 2502.710 2282.950 2503.930 2283.250 ;
        RECT 2502.710 2150.650 2503.010 2282.950 ;
        RECT 2502.710 2150.350 2504.850 2150.650 ;
        RECT 2504.550 2072.450 2504.850 2150.350 ;
        RECT 2502.710 2072.150 2504.850 2072.450 ;
        RECT 2502.710 1950.050 2503.010 2072.150 ;
        RECT 2502.710 1949.750 2503.930 1950.050 ;
        RECT 2503.630 1868.450 2503.930 1949.750 ;
        RECT 2501.790 1868.150 2503.930 1868.450 ;
        RECT 2501.790 1803.850 2502.090 1868.150 ;
        RECT 2501.790 1803.550 2503.010 1803.850 ;
        RECT 2502.710 1667.850 2503.010 1803.550 ;
        RECT 2501.790 1667.550 2503.010 1667.850 ;
        RECT 2501.790 1664.450 2502.090 1667.550 ;
        RECT 2500.870 1664.150 2502.090 1664.450 ;
        RECT 2500.870 1589.650 2501.170 1664.150 ;
        RECT 2500.870 1589.350 2503.930 1589.650 ;
        RECT 2503.630 1572.650 2503.930 1589.350 ;
        RECT 2502.710 1572.350 2503.930 1572.650 ;
        RECT 2502.710 1565.850 2503.010 1572.350 ;
        RECT 2502.710 1565.550 2503.930 1565.850 ;
        RECT 2503.630 1484.250 2503.930 1565.550 ;
        RECT 2502.710 1483.950 2503.930 1484.250 ;
        RECT 2502.710 1389.050 2503.010 1483.950 ;
        RECT 2500.870 1388.750 2503.010 1389.050 ;
        RECT 2500.870 1232.650 2501.170 1388.750 ;
        RECT 2500.870 1232.350 2503.930 1232.650 ;
        RECT 2503.630 1229.690 2503.930 1232.350 ;
        RECT 2489.390 1228.510 2490.570 1229.690 ;
        RECT 2503.190 1228.510 2504.370 1229.690 ;
        RECT 2489.830 923.690 2490.130 1228.510 ;
        RECT 2489.390 922.510 2490.570 923.690 ;
        RECT 2505.950 922.510 2507.130 923.690 ;
        RECT 2506.390 919.850 2506.690 922.510 ;
        RECT 2507.295 919.850 2507.625 919.865 ;
        RECT 2506.390 919.550 2507.625 919.850 ;
        RECT 2507.295 919.535 2507.625 919.550 ;
        RECT 2510.055 613.535 2510.385 613.865 ;
        RECT 2510.070 580.290 2510.370 613.535 ;
        RECT 2498.590 579.110 2499.770 580.290 ;
        RECT 2509.630 579.110 2510.810 580.290 ;
        RECT 2499.030 486.025 2499.330 579.110 ;
        RECT 2499.015 485.695 2499.345 486.025 ;
      LAYER met5 ;
        RECT 2489.180 1228.300 2504.580 1229.900 ;
        RECT 2489.180 922.300 2507.340 923.900 ;
        RECT 2498.380 578.900 2511.020 580.500 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 390.220 1228.130 390.280 ;
        RECT 2509.370 390.220 2509.690 390.280 ;
        RECT 1227.810 390.080 2509.690 390.220 ;
        RECT 1227.810 390.020 1228.130 390.080 ;
        RECT 2509.370 390.020 2509.690 390.080 ;
      LAYER via ;
        RECT 1227.840 390.020 1228.100 390.280 ;
        RECT 2509.400 390.020 2509.660 390.280 ;
      LAYER met2 ;
        RECT 2509.390 609.435 2509.670 609.805 ;
        RECT 2509.460 390.310 2509.600 609.435 ;
        RECT 1227.840 389.990 1228.100 390.310 ;
        RECT 2509.400 389.990 2509.660 390.310 ;
        RECT 1227.900 2.400 1228.040 389.990 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
      LAYER via2 ;
        RECT 2509.390 609.480 2509.670 609.760 ;
      LAYER met3 ;
        RECT 2506.000 612.040 2510.000 612.640 ;
        RECT 2509.150 609.785 2509.450 612.040 ;
        RECT 2509.150 609.470 2509.695 609.785 ;
        RECT 2509.365 609.455 2509.695 609.470 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1173.240 2520.730 1173.300 ;
        RECT 2583.430 1173.240 2583.750 1173.300 ;
        RECT 2520.410 1173.100 2583.750 1173.240 ;
        RECT 2520.410 1173.040 2520.730 1173.100 ;
        RECT 2583.430 1173.040 2583.750 1173.100 ;
        RECT 1248.510 467.740 1248.830 467.800 ;
        RECT 2583.430 467.740 2583.750 467.800 ;
        RECT 1248.510 467.600 2583.750 467.740 ;
        RECT 1248.510 467.540 1248.830 467.600 ;
        RECT 2583.430 467.540 2583.750 467.600 ;
        RECT 1245.750 16.900 1246.070 16.960 ;
        RECT 1248.510 16.900 1248.830 16.960 ;
        RECT 1245.750 16.760 1248.830 16.900 ;
        RECT 1245.750 16.700 1246.070 16.760 ;
        RECT 1248.510 16.700 1248.830 16.760 ;
      LAYER via ;
        RECT 2520.440 1173.040 2520.700 1173.300 ;
        RECT 2583.460 1173.040 2583.720 1173.300 ;
        RECT 1248.540 467.540 1248.800 467.800 ;
        RECT 2583.460 467.540 2583.720 467.800 ;
        RECT 1245.780 16.700 1246.040 16.960 ;
        RECT 1248.540 16.700 1248.800 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1179.275 2520.710 1179.645 ;
        RECT 2520.500 1173.330 2520.640 1179.275 ;
        RECT 2520.440 1173.010 2520.700 1173.330 ;
        RECT 2583.460 1173.010 2583.720 1173.330 ;
        RECT 2583.520 467.830 2583.660 1173.010 ;
        RECT 1248.540 467.510 1248.800 467.830 ;
        RECT 2583.460 467.510 2583.720 467.830 ;
        RECT 1248.600 16.990 1248.740 467.510 ;
        RECT 1245.780 16.670 1246.040 16.990 ;
        RECT 1248.540 16.670 1248.800 16.990 ;
        RECT 1245.840 2.400 1245.980 16.670 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1179.320 2520.710 1179.600 ;
      LAYER met3 ;
        RECT 2506.000 1179.610 2510.000 1179.760 ;
        RECT 2520.405 1179.610 2520.735 1179.625 ;
        RECT 2506.000 1179.310 2520.735 1179.610 ;
        RECT 2506.000 1179.160 2510.000 1179.310 ;
        RECT 2520.405 1179.295 2520.735 1179.310 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1269.210 431.700 1269.530 431.760 ;
        RECT 2521.330 431.700 2521.650 431.760 ;
        RECT 1269.210 431.560 2521.650 431.700 ;
        RECT 1269.210 431.500 1269.530 431.560 ;
        RECT 2521.330 431.500 2521.650 431.560 ;
        RECT 1263.230 18.260 1263.550 18.320 ;
        RECT 1269.210 18.260 1269.530 18.320 ;
        RECT 1263.230 18.120 1269.530 18.260 ;
        RECT 1263.230 18.060 1263.550 18.120 ;
        RECT 1269.210 18.060 1269.530 18.120 ;
      LAYER via ;
        RECT 1269.240 431.500 1269.500 431.760 ;
        RECT 2521.360 431.500 2521.620 431.760 ;
        RECT 1263.260 18.060 1263.520 18.320 ;
        RECT 1269.240 18.060 1269.500 18.320 ;
      LAYER met2 ;
        RECT 2521.350 923.595 2521.630 923.965 ;
        RECT 2521.420 431.790 2521.560 923.595 ;
        RECT 1269.240 431.470 1269.500 431.790 ;
        RECT 2521.360 431.470 2521.620 431.790 ;
        RECT 1269.300 18.350 1269.440 431.470 ;
        RECT 1263.260 18.030 1263.520 18.350 ;
        RECT 1269.240 18.030 1269.500 18.350 ;
        RECT 1263.320 2.400 1263.460 18.030 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 2521.350 923.640 2521.630 923.920 ;
      LAYER met3 ;
        RECT 2506.000 923.930 2510.000 924.080 ;
        RECT 2521.325 923.930 2521.655 923.945 ;
        RECT 2506.000 923.630 2521.655 923.930 ;
        RECT 2506.000 923.480 2510.000 923.630 ;
        RECT 2521.325 923.615 2521.655 923.630 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.550 334.800 1282.870 334.860 ;
        RECT 1518.070 334.800 1518.390 334.860 ;
        RECT 1282.550 334.660 1518.390 334.800 ;
        RECT 1282.550 334.600 1282.870 334.660 ;
        RECT 1518.070 334.600 1518.390 334.660 ;
      LAYER via ;
        RECT 1282.580 334.600 1282.840 334.860 ;
        RECT 1518.100 334.600 1518.360 334.860 ;
      LAYER met2 ;
        RECT 1524.210 510.410 1524.490 514.000 ;
        RECT 1518.160 510.270 1524.490 510.410 ;
        RECT 1518.160 334.890 1518.300 510.270 ;
        RECT 1524.210 510.000 1524.490 510.270 ;
        RECT 1282.580 334.570 1282.840 334.890 ;
        RECT 1518.100 334.570 1518.360 334.890 ;
        RECT 1282.640 17.410 1282.780 334.570 ;
        RECT 1281.260 17.270 1282.780 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 307.260 1304.030 307.320 ;
        RECT 2511.670 307.260 2511.990 307.320 ;
        RECT 1303.710 307.120 2511.990 307.260 ;
        RECT 1303.710 307.060 1304.030 307.120 ;
        RECT 2511.670 307.060 2511.990 307.120 ;
        RECT 1299.110 29.480 1299.430 29.540 ;
        RECT 1303.710 29.480 1304.030 29.540 ;
        RECT 1299.110 29.340 1304.030 29.480 ;
        RECT 1299.110 29.280 1299.430 29.340 ;
        RECT 1303.710 29.280 1304.030 29.340 ;
      LAYER via ;
        RECT 1303.740 307.060 1304.000 307.320 ;
        RECT 2511.700 307.060 2511.960 307.320 ;
        RECT 1299.140 29.280 1299.400 29.540 ;
        RECT 1303.740 29.280 1304.000 29.540 ;
      LAYER met2 ;
        RECT 2511.690 2256.395 2511.970 2256.765 ;
        RECT 2511.760 307.350 2511.900 2256.395 ;
        RECT 1303.740 307.030 1304.000 307.350 ;
        RECT 2511.700 307.030 2511.960 307.350 ;
        RECT 1303.800 29.570 1303.940 307.030 ;
        RECT 1299.140 29.250 1299.400 29.570 ;
        RECT 1303.740 29.250 1304.000 29.570 ;
        RECT 1299.200 2.400 1299.340 29.250 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
      LAYER via2 ;
        RECT 2511.690 2256.440 2511.970 2256.720 ;
      LAYER met3 ;
        RECT 2506.000 2256.730 2510.000 2256.880 ;
        RECT 2511.665 2256.730 2511.995 2256.745 ;
        RECT 2506.000 2256.430 2511.995 2256.730 ;
        RECT 2506.000 2256.280 2510.000 2256.430 ;
        RECT 2511.665 2256.415 2511.995 2256.430 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 358.410 3018.080 358.730 3018.140 ;
        RECT 628.890 3018.080 629.210 3018.140 ;
        RECT 358.410 3017.940 629.210 3018.080 ;
        RECT 358.410 3017.880 358.730 3017.940 ;
        RECT 628.890 3017.880 629.210 3017.940 ;
      LAYER via ;
        RECT 358.440 3017.880 358.700 3018.140 ;
        RECT 628.920 3017.880 629.180 3018.140 ;
      LAYER met2 ;
        RECT 358.440 3017.850 358.700 3018.170 ;
        RECT 628.920 3017.850 629.180 3018.170 ;
        RECT 358.500 18.205 358.640 3017.850 ;
        RECT 628.980 3010.000 629.120 3017.850 ;
        RECT 628.980 3009.340 629.330 3010.000 ;
        RECT 629.050 3006.000 629.330 3009.340 ;
        RECT 358.430 17.835 358.710 18.205 ;
        RECT 1316.610 17.835 1316.890 18.205 ;
        RECT 1316.680 16.050 1316.820 17.835 ;
        RECT 1316.680 15.910 1317.280 16.050 ;
        RECT 1317.140 2.400 1317.280 15.910 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 358.430 17.880 358.710 18.160 ;
        RECT 1316.610 17.880 1316.890 18.160 ;
      LAYER met3 ;
        RECT 358.405 18.170 358.735 18.185 ;
        RECT 1316.585 18.170 1316.915 18.185 ;
        RECT 358.405 17.870 1316.915 18.170 ;
        RECT 358.405 17.855 358.735 17.870 ;
        RECT 1316.585 17.855 1316.915 17.870 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.790 356.475 1332.070 356.845 ;
        RECT 1331.860 17.410 1332.000 356.475 ;
        RECT 1331.860 17.270 1335.220 17.410 ;
        RECT 1335.080 2.400 1335.220 17.270 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
      LAYER via2 ;
        RECT 1331.790 356.520 1332.070 356.800 ;
      LAYER met3 ;
        RECT 392.190 2942.170 392.570 2942.180 ;
        RECT 410.000 2942.170 414.000 2942.320 ;
        RECT 392.190 2941.870 414.000 2942.170 ;
        RECT 392.190 2941.860 392.570 2941.870 ;
        RECT 410.000 2941.720 414.000 2941.870 ;
        RECT 392.190 356.810 392.570 356.820 ;
        RECT 1331.765 356.810 1332.095 356.825 ;
        RECT 392.190 356.510 1332.095 356.810 ;
        RECT 392.190 356.500 392.570 356.510 ;
        RECT 1331.765 356.495 1332.095 356.510 ;
      LAYER via3 ;
        RECT 392.220 2941.860 392.540 2942.180 ;
        RECT 392.220 356.500 392.540 356.820 ;
      LAYER met4 ;
        RECT 392.215 2941.855 392.545 2942.185 ;
        RECT 392.230 356.825 392.530 2941.855 ;
        RECT 392.215 356.495 392.545 356.825 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 33.220 692.690 33.280 ;
        RECT 1283.470 33.220 1283.790 33.280 ;
        RECT 692.370 33.080 1283.790 33.220 ;
        RECT 692.370 33.020 692.690 33.080 ;
        RECT 1283.470 33.020 1283.790 33.080 ;
      LAYER via ;
        RECT 692.400 33.020 692.660 33.280 ;
        RECT 1283.500 33.020 1283.760 33.280 ;
      LAYER met2 ;
        RECT 1289.610 510.410 1289.890 514.000 ;
        RECT 1283.560 510.270 1289.890 510.410 ;
        RECT 1283.560 33.310 1283.700 510.270 ;
        RECT 1289.610 510.000 1289.890 510.270 ;
        RECT 692.400 32.990 692.660 33.310 ;
        RECT 1283.500 32.990 1283.760 33.310 ;
        RECT 692.460 2.400 692.600 32.990 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.250 3024.540 2062.570 3024.600 ;
        RECT 2566.870 3024.540 2567.190 3024.600 ;
        RECT 2062.250 3024.400 2567.190 3024.540 ;
        RECT 2062.250 3024.340 2062.570 3024.400 ;
        RECT 2566.870 3024.340 2567.190 3024.400 ;
        RECT 1352.470 18.600 1352.790 18.660 ;
        RECT 2566.870 18.600 2567.190 18.660 ;
        RECT 1352.470 18.460 2567.190 18.600 ;
        RECT 1352.470 18.400 1352.790 18.460 ;
        RECT 2566.870 18.400 2567.190 18.460 ;
      LAYER via ;
        RECT 2062.280 3024.340 2062.540 3024.600 ;
        RECT 2566.900 3024.340 2567.160 3024.600 ;
        RECT 1352.500 18.400 1352.760 18.660 ;
        RECT 2566.900 18.400 2567.160 18.660 ;
      LAYER met2 ;
        RECT 2062.280 3024.310 2062.540 3024.630 ;
        RECT 2566.900 3024.310 2567.160 3024.630 ;
        RECT 2062.340 3010.000 2062.480 3024.310 ;
        RECT 2062.340 3009.340 2062.690 3010.000 ;
        RECT 2062.410 3006.000 2062.690 3009.340 ;
        RECT 2566.960 18.690 2567.100 3024.310 ;
        RECT 1352.500 18.370 1352.760 18.690 ;
        RECT 2566.900 18.370 2567.160 18.690 ;
        RECT 1352.560 2.400 1352.700 18.370 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 20.300 1370.730 20.360 ;
        RECT 1372.710 20.300 1373.030 20.360 ;
        RECT 1370.410 20.160 1373.030 20.300 ;
        RECT 1370.410 20.100 1370.730 20.160 ;
        RECT 1372.710 20.100 1373.030 20.160 ;
      LAYER via ;
        RECT 1370.440 20.100 1370.700 20.360 ;
        RECT 1372.740 20.100 1373.000 20.360 ;
      LAYER met2 ;
        RECT 1926.110 3031.595 1926.390 3031.965 ;
        RECT 1926.180 3010.000 1926.320 3031.595 ;
        RECT 1926.180 3009.340 1926.530 3010.000 ;
        RECT 1926.250 3006.000 1926.530 3009.340 ;
        RECT 1372.730 512.195 1373.010 512.565 ;
        RECT 1372.800 20.390 1372.940 512.195 ;
        RECT 1370.440 20.070 1370.700 20.390 ;
        RECT 1372.740 20.070 1373.000 20.390 ;
        RECT 1370.500 2.400 1370.640 20.070 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
      LAYER via2 ;
        RECT 1926.110 3031.640 1926.390 3031.920 ;
        RECT 1372.730 512.240 1373.010 512.520 ;
      LAYER met3 ;
        RECT 1926.085 3031.930 1926.415 3031.945 ;
        RECT 2511.870 3031.930 2512.250 3031.940 ;
        RECT 1926.085 3031.630 2512.250 3031.930 ;
        RECT 1926.085 3031.615 1926.415 3031.630 ;
        RECT 2511.870 3031.620 2512.250 3031.630 ;
        RECT 2511.870 513.890 2512.250 513.900 ;
        RECT 1372.950 513.590 2512.250 513.890 ;
        RECT 1372.950 512.545 1373.250 513.590 ;
        RECT 2511.870 513.580 2512.250 513.590 ;
        RECT 1372.705 512.230 1373.250 512.545 ;
        RECT 1372.705 512.215 1373.035 512.230 ;
      LAYER via3 ;
        RECT 2511.900 3031.620 2512.220 3031.940 ;
        RECT 2511.900 513.580 2512.220 513.900 ;
      LAYER met4 ;
        RECT 2511.895 3031.615 2512.225 3031.945 ;
        RECT 2511.910 513.905 2512.210 3031.615 ;
        RECT 2511.895 513.575 2512.225 513.905 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.410 459.240 1393.730 459.300 ;
        RECT 2525.470 459.240 2525.790 459.300 ;
        RECT 1393.410 459.100 2525.790 459.240 ;
        RECT 1393.410 459.040 1393.730 459.100 ;
        RECT 2525.470 459.040 2525.790 459.100 ;
        RECT 1388.350 16.220 1388.670 16.280 ;
        RECT 1393.410 16.220 1393.730 16.280 ;
        RECT 1388.350 16.080 1393.730 16.220 ;
        RECT 1388.350 16.020 1388.670 16.080 ;
        RECT 1393.410 16.020 1393.730 16.080 ;
      LAYER via ;
        RECT 1393.440 459.040 1393.700 459.300 ;
        RECT 2525.500 459.040 2525.760 459.300 ;
        RECT 1388.380 16.020 1388.640 16.280 ;
        RECT 1393.440 16.020 1393.700 16.280 ;
      LAYER met2 ;
        RECT 2525.490 1983.035 2525.770 1983.405 ;
        RECT 2525.560 459.330 2525.700 1983.035 ;
        RECT 1393.440 459.010 1393.700 459.330 ;
        RECT 2525.500 459.010 2525.760 459.330 ;
        RECT 1393.500 16.310 1393.640 459.010 ;
        RECT 1388.380 15.990 1388.640 16.310 ;
        RECT 1393.440 15.990 1393.700 16.310 ;
        RECT 1388.440 2.400 1388.580 15.990 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
      LAYER via2 ;
        RECT 2525.490 1983.080 2525.770 1983.360 ;
      LAYER met3 ;
        RECT 2506.000 1983.370 2510.000 1983.520 ;
        RECT 2525.465 1983.370 2525.795 1983.385 ;
        RECT 2506.000 1983.070 2525.795 1983.370 ;
        RECT 2506.000 1982.920 2510.000 1983.070 ;
        RECT 2525.465 1983.055 2525.795 1983.070 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.145 2209.745 414.315 2221.815 ;
        RECT 414.145 1471.265 414.315 1473.815 ;
        RECT 414.605 1038.445 414.775 1095.055 ;
        RECT 414.145 791.945 414.315 866.915 ;
        RECT 413.685 717.825 413.855 725.135 ;
        RECT 456.465 512.125 456.635 513.995 ;
        RECT 520.865 512.125 521.035 513.995 ;
        RECT 569.165 512.125 569.335 513.995 ;
        RECT 603.665 512.125 603.835 513.995 ;
        RECT 636.785 512.125 636.955 513.995 ;
        RECT 713.605 512.125 713.775 513.995 ;
        RECT 724.645 512.465 724.815 513.995 ;
        RECT 766.045 511.785 766.215 512.635 ;
        RECT 813.885 511.785 814.055 513.995 ;
        RECT 814.345 512.465 814.515 513.995 ;
        RECT 862.645 511.785 862.815 512.635 ;
        RECT 910.485 511.785 910.655 513.995 ;
        RECT 966.145 513.145 966.315 513.995 ;
        RECT 1076.085 513.485 1076.715 513.655 ;
        RECT 1111.045 512.465 1111.215 513.315 ;
        RECT 1134.965 512.465 1135.135 513.655 ;
        RECT 1402.685 496.485 1402.855 513.655 ;
        RECT 1402.225 386.325 1402.395 434.775 ;
        RECT 1401.765 241.485 1401.935 289.595 ;
        RECT 1401.765 158.525 1401.935 193.035 ;
      LAYER mcon ;
        RECT 414.145 2221.645 414.315 2221.815 ;
        RECT 414.145 1473.645 414.315 1473.815 ;
        RECT 414.605 1094.885 414.775 1095.055 ;
        RECT 414.145 866.745 414.315 866.915 ;
        RECT 413.685 724.965 413.855 725.135 ;
        RECT 456.465 513.825 456.635 513.995 ;
        RECT 520.865 513.825 521.035 513.995 ;
        RECT 569.165 513.825 569.335 513.995 ;
        RECT 603.665 513.825 603.835 513.995 ;
        RECT 636.785 513.825 636.955 513.995 ;
        RECT 713.605 513.825 713.775 513.995 ;
        RECT 724.645 513.825 724.815 513.995 ;
        RECT 813.885 513.825 814.055 513.995 ;
        RECT 766.045 512.465 766.215 512.635 ;
        RECT 814.345 513.825 814.515 513.995 ;
        RECT 910.485 513.825 910.655 513.995 ;
        RECT 862.645 512.465 862.815 512.635 ;
        RECT 966.145 513.825 966.315 513.995 ;
        RECT 1076.545 513.485 1076.715 513.655 ;
        RECT 1134.965 513.485 1135.135 513.655 ;
        RECT 1111.045 513.145 1111.215 513.315 ;
        RECT 1402.685 513.485 1402.855 513.655 ;
        RECT 1402.225 434.605 1402.395 434.775 ;
        RECT 1401.765 289.425 1401.935 289.595 ;
        RECT 1401.765 192.865 1401.935 193.035 ;
      LAYER met1 ;
        RECT 417.290 3010.260 417.610 3010.320 ;
        RECT 1134.430 3010.260 1134.750 3010.320 ;
        RECT 417.290 3010.120 1134.750 3010.260 ;
        RECT 417.290 3010.060 417.610 3010.120 ;
        RECT 1134.430 3010.060 1134.750 3010.120 ;
        RECT 414.085 2221.800 414.375 2221.845 ;
        RECT 414.530 2221.800 414.850 2221.860 ;
        RECT 414.085 2221.660 414.850 2221.800 ;
        RECT 414.085 2221.615 414.375 2221.660 ;
        RECT 414.530 2221.600 414.850 2221.660 ;
        RECT 414.085 2209.900 414.375 2209.945 ;
        RECT 414.530 2209.900 414.850 2209.960 ;
        RECT 414.085 2209.760 414.850 2209.900 ;
        RECT 414.085 2209.715 414.375 2209.760 ;
        RECT 414.530 2209.700 414.850 2209.760 ;
        RECT 414.085 1473.800 414.375 1473.845 ;
        RECT 414.530 1473.800 414.850 1473.860 ;
        RECT 414.085 1473.660 414.850 1473.800 ;
        RECT 414.085 1473.615 414.375 1473.660 ;
        RECT 414.530 1473.600 414.850 1473.660 ;
        RECT 414.085 1471.420 414.375 1471.465 ;
        RECT 414.530 1471.420 414.850 1471.480 ;
        RECT 414.085 1471.280 414.850 1471.420 ;
        RECT 414.085 1471.235 414.375 1471.280 ;
        RECT 414.530 1471.220 414.850 1471.280 ;
        RECT 414.530 1095.040 414.850 1095.100 ;
        RECT 414.335 1094.900 414.850 1095.040 ;
        RECT 414.530 1094.840 414.850 1094.900 ;
        RECT 414.530 1038.600 414.850 1038.660 ;
        RECT 414.335 1038.460 414.850 1038.600 ;
        RECT 414.530 1038.400 414.850 1038.460 ;
        RECT 414.085 866.900 414.375 866.945 ;
        RECT 414.530 866.900 414.850 866.960 ;
        RECT 414.085 866.760 414.850 866.900 ;
        RECT 414.085 866.715 414.375 866.760 ;
        RECT 414.530 866.700 414.850 866.760 ;
        RECT 414.085 792.100 414.375 792.145 ;
        RECT 414.530 792.100 414.850 792.160 ;
        RECT 414.085 791.960 414.850 792.100 ;
        RECT 414.085 791.915 414.375 791.960 ;
        RECT 414.530 791.900 414.850 791.960 ;
        RECT 413.625 725.120 413.915 725.165 ;
        RECT 414.530 725.120 414.850 725.180 ;
        RECT 413.625 724.980 414.850 725.120 ;
        RECT 413.625 724.935 413.915 724.980 ;
        RECT 414.530 724.920 414.850 724.980 ;
        RECT 413.625 717.980 413.915 718.025 ;
        RECT 414.530 717.980 414.850 718.040 ;
        RECT 413.625 717.840 414.850 717.980 ;
        RECT 413.625 717.795 413.915 717.840 ;
        RECT 414.530 717.780 414.850 717.840 ;
        RECT 713.620 514.180 724.800 514.320 ;
        RECT 413.610 513.980 413.930 514.040 ;
        RECT 713.620 514.025 713.760 514.180 ;
        RECT 724.660 514.025 724.800 514.180 ;
        RECT 813.900 514.180 814.500 514.320 ;
        RECT 813.900 514.025 814.040 514.180 ;
        RECT 814.360 514.025 814.500 514.180 ;
        RECT 937.180 514.180 966.300 514.320 ;
        RECT 456.405 513.980 456.695 514.025 ;
        RECT 413.610 513.840 456.695 513.980 ;
        RECT 413.610 513.780 413.930 513.840 ;
        RECT 456.405 513.795 456.695 513.840 ;
        RECT 520.805 513.980 521.095 514.025 ;
        RECT 569.105 513.980 569.395 514.025 ;
        RECT 520.805 513.840 569.395 513.980 ;
        RECT 520.805 513.795 521.095 513.840 ;
        RECT 569.105 513.795 569.395 513.840 ;
        RECT 603.605 513.980 603.895 514.025 ;
        RECT 636.725 513.980 637.015 514.025 ;
        RECT 603.605 513.840 637.015 513.980 ;
        RECT 603.605 513.795 603.895 513.840 ;
        RECT 636.725 513.795 637.015 513.840 ;
        RECT 713.545 513.795 713.835 514.025 ;
        RECT 724.585 513.795 724.875 514.025 ;
        RECT 813.825 513.795 814.115 514.025 ;
        RECT 814.285 513.795 814.575 514.025 ;
        RECT 910.425 513.980 910.715 514.025 ;
        RECT 937.180 513.980 937.320 514.180 ;
        RECT 966.160 514.025 966.300 514.180 ;
        RECT 910.425 513.840 937.320 513.980 ;
        RECT 910.425 513.795 910.715 513.840 ;
        RECT 966.085 513.795 966.375 514.025 ;
        RECT 1008.480 513.840 1027.940 513.980 ;
        RECT 966.085 513.300 966.375 513.345 ;
        RECT 1008.480 513.300 1008.620 513.840 ;
        RECT 1027.800 513.640 1027.940 513.840 ;
        RECT 1173.160 513.840 1221.600 513.980 ;
        RECT 1076.025 513.640 1076.315 513.685 ;
        RECT 1027.800 513.500 1076.315 513.640 ;
        RECT 1076.025 513.455 1076.315 513.500 ;
        RECT 1076.485 513.640 1076.775 513.685 ;
        RECT 1134.905 513.640 1135.195 513.685 ;
        RECT 1173.160 513.640 1173.300 513.840 ;
        RECT 1076.485 513.500 1082.680 513.640 ;
        RECT 1076.485 513.455 1076.775 513.500 ;
        RECT 966.085 513.160 1008.620 513.300 ;
        RECT 1082.540 513.300 1082.680 513.500 ;
        RECT 1134.905 513.500 1173.300 513.640 ;
        RECT 1221.460 513.640 1221.600 513.840 ;
        RECT 1269.760 513.840 1318.200 513.980 ;
        RECT 1269.760 513.640 1269.900 513.840 ;
        RECT 1221.460 513.500 1269.900 513.640 ;
        RECT 1318.060 513.640 1318.200 513.840 ;
        RECT 1402.625 513.640 1402.915 513.685 ;
        RECT 1318.060 513.500 1402.915 513.640 ;
        RECT 1134.905 513.455 1135.195 513.500 ;
        RECT 1402.625 513.455 1402.915 513.500 ;
        RECT 1110.985 513.300 1111.275 513.345 ;
        RECT 1082.540 513.160 1111.275 513.300 ;
        RECT 966.085 513.115 966.375 513.160 ;
        RECT 1110.985 513.115 1111.275 513.160 ;
        RECT 724.585 512.620 724.875 512.665 ;
        RECT 765.985 512.620 766.275 512.665 ;
        RECT 724.585 512.480 766.275 512.620 ;
        RECT 724.585 512.435 724.875 512.480 ;
        RECT 765.985 512.435 766.275 512.480 ;
        RECT 814.285 512.620 814.575 512.665 ;
        RECT 862.585 512.620 862.875 512.665 ;
        RECT 814.285 512.480 862.875 512.620 ;
        RECT 814.285 512.435 814.575 512.480 ;
        RECT 862.585 512.435 862.875 512.480 ;
        RECT 1110.985 512.620 1111.275 512.665 ;
        RECT 1134.905 512.620 1135.195 512.665 ;
        RECT 1110.985 512.480 1135.195 512.620 ;
        RECT 1110.985 512.435 1111.275 512.480 ;
        RECT 1134.905 512.435 1135.195 512.480 ;
        RECT 456.405 512.280 456.695 512.325 ;
        RECT 520.805 512.280 521.095 512.325 ;
        RECT 456.405 512.140 521.095 512.280 ;
        RECT 456.405 512.095 456.695 512.140 ;
        RECT 520.805 512.095 521.095 512.140 ;
        RECT 569.105 512.280 569.395 512.325 ;
        RECT 603.605 512.280 603.895 512.325 ;
        RECT 569.105 512.140 603.895 512.280 ;
        RECT 569.105 512.095 569.395 512.140 ;
        RECT 603.605 512.095 603.895 512.140 ;
        RECT 636.725 512.280 637.015 512.325 ;
        RECT 713.545 512.280 713.835 512.325 ;
        RECT 636.725 512.140 713.835 512.280 ;
        RECT 636.725 512.095 637.015 512.140 ;
        RECT 713.545 512.095 713.835 512.140 ;
        RECT 765.985 511.940 766.275 511.985 ;
        RECT 813.825 511.940 814.115 511.985 ;
        RECT 765.985 511.800 814.115 511.940 ;
        RECT 765.985 511.755 766.275 511.800 ;
        RECT 813.825 511.755 814.115 511.800 ;
        RECT 862.585 511.940 862.875 511.985 ;
        RECT 910.425 511.940 910.715 511.985 ;
        RECT 862.585 511.800 910.715 511.940 ;
        RECT 862.585 511.755 862.875 511.800 ;
        RECT 910.425 511.755 910.715 511.800 ;
        RECT 1402.610 496.640 1402.930 496.700 ;
        RECT 1402.415 496.500 1402.930 496.640 ;
        RECT 1402.610 496.440 1402.930 496.500 ;
        RECT 1402.165 434.760 1402.455 434.805 ;
        RECT 1402.610 434.760 1402.930 434.820 ;
        RECT 1402.165 434.620 1402.930 434.760 ;
        RECT 1402.165 434.575 1402.455 434.620 ;
        RECT 1402.610 434.560 1402.930 434.620 ;
        RECT 1402.150 386.480 1402.470 386.540 ;
        RECT 1401.955 386.340 1402.470 386.480 ;
        RECT 1402.150 386.280 1402.470 386.340 ;
        RECT 1401.230 352.140 1401.550 352.200 ;
        RECT 1401.230 352.000 1401.920 352.140 ;
        RECT 1401.230 351.940 1401.550 352.000 ;
        RECT 1401.780 351.860 1401.920 352.000 ;
        RECT 1401.690 351.600 1402.010 351.860 ;
        RECT 1401.705 289.580 1401.995 289.625 ;
        RECT 1402.150 289.580 1402.470 289.640 ;
        RECT 1401.705 289.440 1402.470 289.580 ;
        RECT 1401.705 289.395 1401.995 289.440 ;
        RECT 1402.150 289.380 1402.470 289.440 ;
        RECT 1401.690 241.640 1402.010 241.700 ;
        RECT 1401.495 241.500 1402.010 241.640 ;
        RECT 1401.690 241.440 1402.010 241.500 ;
        RECT 1401.705 193.020 1401.995 193.065 ;
        RECT 1402.150 193.020 1402.470 193.080 ;
        RECT 1401.705 192.880 1402.470 193.020 ;
        RECT 1401.705 192.835 1401.995 192.880 ;
        RECT 1402.150 192.820 1402.470 192.880 ;
        RECT 1401.690 158.680 1402.010 158.740 ;
        RECT 1401.495 158.540 1402.010 158.680 ;
        RECT 1401.690 158.480 1402.010 158.540 ;
        RECT 1401.230 62.120 1401.550 62.180 ;
        RECT 1405.830 62.120 1406.150 62.180 ;
        RECT 1401.230 61.980 1406.150 62.120 ;
        RECT 1401.230 61.920 1401.550 61.980 ;
        RECT 1405.830 61.920 1406.150 61.980 ;
      LAYER via ;
        RECT 417.320 3010.060 417.580 3010.320 ;
        RECT 1134.460 3010.060 1134.720 3010.320 ;
        RECT 414.560 2221.600 414.820 2221.860 ;
        RECT 414.560 2209.700 414.820 2209.960 ;
        RECT 414.560 1473.600 414.820 1473.860 ;
        RECT 414.560 1471.220 414.820 1471.480 ;
        RECT 414.560 1094.840 414.820 1095.100 ;
        RECT 414.560 1038.400 414.820 1038.660 ;
        RECT 414.560 866.700 414.820 866.960 ;
        RECT 414.560 791.900 414.820 792.160 ;
        RECT 414.560 724.920 414.820 725.180 ;
        RECT 414.560 717.780 414.820 718.040 ;
        RECT 413.640 513.780 413.900 514.040 ;
        RECT 1402.640 496.440 1402.900 496.700 ;
        RECT 1402.640 434.560 1402.900 434.820 ;
        RECT 1402.180 386.280 1402.440 386.540 ;
        RECT 1401.260 351.940 1401.520 352.200 ;
        RECT 1401.720 351.600 1401.980 351.860 ;
        RECT 1402.180 289.380 1402.440 289.640 ;
        RECT 1401.720 241.440 1401.980 241.700 ;
        RECT 1402.180 192.820 1402.440 193.080 ;
        RECT 1401.720 158.480 1401.980 158.740 ;
        RECT 1401.260 61.920 1401.520 62.180 ;
        RECT 1405.860 61.920 1406.120 62.180 ;
      LAYER met2 ;
        RECT 417.320 3010.030 417.580 3010.350 ;
        RECT 1134.460 3010.030 1134.720 3010.350 ;
        RECT 417.380 3006.010 417.520 3010.030 ;
        RECT 1134.520 3009.410 1134.660 3010.030 ;
        RECT 1135.970 3009.410 1136.250 3010.000 ;
        RECT 1134.520 3009.270 1136.250 3009.410 ;
        RECT 417.380 3005.870 417.980 3006.010 ;
        RECT 1135.970 3006.000 1136.250 3009.270 ;
        RECT 417.840 2531.370 417.980 3005.870 ;
        RECT 414.160 2531.230 417.980 2531.370 ;
        RECT 414.160 2496.010 414.300 2531.230 ;
        RECT 414.160 2495.870 416.140 2496.010 ;
        RECT 416.000 2466.090 416.140 2495.870 ;
        RECT 414.620 2465.950 416.140 2466.090 ;
        RECT 414.620 2374.290 414.760 2465.950 ;
        RECT 414.620 2374.150 418.440 2374.290 ;
        RECT 418.300 2332.130 418.440 2374.150 ;
        RECT 417.840 2331.990 418.440 2332.130 ;
        RECT 417.840 2317.850 417.980 2331.990 ;
        RECT 416.920 2317.710 417.980 2317.850 ;
        RECT 416.920 2270.250 417.060 2317.710 ;
        RECT 416.920 2270.110 417.980 2270.250 ;
        RECT 417.840 2255.970 417.980 2270.110 ;
        RECT 417.840 2255.830 418.440 2255.970 ;
        RECT 418.300 2238.290 418.440 2255.830 ;
        RECT 414.620 2238.150 418.440 2238.290 ;
        RECT 414.620 2221.890 414.760 2238.150 ;
        RECT 414.560 2221.570 414.820 2221.890 ;
        RECT 414.560 2209.730 414.820 2209.990 ;
        RECT 414.560 2209.670 416.140 2209.730 ;
        RECT 414.620 2209.590 416.140 2209.670 ;
        RECT 416.000 2160.090 416.140 2209.590 ;
        RECT 416.000 2159.950 417.520 2160.090 ;
        RECT 417.380 2115.210 417.520 2159.950 ;
        RECT 416.920 2115.070 417.520 2115.210 ;
        RECT 416.920 2109.090 417.060 2115.070 ;
        RECT 416.920 2108.950 417.520 2109.090 ;
        RECT 417.380 2092.090 417.520 2108.950 ;
        RECT 416.920 2091.950 417.520 2092.090 ;
        RECT 416.920 2063.360 417.060 2091.950 ;
        RECT 416.920 2063.220 417.520 2063.360 ;
        RECT 417.380 2054.690 417.520 2063.220 ;
        RECT 416.000 2054.550 417.520 2054.690 ;
        RECT 416.000 2051.970 416.140 2054.550 ;
        RECT 416.000 2051.830 417.060 2051.970 ;
        RECT 416.920 2028.850 417.060 2051.830 ;
        RECT 416.920 2028.710 417.980 2028.850 ;
        RECT 417.840 2014.570 417.980 2028.710 ;
        RECT 416.920 2014.430 417.980 2014.570 ;
        RECT 416.920 1994.170 417.060 2014.430 ;
        RECT 416.460 1994.030 417.060 1994.170 ;
        RECT 416.460 1973.090 416.600 1994.030 ;
        RECT 416.460 1972.950 417.060 1973.090 ;
        RECT 416.920 1932.120 417.060 1972.950 ;
        RECT 416.920 1931.980 417.980 1932.120 ;
        RECT 417.840 1930.930 417.980 1931.980 ;
        RECT 414.620 1930.790 417.980 1930.930 ;
        RECT 414.620 1874.490 414.760 1930.790 ;
        RECT 414.620 1874.350 417.060 1874.490 ;
        RECT 416.920 1849.330 417.060 1874.350 ;
        RECT 416.920 1849.190 417.980 1849.330 ;
        RECT 417.840 1803.770 417.980 1849.190 ;
        RECT 416.920 1803.630 417.980 1803.770 ;
        RECT 416.920 1740.530 417.060 1803.630 ;
        RECT 416.920 1740.390 417.980 1740.530 ;
        RECT 417.840 1711.970 417.980 1740.390 ;
        RECT 414.620 1711.830 417.980 1711.970 ;
        RECT 414.620 1684.770 414.760 1711.830 ;
        RECT 414.620 1684.630 417.520 1684.770 ;
        RECT 417.380 1666.410 417.520 1684.630 ;
        RECT 416.920 1666.270 417.520 1666.410 ;
        RECT 416.920 1618.130 417.060 1666.270 ;
        RECT 416.460 1617.990 417.060 1618.130 ;
        RECT 416.460 1606.570 416.600 1617.990 ;
        RECT 416.460 1606.430 417.520 1606.570 ;
        RECT 417.380 1593.650 417.520 1606.430 ;
        RECT 416.920 1593.510 417.520 1593.650 ;
        RECT 416.920 1590.930 417.060 1593.510 ;
        RECT 416.920 1590.790 417.520 1590.930 ;
        RECT 417.380 1569.850 417.520 1590.790 ;
        RECT 416.920 1569.710 417.520 1569.850 ;
        RECT 416.920 1560.330 417.060 1569.710 ;
        RECT 416.920 1560.190 417.520 1560.330 ;
        RECT 417.380 1510.010 417.520 1560.190 ;
        RECT 416.920 1509.870 417.520 1510.010 ;
        RECT 416.920 1509.330 417.060 1509.870 ;
        RECT 416.460 1509.190 417.060 1509.330 ;
        RECT 416.460 1497.090 416.600 1509.190 ;
        RECT 414.620 1496.950 416.600 1497.090 ;
        RECT 414.620 1473.890 414.760 1496.950 ;
        RECT 414.560 1473.570 414.820 1473.890 ;
        RECT 414.560 1471.190 414.820 1471.510 ;
        RECT 414.620 1462.410 414.760 1471.190 ;
        RECT 414.620 1462.270 415.680 1462.410 ;
        RECT 415.540 1369.930 415.680 1462.270 ;
        RECT 414.160 1369.790 415.680 1369.930 ;
        RECT 414.160 1361.770 414.300 1369.790 ;
        RECT 414.160 1361.630 416.140 1361.770 ;
        RECT 416.000 1304.650 416.140 1361.630 ;
        RECT 416.000 1304.510 417.060 1304.650 ;
        RECT 416.920 1265.210 417.060 1304.510 ;
        RECT 416.920 1265.070 417.520 1265.210 ;
        RECT 417.380 1248.890 417.520 1265.070 ;
        RECT 416.460 1248.750 417.520 1248.890 ;
        RECT 416.460 1242.770 416.600 1248.750 ;
        RECT 416.460 1242.630 417.520 1242.770 ;
        RECT 417.380 1183.610 417.520 1242.630 ;
        RECT 417.380 1183.470 417.980 1183.610 ;
        RECT 417.840 1097.250 417.980 1183.470 ;
        RECT 414.620 1097.110 417.980 1097.250 ;
        RECT 414.620 1095.130 414.760 1097.110 ;
        RECT 414.560 1094.810 414.820 1095.130 ;
        RECT 414.620 1038.690 415.680 1038.770 ;
        RECT 414.560 1038.630 415.680 1038.690 ;
        RECT 414.560 1038.370 414.820 1038.630 ;
        RECT 415.540 1035.370 415.680 1038.630 ;
        RECT 415.540 1035.230 416.600 1035.370 ;
        RECT 416.460 965.330 416.600 1035.230 ;
        RECT 416.460 965.190 417.980 965.330 ;
        RECT 417.840 936.090 417.980 965.190 ;
        RECT 414.160 935.950 417.980 936.090 ;
        RECT 414.160 914.330 414.300 935.950 ;
        RECT 414.160 914.190 415.220 914.330 ;
        RECT 415.080 895.290 415.220 914.190 ;
        RECT 415.080 895.150 415.680 895.290 ;
        RECT 415.540 868.770 415.680 895.150 ;
        RECT 415.540 868.630 416.140 868.770 ;
        RECT 416.000 867.410 416.140 868.630 ;
        RECT 415.540 867.270 416.140 867.410 ;
        RECT 414.560 866.730 414.820 866.990 ;
        RECT 415.540 866.730 415.680 867.270 ;
        RECT 414.560 866.670 415.680 866.730 ;
        RECT 414.620 866.590 415.680 866.670 ;
        RECT 414.560 791.930 414.820 792.190 ;
        RECT 414.560 791.870 417.060 791.930 ;
        RECT 414.620 791.790 417.060 791.870 ;
        RECT 416.920 789.890 417.060 791.790 ;
        RECT 416.920 789.750 418.440 789.890 ;
        RECT 414.620 725.210 417.520 725.290 ;
        RECT 414.560 725.150 417.520 725.210 ;
        RECT 414.560 724.890 414.820 725.150 ;
        RECT 417.380 724.610 417.520 725.150 ;
        RECT 418.300 724.610 418.440 789.750 ;
        RECT 417.380 724.470 418.440 724.610 ;
        RECT 414.560 717.810 414.820 718.070 ;
        RECT 414.560 717.750 415.220 717.810 ;
        RECT 414.620 717.670 415.220 717.750 ;
        RECT 415.080 700.810 415.220 717.670 ;
        RECT 414.160 700.670 415.220 700.810 ;
        RECT 414.160 686.530 414.300 700.670 ;
        RECT 413.700 686.390 414.300 686.530 ;
        RECT 413.700 514.070 413.840 686.390 ;
        RECT 413.640 513.750 413.900 514.070 ;
        RECT 1402.640 496.410 1402.900 496.730 ;
        RECT 1402.700 483.210 1402.840 496.410 ;
        RECT 1402.700 483.070 1403.300 483.210 ;
        RECT 1403.160 448.530 1403.300 483.070 ;
        RECT 1402.700 448.390 1403.300 448.530 ;
        RECT 1402.700 434.850 1402.840 448.390 ;
        RECT 1402.640 434.530 1402.900 434.850 ;
        RECT 1402.180 386.250 1402.440 386.570 ;
        RECT 1402.240 386.085 1402.380 386.250 ;
        RECT 1401.250 385.715 1401.530 386.085 ;
        RECT 1402.170 385.715 1402.450 386.085 ;
        RECT 1401.320 352.230 1401.460 385.715 ;
        RECT 1401.260 351.910 1401.520 352.230 ;
        RECT 1401.720 351.570 1401.980 351.890 ;
        RECT 1401.780 303.690 1401.920 351.570 ;
        RECT 1401.780 303.550 1402.380 303.690 ;
        RECT 1402.240 289.670 1402.380 303.550 ;
        RECT 1402.180 289.350 1402.440 289.670 ;
        RECT 1401.720 241.410 1401.980 241.730 ;
        RECT 1401.780 207.130 1401.920 241.410 ;
        RECT 1401.780 206.990 1402.380 207.130 ;
        RECT 1402.240 193.110 1402.380 206.990 ;
        RECT 1402.180 192.790 1402.440 193.110 ;
        RECT 1401.720 158.450 1401.980 158.770 ;
        RECT 1401.780 110.570 1401.920 158.450 ;
        RECT 1401.780 110.430 1402.380 110.570 ;
        RECT 1402.240 62.290 1402.380 110.430 ;
        RECT 1401.320 62.210 1402.380 62.290 ;
        RECT 1401.260 62.150 1402.380 62.210 ;
        RECT 1401.260 61.890 1401.520 62.150 ;
        RECT 1405.860 61.890 1406.120 62.210 ;
        RECT 1401.320 61.735 1401.460 61.890 ;
        RECT 1405.920 61.610 1406.060 61.890 ;
        RECT 1405.920 61.470 1406.520 61.610 ;
        RECT 1406.380 2.400 1406.520 61.470 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
      LAYER via2 ;
        RECT 1401.250 385.760 1401.530 386.040 ;
        RECT 1402.170 385.760 1402.450 386.040 ;
      LAYER met3 ;
        RECT 1401.225 386.050 1401.555 386.065 ;
        RECT 1402.145 386.050 1402.475 386.065 ;
        RECT 1401.225 385.750 1402.475 386.050 ;
        RECT 1401.225 385.735 1401.555 385.750 ;
        RECT 1402.145 385.735 1402.475 385.750 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1131.210 355.540 1131.530 355.600 ;
        RECT 1421.470 355.540 1421.790 355.600 ;
        RECT 1131.210 355.400 1421.790 355.540 ;
        RECT 1131.210 355.340 1131.530 355.400 ;
        RECT 1421.470 355.340 1421.790 355.400 ;
      LAYER via ;
        RECT 1131.240 355.340 1131.500 355.600 ;
        RECT 1421.500 355.340 1421.760 355.600 ;
      LAYER met2 ;
        RECT 1128.610 510.410 1128.890 514.000 ;
        RECT 1128.610 510.270 1131.440 510.410 ;
        RECT 1128.610 510.000 1128.890 510.270 ;
        RECT 1131.300 355.630 1131.440 510.270 ;
        RECT 1131.240 355.310 1131.500 355.630 ;
        RECT 1421.500 355.310 1421.760 355.630 ;
        RECT 1421.560 17.410 1421.700 355.310 ;
        RECT 1421.560 17.270 1424.000 17.410 ;
        RECT 1423.860 2.400 1424.000 17.270 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 391.070 418.100 391.390 418.160 ;
        RECT 1435.270 418.100 1435.590 418.160 ;
        RECT 391.070 417.960 1435.590 418.100 ;
        RECT 391.070 417.900 391.390 417.960 ;
        RECT 1435.270 417.900 1435.590 417.960 ;
        RECT 1435.270 16.900 1435.590 16.960 ;
        RECT 1441.710 16.900 1442.030 16.960 ;
        RECT 1435.270 16.760 1442.030 16.900 ;
        RECT 1435.270 16.700 1435.590 16.760 ;
        RECT 1441.710 16.700 1442.030 16.760 ;
      LAYER via ;
        RECT 391.100 417.900 391.360 418.160 ;
        RECT 1435.300 417.900 1435.560 418.160 ;
        RECT 1435.300 16.700 1435.560 16.960 ;
        RECT 1441.740 16.700 1442.000 16.960 ;
      LAYER met2 ;
        RECT 391.090 1535.595 391.370 1535.965 ;
        RECT 391.160 418.190 391.300 1535.595 ;
        RECT 391.100 417.870 391.360 418.190 ;
        RECT 1435.300 417.870 1435.560 418.190 ;
        RECT 1435.360 16.990 1435.500 417.870 ;
        RECT 1435.300 16.670 1435.560 16.990 ;
        RECT 1441.740 16.670 1442.000 16.990 ;
        RECT 1441.800 2.400 1441.940 16.670 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
      LAYER via2 ;
        RECT 391.090 1535.640 391.370 1535.920 ;
      LAYER met3 ;
        RECT 391.065 1535.930 391.395 1535.945 ;
        RECT 410.000 1535.930 414.000 1536.080 ;
        RECT 391.065 1535.630 414.000 1535.930 ;
        RECT 391.065 1535.615 391.395 1535.630 ;
        RECT 410.000 1535.480 414.000 1535.630 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2408.630 474.880 2408.950 474.940 ;
        RECT 2422.430 474.880 2422.750 474.940 ;
        RECT 2408.630 474.740 2422.750 474.880 ;
        RECT 2408.630 474.680 2408.950 474.740 ;
        RECT 2422.430 474.680 2422.750 474.740 ;
        RECT 2403.570 455.500 2403.890 455.560 ;
        RECT 2408.630 455.500 2408.950 455.560 ;
        RECT 2403.570 455.360 2408.950 455.500 ;
        RECT 2403.570 455.300 2403.890 455.360 ;
        RECT 2408.630 455.300 2408.950 455.360 ;
        RECT 2387.470 427.960 2387.790 428.020 ;
        RECT 2403.570 427.960 2403.890 428.020 ;
        RECT 2387.470 427.820 2403.890 427.960 ;
        RECT 2387.470 427.760 2387.790 427.820 ;
        RECT 2403.570 427.760 2403.890 427.820 ;
        RECT 2366.310 396.680 2366.630 396.740 ;
        RECT 2387.010 396.680 2387.330 396.740 ;
        RECT 2366.310 396.540 2387.330 396.680 ;
        RECT 2366.310 396.480 2366.630 396.540 ;
        RECT 2387.010 396.480 2387.330 396.540 ;
        RECT 2352.970 383.760 2353.290 383.820 ;
        RECT 2366.310 383.760 2366.630 383.820 ;
        RECT 2352.970 383.620 2366.630 383.760 ;
        RECT 2352.970 383.560 2353.290 383.620 ;
        RECT 2366.310 383.560 2366.630 383.620 ;
        RECT 2344.690 345.340 2345.010 345.400 ;
        RECT 2352.510 345.340 2352.830 345.400 ;
        RECT 2344.690 345.200 2352.830 345.340 ;
        RECT 2344.690 345.140 2345.010 345.200 ;
        RECT 2352.510 345.140 2352.830 345.200 ;
        RECT 2335.950 336.160 2336.270 336.220 ;
        RECT 2344.690 336.160 2345.010 336.220 ;
        RECT 2335.950 336.020 2345.010 336.160 ;
        RECT 2335.950 335.960 2336.270 336.020 ;
        RECT 2344.690 335.960 2345.010 336.020 ;
        RECT 2325.830 310.660 2326.150 310.720 ;
        RECT 2335.950 310.660 2336.270 310.720 ;
        RECT 2325.830 310.520 2336.270 310.660 ;
        RECT 2325.830 310.460 2326.150 310.520 ;
        RECT 2335.950 310.460 2336.270 310.520 ;
        RECT 2312.030 289.240 2312.350 289.300 ;
        RECT 2325.830 289.240 2326.150 289.300 ;
        RECT 2312.030 289.100 2326.150 289.240 ;
        RECT 2312.030 289.040 2312.350 289.100 ;
        RECT 2325.830 289.040 2326.150 289.100 ;
        RECT 2307.890 248.440 2308.210 248.500 ;
        RECT 2312.030 248.440 2312.350 248.500 ;
        RECT 2307.890 248.300 2312.350 248.440 ;
        RECT 2307.890 248.240 2308.210 248.300 ;
        RECT 2312.030 248.240 2312.350 248.300 ;
        RECT 2307.890 220.900 2308.210 220.960 ;
        RECT 2297.860 220.760 2308.210 220.900 ;
        RECT 2280.290 220.220 2280.610 220.280 ;
        RECT 2297.860 220.220 2298.000 220.760 ;
        RECT 2307.890 220.700 2308.210 220.760 ;
        RECT 2280.290 220.080 2298.000 220.220 ;
        RECT 2280.290 220.020 2280.610 220.080 ;
        RECT 2262.810 111.080 2263.130 111.140 ;
        RECT 2280.290 111.080 2280.610 111.140 ;
        RECT 2262.810 110.940 2280.610 111.080 ;
        RECT 2262.810 110.880 2263.130 110.940 ;
        RECT 2280.290 110.880 2280.610 110.940 ;
        RECT 2245.790 100.200 2246.110 100.260 ;
        RECT 2262.810 100.200 2263.130 100.260 ;
        RECT 2245.790 100.060 2263.130 100.200 ;
        RECT 2245.790 100.000 2246.110 100.060 ;
        RECT 2262.810 100.000 2263.130 100.060 ;
        RECT 2237.050 38.320 2237.370 38.380 ;
        RECT 2245.790 38.320 2246.110 38.380 ;
        RECT 2237.050 38.180 2246.110 38.320 ;
        RECT 2237.050 38.120 2237.370 38.180 ;
        RECT 2245.790 38.120 2246.110 38.180 ;
        RECT 1459.650 24.720 1459.970 24.780 ;
        RECT 2237.050 24.720 2237.370 24.780 ;
        RECT 1459.650 24.580 2237.370 24.720 ;
        RECT 1459.650 24.520 1459.970 24.580 ;
        RECT 2237.050 24.520 2237.370 24.580 ;
      LAYER via ;
        RECT 2408.660 474.680 2408.920 474.940 ;
        RECT 2422.460 474.680 2422.720 474.940 ;
        RECT 2403.600 455.300 2403.860 455.560 ;
        RECT 2408.660 455.300 2408.920 455.560 ;
        RECT 2387.500 427.760 2387.760 428.020 ;
        RECT 2403.600 427.760 2403.860 428.020 ;
        RECT 2366.340 396.480 2366.600 396.740 ;
        RECT 2387.040 396.480 2387.300 396.740 ;
        RECT 2353.000 383.560 2353.260 383.820 ;
        RECT 2366.340 383.560 2366.600 383.820 ;
        RECT 2344.720 345.140 2344.980 345.400 ;
        RECT 2352.540 345.140 2352.800 345.400 ;
        RECT 2335.980 335.960 2336.240 336.220 ;
        RECT 2344.720 335.960 2344.980 336.220 ;
        RECT 2325.860 310.460 2326.120 310.720 ;
        RECT 2335.980 310.460 2336.240 310.720 ;
        RECT 2312.060 289.040 2312.320 289.300 ;
        RECT 2325.860 289.040 2326.120 289.300 ;
        RECT 2307.920 248.240 2308.180 248.500 ;
        RECT 2312.060 248.240 2312.320 248.500 ;
        RECT 2280.320 220.020 2280.580 220.280 ;
        RECT 2307.920 220.700 2308.180 220.960 ;
        RECT 2262.840 110.880 2263.100 111.140 ;
        RECT 2280.320 110.880 2280.580 111.140 ;
        RECT 2245.820 100.000 2246.080 100.260 ;
        RECT 2262.840 100.000 2263.100 100.260 ;
        RECT 2237.080 38.120 2237.340 38.380 ;
        RECT 2245.820 38.120 2246.080 38.380 ;
        RECT 1459.680 24.520 1459.940 24.780 ;
        RECT 2237.080 24.520 2237.340 24.780 ;
      LAYER met2 ;
        RECT 1469.790 3037.035 1470.070 3037.405 ;
        RECT 1469.860 3010.000 1470.000 3037.035 ;
        RECT 1469.860 3009.340 1470.210 3010.000 ;
        RECT 1469.930 3006.000 1470.210 3009.340 ;
        RECT 2422.450 482.955 2422.730 483.325 ;
        RECT 2422.520 474.970 2422.660 482.955 ;
        RECT 2408.660 474.650 2408.920 474.970 ;
        RECT 2422.460 474.650 2422.720 474.970 ;
        RECT 2408.720 455.590 2408.860 474.650 ;
        RECT 2403.600 455.270 2403.860 455.590 ;
        RECT 2408.660 455.270 2408.920 455.590 ;
        RECT 2403.660 428.050 2403.800 455.270 ;
        RECT 2387.500 427.730 2387.760 428.050 ;
        RECT 2403.600 427.730 2403.860 428.050 ;
        RECT 2387.560 407.730 2387.700 427.730 ;
        RECT 2387.100 407.590 2387.700 407.730 ;
        RECT 2387.100 396.770 2387.240 407.590 ;
        RECT 2366.340 396.450 2366.600 396.770 ;
        RECT 2387.040 396.450 2387.300 396.770 ;
        RECT 2366.400 383.850 2366.540 396.450 ;
        RECT 2353.000 383.530 2353.260 383.850 ;
        RECT 2366.340 383.530 2366.600 383.850 ;
        RECT 2353.060 366.250 2353.200 383.530 ;
        RECT 2352.600 366.110 2353.200 366.250 ;
        RECT 2352.600 345.430 2352.740 366.110 ;
        RECT 2344.720 345.110 2344.980 345.430 ;
        RECT 2352.540 345.110 2352.800 345.430 ;
        RECT 2344.780 336.250 2344.920 345.110 ;
        RECT 2335.980 335.930 2336.240 336.250 ;
        RECT 2344.720 335.930 2344.980 336.250 ;
        RECT 2336.040 310.750 2336.180 335.930 ;
        RECT 2325.860 310.430 2326.120 310.750 ;
        RECT 2335.980 310.430 2336.240 310.750 ;
        RECT 2325.920 289.330 2326.060 310.430 ;
        RECT 2312.060 289.010 2312.320 289.330 ;
        RECT 2325.860 289.010 2326.120 289.330 ;
        RECT 2312.120 248.530 2312.260 289.010 ;
        RECT 2307.920 248.210 2308.180 248.530 ;
        RECT 2312.060 248.210 2312.320 248.530 ;
        RECT 2307.980 220.990 2308.120 248.210 ;
        RECT 2307.920 220.670 2308.180 220.990 ;
        RECT 2280.320 219.990 2280.580 220.310 ;
        RECT 2280.380 111.170 2280.520 219.990 ;
        RECT 2262.840 110.850 2263.100 111.170 ;
        RECT 2280.320 110.850 2280.580 111.170 ;
        RECT 2262.900 100.290 2263.040 110.850 ;
        RECT 2245.820 99.970 2246.080 100.290 ;
        RECT 2262.840 99.970 2263.100 100.290 ;
        RECT 2245.880 38.410 2246.020 99.970 ;
        RECT 2237.080 38.090 2237.340 38.410 ;
        RECT 2245.820 38.090 2246.080 38.410 ;
        RECT 2237.140 24.810 2237.280 38.090 ;
        RECT 1459.680 24.490 1459.940 24.810 ;
        RECT 2237.080 24.490 2237.340 24.810 ;
        RECT 1459.740 2.400 1459.880 24.490 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
      LAYER via2 ;
        RECT 1469.790 3037.080 1470.070 3037.360 ;
        RECT 2422.450 483.000 2422.730 483.280 ;
      LAYER met3 ;
        RECT 1469.765 3037.370 1470.095 3037.385 ;
        RECT 2439.190 3037.370 2439.570 3037.380 ;
        RECT 1469.765 3037.070 2439.570 3037.370 ;
        RECT 1469.765 3037.055 1470.095 3037.070 ;
        RECT 2439.190 3037.060 2439.570 3037.070 ;
        RECT 2439.190 3000.650 2439.570 3000.660 ;
        RECT 2441.030 3000.650 2441.410 3000.660 ;
        RECT 2439.190 3000.350 2441.410 3000.650 ;
        RECT 2439.190 3000.340 2439.570 3000.350 ;
        RECT 2441.030 3000.340 2441.410 3000.350 ;
        RECT 2422.425 483.290 2422.755 483.305 ;
        RECT 2439.190 483.290 2439.570 483.300 ;
        RECT 2422.425 482.990 2439.570 483.290 ;
        RECT 2422.425 482.975 2422.755 482.990 ;
        RECT 2439.190 482.980 2439.570 482.990 ;
      LAYER via3 ;
        RECT 2439.220 3037.060 2439.540 3037.380 ;
        RECT 2439.220 3000.340 2439.540 3000.660 ;
        RECT 2441.060 3000.340 2441.380 3000.660 ;
        RECT 2439.220 482.980 2439.540 483.300 ;
      LAYER met4 ;
        RECT 2439.215 3037.055 2439.545 3037.385 ;
        RECT 2439.230 3000.665 2439.530 3037.055 ;
        RECT 2439.215 3000.335 2439.545 3000.665 ;
        RECT 2441.055 3000.335 2441.385 3000.665 ;
        RECT 2441.070 2980.250 2441.370 3000.335 ;
        RECT 2439.230 2979.950 2441.370 2980.250 ;
        RECT 2439.230 2738.850 2439.530 2979.950 ;
        RECT 2437.390 2738.550 2439.530 2738.850 ;
        RECT 2437.390 2691.250 2437.690 2738.550 ;
        RECT 2437.390 2690.950 2439.530 2691.250 ;
        RECT 2439.230 2256.050 2439.530 2690.950 ;
        RECT 2437.390 2255.750 2439.530 2256.050 ;
        RECT 2437.390 2208.450 2437.690 2255.750 ;
        RECT 2437.390 2208.150 2439.530 2208.450 ;
        RECT 2439.230 2021.450 2439.530 2208.150 ;
        RECT 2439.230 2021.150 2441.370 2021.450 ;
        RECT 2441.070 2007.850 2441.370 2021.150 ;
        RECT 2440.150 2007.550 2441.370 2007.850 ;
        RECT 2440.150 1977.250 2440.450 2007.550 ;
        RECT 2439.230 1976.950 2440.450 1977.250 ;
        RECT 2439.230 1871.850 2439.530 1976.950 ;
        RECT 2438.310 1871.550 2439.530 1871.850 ;
        RECT 2438.310 1831.050 2438.610 1871.550 ;
        RECT 2438.310 1830.750 2439.530 1831.050 ;
        RECT 2439.230 1623.650 2439.530 1830.750 ;
        RECT 2439.230 1623.350 2441.370 1623.650 ;
        RECT 2441.070 1589.650 2441.370 1623.350 ;
        RECT 2439.230 1589.350 2441.370 1589.650 ;
        RECT 2439.230 1545.450 2439.530 1589.350 ;
        RECT 2439.230 1545.150 2441.370 1545.450 ;
        RECT 2441.070 1497.850 2441.370 1545.150 ;
        RECT 2439.230 1497.550 2441.370 1497.850 ;
        RECT 2439.230 1304.050 2439.530 1497.550 ;
        RECT 2438.310 1303.750 2439.530 1304.050 ;
        RECT 2438.310 1256.450 2438.610 1303.750 ;
        RECT 2438.310 1256.150 2439.530 1256.450 ;
        RECT 2439.230 483.305 2439.530 1256.150 ;
        RECT 2439.215 482.975 2439.545 483.305 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2481.330 3006.690 2481.610 3006.805 ;
        RECT 2482.850 3006.690 2483.130 3010.000 ;
        RECT 2481.330 3006.550 2483.130 3006.690 ;
        RECT 2481.330 3006.435 2481.610 3006.550 ;
        RECT 2482.850 3006.000 2483.130 3006.550 ;
        RECT 1477.610 37.555 1477.890 37.925 ;
        RECT 1477.680 2.400 1477.820 37.555 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
      LAYER via2 ;
        RECT 2481.330 3006.480 2481.610 3006.760 ;
        RECT 1477.610 37.600 1477.890 37.880 ;
      LAYER met3 ;
        RECT 2474.150 3006.770 2474.530 3006.780 ;
        RECT 2481.305 3006.770 2481.635 3006.785 ;
        RECT 2474.150 3006.470 2481.635 3006.770 ;
        RECT 2474.150 3006.460 2474.530 3006.470 ;
        RECT 2481.305 3006.455 2481.635 3006.470 ;
        RECT 1477.585 37.890 1477.915 37.905 ;
        RECT 2474.150 37.890 2474.530 37.900 ;
        RECT 1477.585 37.590 2474.530 37.890 ;
        RECT 1477.585 37.575 1477.915 37.590 ;
        RECT 2474.150 37.580 2474.530 37.590 ;
      LAYER via3 ;
        RECT 2474.180 3006.460 2474.500 3006.780 ;
        RECT 2474.180 37.580 2474.500 37.900 ;
      LAYER met4 ;
        RECT 2474.175 3006.455 2474.505 3006.785 ;
        RECT 2474.190 2228.850 2474.490 3006.455 ;
        RECT 2473.270 2228.550 2474.490 2228.850 ;
        RECT 2473.270 2218.650 2473.570 2228.550 ;
        RECT 2473.270 2218.350 2474.490 2218.650 ;
        RECT 2474.190 2143.850 2474.490 2218.350 ;
        RECT 2474.190 2143.550 2476.330 2143.850 ;
        RECT 2476.030 2099.650 2476.330 2143.550 ;
        RECT 2474.190 2099.350 2476.330 2099.650 ;
        RECT 2474.190 1790.690 2474.490 2099.350 ;
        RECT 2473.750 1789.510 2474.930 1790.690 ;
        RECT 2477.430 1789.510 2478.610 1790.690 ;
        RECT 2477.870 1715.450 2478.170 1789.510 ;
        RECT 2476.950 1715.150 2478.170 1715.450 ;
        RECT 2476.950 1640.650 2477.250 1715.150 ;
        RECT 2476.030 1640.350 2477.250 1640.650 ;
        RECT 2476.030 1637.250 2476.330 1640.350 ;
        RECT 2474.190 1636.950 2476.330 1637.250 ;
        RECT 2474.190 1521.650 2474.490 1636.950 ;
        RECT 2474.190 1521.350 2475.410 1521.650 ;
        RECT 2475.110 1511.450 2475.410 1521.350 ;
        RECT 2474.190 1511.150 2475.410 1511.450 ;
        RECT 2474.190 1433.250 2474.490 1511.150 ;
        RECT 2473.270 1432.950 2474.490 1433.250 ;
        RECT 2473.270 1409.890 2473.570 1432.950 ;
        RECT 2472.830 1408.710 2474.010 1409.890 ;
        RECT 2474.670 1401.910 2475.850 1403.090 ;
        RECT 2475.110 1385.650 2475.410 1401.910 ;
        RECT 2474.190 1385.350 2475.410 1385.650 ;
        RECT 2474.190 1335.090 2474.490 1385.350 ;
        RECT 2473.750 1333.910 2474.930 1335.090 ;
        RECT 2481.110 1333.910 2482.290 1335.090 ;
        RECT 2481.550 1321.490 2481.850 1333.910 ;
        RECT 2473.750 1320.310 2474.930 1321.490 ;
        RECT 2481.110 1320.310 2482.290 1321.490 ;
        RECT 2474.190 1293.850 2474.490 1320.310 ;
        RECT 2471.430 1293.550 2474.490 1293.850 ;
        RECT 2471.430 1259.850 2471.730 1293.550 ;
        RECT 2471.430 1259.550 2474.490 1259.850 ;
        RECT 2474.190 1045.650 2474.490 1259.550 ;
        RECT 2474.190 1045.350 2476.330 1045.650 ;
        RECT 2476.030 981.050 2476.330 1045.350 ;
        RECT 2474.190 980.750 2476.330 981.050 ;
        RECT 2474.190 885.850 2474.490 980.750 ;
        RECT 2474.190 885.550 2476.330 885.850 ;
        RECT 2476.030 879.050 2476.330 885.550 ;
        RECT 2474.190 878.750 2476.330 879.050 ;
        RECT 2474.190 828.490 2474.490 878.750 ;
        RECT 2465.470 827.310 2466.650 828.490 ;
        RECT 2473.750 827.310 2474.930 828.490 ;
        RECT 2465.910 780.890 2466.210 827.310 ;
        RECT 2465.470 779.710 2466.650 780.890 ;
        RECT 2474.670 779.710 2475.850 780.890 ;
        RECT 2475.110 773.650 2475.410 779.710 ;
        RECT 2474.190 773.350 2475.410 773.650 ;
        RECT 2474.190 654.650 2474.490 773.350 ;
        RECT 2474.190 654.350 2477.250 654.650 ;
        RECT 2476.950 603.650 2477.250 654.350 ;
        RECT 2474.190 603.350 2477.250 603.650 ;
        RECT 2474.190 600.250 2474.490 603.350 ;
        RECT 2473.270 599.950 2474.490 600.250 ;
        RECT 2473.270 552.650 2473.570 599.950 ;
        RECT 2473.270 552.350 2474.490 552.650 ;
        RECT 2474.190 37.905 2474.490 552.350 ;
        RECT 2474.175 37.575 2474.505 37.905 ;
      LAYER met5 ;
        RECT 2473.540 1789.300 2478.820 1790.900 ;
        RECT 2472.620 1403.300 2474.220 1410.100 ;
        RECT 2472.620 1401.700 2476.060 1403.300 ;
        RECT 2473.540 1333.700 2482.500 1335.300 ;
        RECT 2473.540 1320.100 2482.500 1321.700 ;
        RECT 2465.260 827.100 2475.140 828.700 ;
        RECT 2465.260 779.500 2476.060 781.100 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 410.850 3011.280 411.170 3011.340 ;
        RECT 715.370 3011.280 715.690 3011.340 ;
        RECT 410.850 3011.140 715.690 3011.280 ;
        RECT 410.850 3011.080 411.170 3011.140 ;
        RECT 715.370 3011.080 715.690 3011.140 ;
        RECT 348.290 776.120 348.610 776.180 ;
        RECT 410.850 776.120 411.170 776.180 ;
        RECT 348.290 775.980 411.170 776.120 ;
        RECT 348.290 775.920 348.610 775.980 ;
        RECT 410.850 775.920 411.170 775.980 ;
      LAYER via ;
        RECT 410.880 3011.080 411.140 3011.340 ;
        RECT 715.400 3011.080 715.660 3011.340 ;
        RECT 348.320 775.920 348.580 776.180 ;
        RECT 410.880 775.920 411.140 776.180 ;
      LAYER met2 ;
        RECT 410.880 3011.050 411.140 3011.370 ;
        RECT 715.400 3011.050 715.660 3011.370 ;
        RECT 410.940 776.210 411.080 3011.050 ;
        RECT 715.460 3010.000 715.600 3011.050 ;
        RECT 715.460 3009.340 715.810 3010.000 ;
        RECT 715.530 3006.000 715.810 3009.340 ;
        RECT 348.320 775.890 348.580 776.210 ;
        RECT 410.880 775.890 411.140 776.210 ;
        RECT 348.380 19.565 348.520 775.890 ;
        RECT 348.310 19.195 348.590 19.565 ;
        RECT 366.250 19.195 366.530 19.565 ;
        RECT 366.320 17.525 366.460 19.195 ;
        RECT 366.250 17.155 366.530 17.525 ;
        RECT 1495.550 17.155 1495.830 17.525 ;
        RECT 1495.620 2.400 1495.760 17.155 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
      LAYER via2 ;
        RECT 348.310 19.240 348.590 19.520 ;
        RECT 366.250 19.240 366.530 19.520 ;
        RECT 366.250 17.200 366.530 17.480 ;
        RECT 1495.550 17.200 1495.830 17.480 ;
      LAYER met3 ;
        RECT 348.285 19.530 348.615 19.545 ;
        RECT 366.225 19.530 366.555 19.545 ;
        RECT 348.285 19.230 366.555 19.530 ;
        RECT 348.285 19.215 348.615 19.230 ;
        RECT 366.225 19.215 366.555 19.230 ;
        RECT 366.225 17.490 366.555 17.505 ;
        RECT 1495.525 17.490 1495.855 17.505 ;
        RECT 366.225 17.190 1495.855 17.490 ;
        RECT 366.225 17.175 366.555 17.190 ;
        RECT 1495.525 17.175 1495.855 17.190 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.250 510.410 1512.530 514.000 ;
        RECT 1511.260 510.270 1512.530 510.410 ;
        RECT 1511.260 17.410 1511.400 510.270 ;
        RECT 1512.250 510.000 1512.530 510.270 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 328.510 890.360 328.830 890.420 ;
        RECT 393.370 890.360 393.690 890.420 ;
        RECT 328.510 890.220 393.690 890.360 ;
        RECT 328.510 890.160 328.830 890.220 ;
        RECT 393.370 890.160 393.690 890.220 ;
        RECT 328.510 62.120 328.830 62.180 ;
        RECT 710.310 62.120 710.630 62.180 ;
        RECT 328.510 61.980 710.630 62.120 ;
        RECT 328.510 61.920 328.830 61.980 ;
        RECT 710.310 61.920 710.630 61.980 ;
      LAYER via ;
        RECT 328.540 890.160 328.800 890.420 ;
        RECT 393.400 890.160 393.660 890.420 ;
        RECT 328.540 61.920 328.800 62.180 ;
        RECT 710.340 61.920 710.600 62.180 ;
      LAYER met2 ;
        RECT 393.390 896.395 393.670 896.765 ;
        RECT 393.460 890.450 393.600 896.395 ;
        RECT 328.540 890.130 328.800 890.450 ;
        RECT 393.400 890.130 393.660 890.450 ;
        RECT 328.600 62.210 328.740 890.130 ;
        RECT 328.540 61.890 328.800 62.210 ;
        RECT 710.340 61.890 710.600 62.210 ;
        RECT 710.400 2.400 710.540 61.890 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 393.390 896.440 393.670 896.720 ;
      LAYER met3 ;
        RECT 393.365 896.730 393.695 896.745 ;
        RECT 410.000 896.730 414.000 896.880 ;
        RECT 393.365 896.430 414.000 896.730 ;
        RECT 393.365 896.415 393.695 896.430 ;
        RECT 410.000 896.280 414.000 896.430 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 390.610 445.300 390.930 445.360 ;
        RECT 1524.970 445.300 1525.290 445.360 ;
        RECT 390.610 445.160 1525.290 445.300 ;
        RECT 390.610 445.100 390.930 445.160 ;
        RECT 1524.970 445.100 1525.290 445.160 ;
        RECT 1524.970 16.900 1525.290 16.960 ;
        RECT 1530.950 16.900 1531.270 16.960 ;
        RECT 1524.970 16.760 1531.270 16.900 ;
        RECT 1524.970 16.700 1525.290 16.760 ;
        RECT 1530.950 16.700 1531.270 16.760 ;
      LAYER via ;
        RECT 390.640 445.100 390.900 445.360 ;
        RECT 1525.000 445.100 1525.260 445.360 ;
        RECT 1525.000 16.700 1525.260 16.960 ;
        RECT 1530.980 16.700 1531.240 16.960 ;
      LAYER met2 ;
        RECT 390.630 1517.915 390.910 1518.285 ;
        RECT 390.700 445.390 390.840 1517.915 ;
        RECT 390.640 445.070 390.900 445.390 ;
        RECT 1525.000 445.070 1525.260 445.390 ;
        RECT 1525.060 16.990 1525.200 445.070 ;
        RECT 1525.000 16.670 1525.260 16.990 ;
        RECT 1530.980 16.670 1531.240 16.990 ;
        RECT 1531.040 2.400 1531.180 16.670 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
      LAYER via2 ;
        RECT 390.630 1517.960 390.910 1518.240 ;
      LAYER met3 ;
        RECT 390.605 1518.250 390.935 1518.265 ;
        RECT 410.000 1518.250 414.000 1518.400 ;
        RECT 390.605 1517.950 414.000 1518.250 ;
        RECT 390.605 1517.935 390.935 1517.950 ;
        RECT 410.000 1517.800 414.000 1517.950 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1545.690 472.075 1545.970 472.445 ;
        RECT 1545.760 17.410 1545.900 472.075 ;
        RECT 1545.760 17.270 1549.120 17.410 ;
        RECT 1548.980 2.400 1549.120 17.270 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
      LAYER via2 ;
        RECT 1545.690 472.120 1545.970 472.400 ;
      LAYER met3 ;
        RECT 391.270 2742.250 391.650 2742.260 ;
        RECT 410.000 2742.250 414.000 2742.400 ;
        RECT 391.270 2741.950 414.000 2742.250 ;
        RECT 391.270 2741.940 391.650 2741.950 ;
        RECT 410.000 2741.800 414.000 2741.950 ;
        RECT 391.270 472.410 391.650 472.420 ;
        RECT 1545.665 472.410 1545.995 472.425 ;
        RECT 391.270 472.110 1545.995 472.410 ;
        RECT 391.270 472.100 391.650 472.110 ;
        RECT 1545.665 472.095 1545.995 472.110 ;
      LAYER via3 ;
        RECT 391.300 2741.940 391.620 2742.260 ;
        RECT 391.300 472.100 391.620 472.420 ;
      LAYER met4 ;
        RECT 391.295 2741.935 391.625 2742.265 ;
        RECT 391.310 472.425 391.610 2741.935 ;
        RECT 391.295 472.095 391.625 472.425 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.510 32.540 1317.830 32.600 ;
        RECT 1566.830 32.540 1567.150 32.600 ;
        RECT 1317.510 32.400 1567.150 32.540 ;
        RECT 1317.510 32.340 1317.830 32.400 ;
        RECT 1566.830 32.340 1567.150 32.400 ;
      LAYER via ;
        RECT 1317.540 32.340 1317.800 32.600 ;
        RECT 1566.860 32.340 1567.120 32.600 ;
      LAYER met2 ;
        RECT 1314.450 510.410 1314.730 514.000 ;
        RECT 1314.450 510.270 1317.740 510.410 ;
        RECT 1314.450 510.000 1314.730 510.270 ;
        RECT 1317.600 32.630 1317.740 510.270 ;
        RECT 1317.540 32.310 1317.800 32.630 ;
        RECT 1566.860 32.310 1567.120 32.630 ;
        RECT 1566.920 2.400 1567.060 32.310 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1586.630 258.555 1586.910 258.925 ;
        RECT 1586.700 17.410 1586.840 258.555 ;
        RECT 1584.860 17.270 1586.840 17.410 ;
        RECT 1584.860 2.400 1585.000 17.270 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 1586.630 258.600 1586.910 258.880 ;
      LAYER met3 ;
        RECT 2506.000 2549.130 2510.000 2549.280 ;
        RECT 2513.710 2549.130 2514.090 2549.140 ;
        RECT 2506.000 2548.830 2514.090 2549.130 ;
        RECT 2506.000 2548.680 2510.000 2548.830 ;
        RECT 2513.710 2548.820 2514.090 2548.830 ;
        RECT 1586.605 258.890 1586.935 258.905 ;
        RECT 2513.710 258.890 2514.090 258.900 ;
        RECT 1586.605 258.590 2514.090 258.890 ;
        RECT 1586.605 258.575 1586.935 258.590 ;
        RECT 2513.710 258.580 2514.090 258.590 ;
      LAYER via3 ;
        RECT 2513.740 2548.820 2514.060 2549.140 ;
        RECT 2513.740 258.580 2514.060 258.900 ;
      LAYER met4 ;
        RECT 2513.735 2548.815 2514.065 2549.145 ;
        RECT 2513.750 258.905 2514.050 2548.815 ;
        RECT 2513.735 258.575 2514.065 258.905 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 408.550 341.940 408.870 342.000 ;
        RECT 1600.870 341.940 1601.190 342.000 ;
        RECT 408.550 341.800 1601.190 341.940 ;
        RECT 408.550 341.740 408.870 341.800 ;
        RECT 1600.870 341.740 1601.190 341.800 ;
      LAYER via ;
        RECT 408.580 341.740 408.840 342.000 ;
        RECT 1600.900 341.740 1601.160 342.000 ;
      LAYER met2 ;
        RECT 408.570 1079.995 408.850 1080.365 ;
        RECT 408.640 342.030 408.780 1079.995 ;
        RECT 408.580 341.710 408.840 342.030 ;
        RECT 1600.900 341.710 1601.160 342.030 ;
        RECT 1600.960 17.410 1601.100 341.710 ;
        RECT 1600.960 17.270 1602.480 17.410 ;
        RECT 1602.340 2.400 1602.480 17.270 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
      LAYER via2 ;
        RECT 408.570 1080.040 408.850 1080.320 ;
      LAYER met3 ;
        RECT 408.545 1080.330 408.875 1080.345 ;
        RECT 410.000 1080.330 414.000 1080.480 ;
        RECT 408.545 1080.030 414.000 1080.330 ;
        RECT 408.545 1080.015 408.875 1080.030 ;
        RECT 410.000 1079.880 414.000 1080.030 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2173.730 3006.690 2174.010 3010.000 ;
        RECT 2175.430 3006.690 2175.710 3006.805 ;
        RECT 2173.730 3006.550 2175.710 3006.690 ;
        RECT 2173.730 3006.000 2174.010 3006.550 ;
        RECT 2175.430 3006.435 2175.710 3006.550 ;
        RECT 1621.130 508.795 1621.410 509.165 ;
        RECT 1621.200 17.410 1621.340 508.795 ;
        RECT 1620.280 17.270 1621.340 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
      LAYER via2 ;
        RECT 2175.430 3006.480 2175.710 3006.760 ;
        RECT 1621.130 508.840 1621.410 509.120 ;
      LAYER met3 ;
        RECT 2175.405 3006.770 2175.735 3006.785 ;
        RECT 2175.405 3006.470 2181.010 3006.770 ;
        RECT 2175.405 3006.455 2175.735 3006.470 ;
        RECT 2180.710 3004.730 2181.010 3006.470 ;
        RECT 2487.950 3004.730 2488.330 3004.740 ;
        RECT 2180.710 3004.430 2488.330 3004.730 ;
        RECT 2487.950 3004.420 2488.330 3004.430 ;
        RECT 1621.105 509.130 1621.435 509.145 ;
        RECT 2445.630 509.130 2446.010 509.140 ;
        RECT 1621.105 508.830 2446.010 509.130 ;
        RECT 1621.105 508.815 1621.435 508.830 ;
        RECT 2445.630 508.820 2446.010 508.830 ;
      LAYER via3 ;
        RECT 2487.980 3004.420 2488.300 3004.740 ;
        RECT 2445.660 508.820 2445.980 509.140 ;
      LAYER met4 ;
        RECT 2487.975 3004.415 2488.305 3004.745 ;
        RECT 2487.990 2925.850 2488.290 3004.415 ;
        RECT 2486.150 2925.550 2488.290 2925.850 ;
        RECT 2486.150 2897.970 2486.450 2925.550 ;
        RECT 2486.150 2897.670 2488.290 2897.970 ;
        RECT 2487.990 2864.650 2488.290 2897.670 ;
        RECT 2487.990 2864.350 2491.050 2864.650 ;
        RECT 2490.750 2830.650 2491.050 2864.350 ;
        RECT 2489.830 2830.350 2491.050 2830.650 ;
        RECT 2489.830 2823.850 2490.130 2830.350 ;
        RECT 2486.150 2823.550 2490.130 2823.850 ;
        RECT 2486.150 2718.450 2486.450 2823.550 ;
        RECT 2486.150 2718.150 2488.290 2718.450 ;
        RECT 2487.990 2711.650 2488.290 2718.150 ;
        RECT 2487.990 2711.350 2490.130 2711.650 ;
        RECT 2489.830 2667.450 2490.130 2711.350 ;
        RECT 2487.990 2667.150 2490.130 2667.450 ;
        RECT 2487.990 2565.450 2488.290 2667.150 ;
        RECT 2486.150 2565.150 2488.290 2565.450 ;
        RECT 2486.150 2470.250 2486.450 2565.150 ;
        RECT 2485.230 2469.950 2486.450 2470.250 ;
        RECT 2485.230 2415.850 2485.530 2469.950 ;
        RECT 2485.230 2415.550 2486.450 2415.850 ;
        RECT 2486.150 2392.050 2486.450 2415.550 ;
        RECT 2486.150 2391.750 2488.290 2392.050 ;
        RECT 2487.990 2375.050 2488.290 2391.750 ;
        RECT 2487.990 2374.750 2491.050 2375.050 ;
        RECT 2487.990 2323.750 2490.130 2324.050 ;
        RECT 2487.990 2262.850 2488.290 2323.750 ;
        RECT 2489.830 2320.650 2490.130 2323.750 ;
        RECT 2490.750 2320.650 2491.050 2374.750 ;
        RECT 2489.830 2320.350 2491.050 2320.650 ;
        RECT 2487.070 2262.550 2488.290 2262.850 ;
        RECT 2487.070 2252.650 2487.370 2262.550 ;
        RECT 2487.070 2252.350 2488.290 2252.650 ;
        RECT 2487.990 2242.450 2488.290 2252.350 ;
        RECT 2487.070 2242.150 2488.290 2242.450 ;
        RECT 2487.070 2239.050 2487.370 2242.150 ;
        RECT 2486.150 2238.750 2487.370 2239.050 ;
        RECT 2486.150 2184.650 2486.450 2238.750 ;
        RECT 2486.150 2184.350 2487.370 2184.650 ;
        RECT 2487.070 2150.650 2487.370 2184.350 ;
        RECT 2486.150 2150.350 2487.370 2150.650 ;
        RECT 2486.150 2109.850 2486.450 2150.350 ;
        RECT 2486.150 2109.550 2487.370 2109.850 ;
        RECT 2487.070 2106.450 2487.370 2109.550 ;
        RECT 2487.070 2106.150 2489.210 2106.450 ;
        RECT 2488.910 2018.490 2489.210 2106.150 ;
        RECT 2488.470 2017.310 2489.650 2018.490 ;
        RECT 2486.630 2013.910 2487.810 2015.090 ;
        RECT 2487.070 1960.250 2487.370 2013.910 ;
        RECT 2486.150 1959.950 2487.370 1960.250 ;
        RECT 2486.150 1950.490 2486.450 1959.950 ;
        RECT 2485.710 1949.310 2486.890 1950.490 ;
        RECT 2493.070 1949.310 2494.250 1950.490 ;
        RECT 2493.510 1909.690 2493.810 1949.310 ;
        RECT 2493.070 1908.510 2494.250 1909.690 ;
        RECT 2485.710 1905.110 2486.890 1906.290 ;
        RECT 2486.150 1892.690 2486.450 1905.110 ;
        RECT 2445.230 1891.510 2446.410 1892.690 ;
        RECT 2485.710 1891.510 2486.890 1892.690 ;
        RECT 2445.670 509.145 2445.970 1891.510 ;
        RECT 2445.655 508.815 2445.985 509.145 ;
      LAYER met5 ;
        RECT 2485.500 2017.100 2489.860 2018.700 ;
        RECT 2485.500 2015.300 2487.100 2017.100 ;
        RECT 2485.500 2013.700 2488.020 2015.300 ;
        RECT 2485.500 1949.100 2494.460 1950.700 ;
        RECT 2485.500 1908.300 2494.460 1909.900 ;
        RECT 2485.500 1904.900 2487.100 1908.300 ;
        RECT 2445.020 1891.300 2487.100 1892.900 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 3036.440 1766.330 3036.500 ;
        RECT 2524.090 3036.440 2524.410 3036.500 ;
        RECT 1766.010 3036.300 2524.410 3036.440 ;
        RECT 1766.010 3036.240 1766.330 3036.300 ;
        RECT 2524.090 3036.240 2524.410 3036.300 ;
        RECT 2524.090 3006.860 2524.410 3006.920 ;
        RECT 2536.510 3006.860 2536.830 3006.920 ;
        RECT 2524.090 3006.720 2536.830 3006.860 ;
        RECT 2524.090 3006.660 2524.410 3006.720 ;
        RECT 2536.510 3006.660 2536.830 3006.720 ;
        RECT 2536.510 2935.800 2536.830 2935.860 ;
        RECT 2616.090 2935.800 2616.410 2935.860 ;
        RECT 2536.510 2935.660 2616.410 2935.800 ;
        RECT 2536.510 2935.600 2536.830 2935.660 ;
        RECT 2616.090 2935.600 2616.410 2935.660 ;
        RECT 2438.990 487.800 2439.310 487.860 ;
        RECT 2616.090 487.800 2616.410 487.860 ;
        RECT 2438.990 487.660 2616.410 487.800 ;
        RECT 2438.990 487.600 2439.310 487.660 ;
        RECT 2616.090 487.600 2616.410 487.660 ;
        RECT 2421.050 475.220 2421.370 475.280 ;
        RECT 2438.990 475.220 2439.310 475.280 ;
        RECT 2421.050 475.080 2439.310 475.220 ;
        RECT 2421.050 475.020 2421.370 475.080 ;
        RECT 2438.990 475.020 2439.310 475.080 ;
        RECT 2411.390 442.580 2411.710 442.640 ;
        RECT 2421.050 442.580 2421.370 442.640 ;
        RECT 2411.390 442.440 2421.370 442.580 ;
        RECT 2411.390 442.380 2411.710 442.440 ;
        RECT 2421.050 442.380 2421.370 442.440 ;
        RECT 2404.490 379.340 2404.810 379.400 ;
        RECT 2411.390 379.340 2411.710 379.400 ;
        RECT 2404.490 379.200 2411.710 379.340 ;
        RECT 2404.490 379.140 2404.810 379.200 ;
        RECT 2411.390 379.140 2411.710 379.200 ;
        RECT 2383.790 313.380 2384.110 313.440 ;
        RECT 2404.490 313.380 2404.810 313.440 ;
        RECT 2383.790 313.240 2404.810 313.380 ;
        RECT 2383.790 313.180 2384.110 313.240 ;
        RECT 2404.490 313.180 2404.810 313.240 ;
        RECT 2369.990 262.380 2370.310 262.440 ;
        RECT 2383.790 262.380 2384.110 262.440 ;
        RECT 2369.990 262.240 2384.110 262.380 ;
        RECT 2369.990 262.180 2370.310 262.240 ;
        RECT 2383.790 262.180 2384.110 262.240 ;
        RECT 2346.530 210.360 2346.850 210.420 ;
        RECT 2369.990 210.360 2370.310 210.420 ;
        RECT 2346.530 210.220 2370.310 210.360 ;
        RECT 2346.530 210.160 2346.850 210.220 ;
        RECT 2369.990 210.160 2370.310 210.220 ;
        RECT 2328.590 200.500 2328.910 200.560 ;
        RECT 2346.530 200.500 2346.850 200.560 ;
        RECT 2328.590 200.360 2346.850 200.500 ;
        RECT 2328.590 200.300 2328.910 200.360 ;
        RECT 2346.530 200.300 2346.850 200.360 ;
        RECT 2314.790 172.620 2315.110 172.680 ;
        RECT 2328.590 172.620 2328.910 172.680 ;
        RECT 2314.790 172.480 2328.910 172.620 ;
        RECT 2314.790 172.420 2315.110 172.480 ;
        RECT 2328.590 172.420 2328.910 172.480 ;
        RECT 2287.190 54.980 2287.510 55.040 ;
        RECT 2314.790 54.980 2315.110 55.040 ;
        RECT 2287.190 54.840 2315.110 54.980 ;
        RECT 2287.190 54.780 2287.510 54.840 ;
        RECT 2314.790 54.780 2315.110 54.840 ;
        RECT 1638.130 25.060 1638.450 25.120 ;
        RECT 2287.190 25.060 2287.510 25.120 ;
        RECT 1638.130 24.920 2287.510 25.060 ;
        RECT 1638.130 24.860 1638.450 24.920 ;
        RECT 2287.190 24.860 2287.510 24.920 ;
      LAYER via ;
        RECT 1766.040 3036.240 1766.300 3036.500 ;
        RECT 2524.120 3036.240 2524.380 3036.500 ;
        RECT 2524.120 3006.660 2524.380 3006.920 ;
        RECT 2536.540 3006.660 2536.800 3006.920 ;
        RECT 2536.540 2935.600 2536.800 2935.860 ;
        RECT 2616.120 2935.600 2616.380 2935.860 ;
        RECT 2439.020 487.600 2439.280 487.860 ;
        RECT 2616.120 487.600 2616.380 487.860 ;
        RECT 2421.080 475.020 2421.340 475.280 ;
        RECT 2439.020 475.020 2439.280 475.280 ;
        RECT 2411.420 442.380 2411.680 442.640 ;
        RECT 2421.080 442.380 2421.340 442.640 ;
        RECT 2404.520 379.140 2404.780 379.400 ;
        RECT 2411.420 379.140 2411.680 379.400 ;
        RECT 2383.820 313.180 2384.080 313.440 ;
        RECT 2404.520 313.180 2404.780 313.440 ;
        RECT 2370.020 262.180 2370.280 262.440 ;
        RECT 2383.820 262.180 2384.080 262.440 ;
        RECT 2346.560 210.160 2346.820 210.420 ;
        RECT 2370.020 210.160 2370.280 210.420 ;
        RECT 2328.620 200.300 2328.880 200.560 ;
        RECT 2346.560 200.300 2346.820 200.560 ;
        RECT 2314.820 172.420 2315.080 172.680 ;
        RECT 2328.620 172.420 2328.880 172.680 ;
        RECT 2287.220 54.780 2287.480 55.040 ;
        RECT 2314.820 54.780 2315.080 55.040 ;
        RECT 1638.160 24.860 1638.420 25.120 ;
        RECT 2287.220 24.860 2287.480 25.120 ;
      LAYER met2 ;
        RECT 1766.040 3036.210 1766.300 3036.530 ;
        RECT 2524.120 3036.210 2524.380 3036.530 ;
        RECT 1766.100 3010.000 1766.240 3036.210 ;
        RECT 1766.100 3009.340 1766.450 3010.000 ;
        RECT 1766.170 3006.000 1766.450 3009.340 ;
        RECT 2524.180 3006.950 2524.320 3036.210 ;
        RECT 2524.120 3006.630 2524.380 3006.950 ;
        RECT 2536.540 3006.630 2536.800 3006.950 ;
        RECT 2536.600 2935.890 2536.740 3006.630 ;
        RECT 2536.540 2935.570 2536.800 2935.890 ;
        RECT 2616.120 2935.570 2616.380 2935.890 ;
        RECT 2616.180 487.890 2616.320 2935.570 ;
        RECT 2439.020 487.570 2439.280 487.890 ;
        RECT 2616.120 487.570 2616.380 487.890 ;
        RECT 2439.080 475.310 2439.220 487.570 ;
        RECT 2421.080 474.990 2421.340 475.310 ;
        RECT 2439.020 474.990 2439.280 475.310 ;
        RECT 2421.140 442.670 2421.280 474.990 ;
        RECT 2411.420 442.350 2411.680 442.670 ;
        RECT 2421.080 442.350 2421.340 442.670 ;
        RECT 2411.480 379.430 2411.620 442.350 ;
        RECT 2404.520 379.110 2404.780 379.430 ;
        RECT 2411.420 379.110 2411.680 379.430 ;
        RECT 2404.580 313.470 2404.720 379.110 ;
        RECT 2383.820 313.150 2384.080 313.470 ;
        RECT 2404.520 313.150 2404.780 313.470 ;
        RECT 2383.880 262.470 2384.020 313.150 ;
        RECT 2370.020 262.150 2370.280 262.470 ;
        RECT 2383.820 262.150 2384.080 262.470 ;
        RECT 2370.080 210.450 2370.220 262.150 ;
        RECT 2346.560 210.130 2346.820 210.450 ;
        RECT 2370.020 210.130 2370.280 210.450 ;
        RECT 2346.620 200.590 2346.760 210.130 ;
        RECT 2328.620 200.270 2328.880 200.590 ;
        RECT 2346.560 200.270 2346.820 200.590 ;
        RECT 2328.680 172.710 2328.820 200.270 ;
        RECT 2314.820 172.390 2315.080 172.710 ;
        RECT 2328.620 172.390 2328.880 172.710 ;
        RECT 2314.880 55.070 2315.020 172.390 ;
        RECT 2287.220 54.750 2287.480 55.070 ;
        RECT 2314.820 54.750 2315.080 55.070 ;
        RECT 2287.280 25.150 2287.420 54.750 ;
        RECT 1638.160 24.830 1638.420 25.150 ;
        RECT 2287.220 24.830 2287.480 25.150 ;
        RECT 1638.220 2.400 1638.360 24.830 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 369.480 1662.830 369.540 ;
        RECT 2508.450 369.480 2508.770 369.540 ;
        RECT 1662.510 369.340 2508.770 369.480 ;
        RECT 1662.510 369.280 1662.830 369.340 ;
        RECT 2508.450 369.280 2508.770 369.340 ;
        RECT 1656.070 20.300 1656.390 20.360 ;
        RECT 1662.510 20.300 1662.830 20.360 ;
        RECT 1656.070 20.160 1662.830 20.300 ;
        RECT 1656.070 20.100 1656.390 20.160 ;
        RECT 1662.510 20.100 1662.830 20.160 ;
      LAYER via ;
        RECT 1662.540 369.280 1662.800 369.540 ;
        RECT 2508.480 369.280 2508.740 369.540 ;
        RECT 1656.100 20.100 1656.360 20.360 ;
        RECT 1662.540 20.100 1662.800 20.360 ;
      LAYER met2 ;
        RECT 2508.470 1359.475 2508.750 1359.845 ;
        RECT 2508.540 369.570 2508.680 1359.475 ;
        RECT 1662.540 369.250 1662.800 369.570 ;
        RECT 2508.480 369.250 2508.740 369.570 ;
        RECT 1662.600 20.390 1662.740 369.250 ;
        RECT 1656.100 20.070 1656.360 20.390 ;
        RECT 1662.540 20.070 1662.800 20.390 ;
        RECT 1656.160 2.400 1656.300 20.070 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
      LAYER via2 ;
        RECT 2508.470 1359.520 2508.750 1359.800 ;
      LAYER met3 ;
        RECT 2506.000 1361.400 2510.000 1362.000 ;
        RECT 2508.230 1359.825 2508.530 1361.400 ;
        RECT 2508.230 1359.510 2508.775 1359.825 ;
        RECT 2508.445 1359.495 2508.775 1359.510 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1400.770 502.420 1401.090 502.480 ;
        RECT 1407.210 502.420 1407.530 502.480 ;
        RECT 1400.770 502.280 1407.530 502.420 ;
        RECT 1400.770 502.220 1401.090 502.280 ;
        RECT 1407.210 502.220 1407.530 502.280 ;
        RECT 1407.210 231.440 1407.530 231.500 ;
        RECT 1669.870 231.440 1670.190 231.500 ;
        RECT 1407.210 231.300 1670.190 231.440 ;
        RECT 1407.210 231.240 1407.530 231.300 ;
        RECT 1669.870 231.240 1670.190 231.300 ;
        RECT 1669.870 96.460 1670.190 96.520 ;
        RECT 1674.010 96.460 1674.330 96.520 ;
        RECT 1669.870 96.320 1674.330 96.460 ;
        RECT 1669.870 96.260 1670.190 96.320 ;
        RECT 1674.010 96.260 1674.330 96.320 ;
      LAYER via ;
        RECT 1400.800 502.220 1401.060 502.480 ;
        RECT 1407.240 502.220 1407.500 502.480 ;
        RECT 1407.240 231.240 1407.500 231.500 ;
        RECT 1669.900 231.240 1670.160 231.500 ;
        RECT 1669.900 96.260 1670.160 96.520 ;
        RECT 1674.040 96.260 1674.300 96.520 ;
      LAYER met2 ;
        RECT 1400.930 510.340 1401.210 514.000 ;
        RECT 1400.860 510.000 1401.210 510.340 ;
        RECT 1400.860 502.510 1401.000 510.000 ;
        RECT 1400.800 502.190 1401.060 502.510 ;
        RECT 1407.240 502.190 1407.500 502.510 ;
        RECT 1407.300 231.530 1407.440 502.190 ;
        RECT 1407.240 231.210 1407.500 231.530 ;
        RECT 1669.900 231.210 1670.160 231.530 ;
        RECT 1669.960 96.550 1670.100 231.210 ;
        RECT 1669.900 96.230 1670.160 96.550 ;
        RECT 1674.040 96.230 1674.300 96.550 ;
        RECT 1674.100 15.880 1674.240 96.230 ;
        RECT 1673.640 15.740 1674.240 15.880 ;
        RECT 1673.640 2.400 1673.780 15.740 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1690.645 48.365 1690.815 96.475 ;
      LAYER mcon ;
        RECT 1690.645 96.305 1690.815 96.475 ;
      LAYER met1 ;
        RECT 397.970 100.200 398.290 100.260 ;
        RECT 1691.030 100.200 1691.350 100.260 ;
        RECT 397.970 100.060 1691.350 100.200 ;
        RECT 397.970 100.000 398.290 100.060 ;
        RECT 1691.030 100.000 1691.350 100.060 ;
        RECT 1690.570 96.460 1690.890 96.520 ;
        RECT 1690.570 96.320 1691.085 96.460 ;
        RECT 1690.570 96.260 1690.890 96.320 ;
        RECT 1690.585 48.520 1690.875 48.565 ;
        RECT 1691.490 48.520 1691.810 48.580 ;
        RECT 1690.585 48.380 1691.810 48.520 ;
        RECT 1690.585 48.335 1690.875 48.380 ;
        RECT 1691.490 48.320 1691.810 48.380 ;
      LAYER via ;
        RECT 398.000 100.000 398.260 100.260 ;
        RECT 1691.060 100.000 1691.320 100.260 ;
        RECT 1690.600 96.260 1690.860 96.520 ;
        RECT 1691.520 48.320 1691.780 48.580 ;
      LAYER met2 ;
        RECT 397.990 1097.675 398.270 1098.045 ;
        RECT 398.060 100.290 398.200 1097.675 ;
        RECT 398.000 99.970 398.260 100.290 ;
        RECT 1691.060 99.970 1691.320 100.290 ;
        RECT 1691.120 96.970 1691.260 99.970 ;
        RECT 1690.660 96.830 1691.260 96.970 ;
        RECT 1690.660 96.550 1690.800 96.830 ;
        RECT 1690.600 96.230 1690.860 96.550 ;
        RECT 1691.520 48.290 1691.780 48.610 ;
        RECT 1691.580 2.400 1691.720 48.290 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
      LAYER via2 ;
        RECT 397.990 1097.720 398.270 1098.000 ;
      LAYER met3 ;
        RECT 397.965 1098.010 398.295 1098.025 ;
        RECT 410.000 1098.010 414.000 1098.160 ;
        RECT 397.965 1097.710 414.000 1098.010 ;
        RECT 397.965 1097.695 398.295 1097.710 ;
        RECT 410.000 1097.560 414.000 1097.710 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2415.260 2519.810 2415.320 ;
        RECT 2610.110 2415.260 2610.430 2415.320 ;
        RECT 2519.490 2415.120 2610.430 2415.260 ;
        RECT 2519.490 2415.060 2519.810 2415.120 ;
        RECT 2610.110 2415.060 2610.430 2415.120 ;
        RECT 731.010 465.700 731.330 465.760 ;
        RECT 2610.110 465.700 2610.430 465.760 ;
        RECT 731.010 465.560 2610.430 465.700 ;
        RECT 731.010 465.500 731.330 465.560 ;
        RECT 2610.110 465.500 2610.430 465.560 ;
        RECT 728.250 20.300 728.570 20.360 ;
        RECT 731.010 20.300 731.330 20.360 ;
        RECT 728.250 20.160 731.330 20.300 ;
        RECT 728.250 20.100 728.570 20.160 ;
        RECT 731.010 20.100 731.330 20.160 ;
      LAYER via ;
        RECT 2519.520 2415.060 2519.780 2415.320 ;
        RECT 2610.140 2415.060 2610.400 2415.320 ;
        RECT 731.040 465.500 731.300 465.760 ;
        RECT 2610.140 465.500 2610.400 465.760 ;
        RECT 728.280 20.100 728.540 20.360 ;
        RECT 731.040 20.100 731.300 20.360 ;
      LAYER met2 ;
        RECT 2519.510 2420.955 2519.790 2421.325 ;
        RECT 2519.580 2415.350 2519.720 2420.955 ;
        RECT 2519.520 2415.030 2519.780 2415.350 ;
        RECT 2610.140 2415.030 2610.400 2415.350 ;
        RECT 2610.200 465.790 2610.340 2415.030 ;
        RECT 731.040 465.470 731.300 465.790 ;
        RECT 2610.140 465.470 2610.400 465.790 ;
        RECT 731.100 20.390 731.240 465.470 ;
        RECT 728.280 20.070 728.540 20.390 ;
        RECT 731.040 20.070 731.300 20.390 ;
        RECT 728.340 2.400 728.480 20.070 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2421.000 2519.790 2421.280 ;
      LAYER met3 ;
        RECT 2506.000 2421.290 2510.000 2421.440 ;
        RECT 2519.485 2421.290 2519.815 2421.305 ;
        RECT 2506.000 2420.990 2519.815 2421.290 ;
        RECT 2506.000 2420.840 2510.000 2420.990 ;
        RECT 2519.485 2420.975 2519.815 2420.990 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1710.810 362.680 1711.130 362.740 ;
        RECT 2449.570 362.680 2449.890 362.740 ;
        RECT 1710.810 362.540 2449.890 362.680 ;
        RECT 1710.810 362.480 1711.130 362.540 ;
        RECT 2449.570 362.480 2449.890 362.540 ;
      LAYER via ;
        RECT 1710.840 362.480 1711.100 362.740 ;
        RECT 2449.600 362.480 2449.860 362.740 ;
      LAYER met2 ;
        RECT 2450.650 510.410 2450.930 514.000 ;
        RECT 2449.660 510.270 2450.930 510.410 ;
        RECT 2449.660 362.770 2449.800 510.270 ;
        RECT 2450.650 510.000 2450.930 510.270 ;
        RECT 1710.840 362.450 1711.100 362.770 ;
        RECT 2449.600 362.450 2449.860 362.770 ;
        RECT 1710.900 17.410 1711.040 362.450 ;
        RECT 1709.520 17.270 1711.040 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2083.025 514.165 2084.115 514.335 ;
        RECT 1931.685 513.145 1931.855 513.995 ;
        RECT 1973.085 513.145 1973.255 513.995 ;
        RECT 2083.025 513.825 2083.195 514.165 ;
        RECT 2083.945 513.825 2084.115 514.165 ;
      LAYER mcon ;
        RECT 1931.685 513.825 1931.855 513.995 ;
        RECT 1973.085 513.825 1973.255 513.995 ;
      LAYER met1 ;
        RECT 1666.650 3023.860 1666.970 3023.920 ;
        RECT 2514.890 3023.860 2515.210 3023.920 ;
        RECT 1666.650 3023.720 2515.210 3023.860 ;
        RECT 1666.650 3023.660 1666.970 3023.720 ;
        RECT 2514.890 3023.660 2515.210 3023.720 ;
        RECT 2514.890 1914.780 2515.210 1914.840 ;
        RECT 2617.010 1914.780 2617.330 1914.840 ;
        RECT 2514.890 1914.640 2617.330 1914.780 ;
        RECT 2514.890 1914.580 2515.210 1914.640 ;
        RECT 2617.010 1914.580 2617.330 1914.640 ;
        RECT 1907.780 514.180 1931.840 514.320 ;
        RECT 1853.040 513.840 1870.200 513.980 ;
        RECT 1852.490 513.300 1852.810 513.360 ;
        RECT 1853.040 513.300 1853.180 513.840 ;
        RECT 1870.060 513.640 1870.200 513.840 ;
        RECT 1907.780 513.640 1907.920 514.180 ;
        RECT 1931.700 514.025 1931.840 514.180 ;
        RECT 1973.100 514.180 1980.140 514.320 ;
        RECT 1973.100 514.025 1973.240 514.180 ;
        RECT 1931.625 513.795 1931.915 514.025 ;
        RECT 1973.025 513.795 1973.315 514.025 ;
        RECT 1980.000 513.980 1980.140 514.180 ;
        RECT 2082.965 513.980 2083.255 514.025 ;
        RECT 1980.000 513.840 2083.255 513.980 ;
        RECT 2082.965 513.795 2083.255 513.840 ;
        RECT 2083.885 513.980 2084.175 514.025 ;
        RECT 2617.010 513.980 2617.330 514.040 ;
        RECT 2083.885 513.840 2617.330 513.980 ;
        RECT 2083.885 513.795 2084.175 513.840 ;
        RECT 2617.010 513.780 2617.330 513.840 ;
        RECT 1870.060 513.500 1907.920 513.640 ;
        RECT 1852.490 513.160 1853.180 513.300 ;
        RECT 1931.625 513.300 1931.915 513.345 ;
        RECT 1973.025 513.300 1973.315 513.345 ;
        RECT 1931.625 513.160 1973.315 513.300 ;
        RECT 1852.490 513.100 1852.810 513.160 ;
        RECT 1931.625 513.115 1931.915 513.160 ;
        RECT 1973.025 513.115 1973.315 513.160 ;
        RECT 1804.190 197.100 1804.510 197.160 ;
        RECT 1852.490 197.100 1852.810 197.160 ;
        RECT 1804.190 196.960 1852.810 197.100 ;
        RECT 1804.190 196.900 1804.510 196.960 ;
        RECT 1852.490 196.900 1852.810 196.960 ;
        RECT 1766.470 162.420 1766.790 162.480 ;
        RECT 1804.190 162.420 1804.510 162.480 ;
        RECT 1766.470 162.280 1804.510 162.420 ;
        RECT 1766.470 162.220 1766.790 162.280 ;
        RECT 1804.190 162.220 1804.510 162.280 ;
        RECT 1755.890 136.240 1756.210 136.300 ;
        RECT 1766.470 136.240 1766.790 136.300 ;
        RECT 1755.890 136.100 1766.790 136.240 ;
        RECT 1755.890 136.040 1756.210 136.100 ;
        RECT 1766.470 136.040 1766.790 136.100 ;
        RECT 1725.070 69.260 1725.390 69.320 ;
        RECT 1755.890 69.260 1756.210 69.320 ;
        RECT 1725.070 69.120 1756.210 69.260 ;
        RECT 1725.070 69.060 1725.390 69.120 ;
        RECT 1755.890 69.060 1756.210 69.120 ;
      LAYER via ;
        RECT 1666.680 3023.660 1666.940 3023.920 ;
        RECT 2514.920 3023.660 2515.180 3023.920 ;
        RECT 2514.920 1914.580 2515.180 1914.840 ;
        RECT 2617.040 1914.580 2617.300 1914.840 ;
        RECT 1852.520 513.100 1852.780 513.360 ;
        RECT 2617.040 513.780 2617.300 514.040 ;
        RECT 1804.220 196.900 1804.480 197.160 ;
        RECT 1852.520 196.900 1852.780 197.160 ;
        RECT 1766.500 162.220 1766.760 162.480 ;
        RECT 1804.220 162.220 1804.480 162.480 ;
        RECT 1755.920 136.040 1756.180 136.300 ;
        RECT 1766.500 136.040 1766.760 136.300 ;
        RECT 1725.100 69.060 1725.360 69.320 ;
        RECT 1755.920 69.060 1756.180 69.320 ;
      LAYER met2 ;
        RECT 1666.680 3023.630 1666.940 3023.950 ;
        RECT 2514.920 3023.630 2515.180 3023.950 ;
        RECT 1666.740 3010.000 1666.880 3023.630 ;
        RECT 1666.740 3009.340 1667.090 3010.000 ;
        RECT 1666.810 3006.000 1667.090 3009.340 ;
        RECT 2514.980 1914.870 2515.120 3023.630 ;
        RECT 2514.920 1914.550 2515.180 1914.870 ;
        RECT 2617.040 1914.550 2617.300 1914.870 ;
        RECT 2617.100 514.070 2617.240 1914.550 ;
        RECT 2617.040 513.750 2617.300 514.070 ;
        RECT 1852.520 513.070 1852.780 513.390 ;
        RECT 1852.580 197.190 1852.720 513.070 ;
        RECT 1804.220 196.870 1804.480 197.190 ;
        RECT 1852.520 196.870 1852.780 197.190 ;
        RECT 1804.280 162.510 1804.420 196.870 ;
        RECT 1766.500 162.190 1766.760 162.510 ;
        RECT 1804.220 162.190 1804.480 162.510 ;
        RECT 1766.560 136.330 1766.700 162.190 ;
        RECT 1755.920 136.010 1756.180 136.330 ;
        RECT 1766.500 136.010 1766.760 136.330 ;
        RECT 1755.980 69.350 1756.120 136.010 ;
        RECT 1725.100 69.030 1725.360 69.350 ;
        RECT 1755.920 69.030 1756.180 69.350 ;
        RECT 1725.160 17.410 1725.300 69.030 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1744.850 341.940 1745.170 342.000 ;
        RECT 2513.050 341.940 2513.370 342.000 ;
        RECT 1744.850 341.800 2513.370 341.940 ;
        RECT 1744.850 341.740 1745.170 341.800 ;
        RECT 2513.050 341.740 2513.370 341.800 ;
      LAYER via ;
        RECT 1744.880 341.740 1745.140 342.000 ;
        RECT 2513.080 341.740 2513.340 342.000 ;
      LAYER met2 ;
        RECT 2513.070 1762.715 2513.350 1763.085 ;
        RECT 2513.140 342.030 2513.280 1762.715 ;
        RECT 1744.880 341.710 1745.140 342.030 ;
        RECT 2513.080 341.710 2513.340 342.030 ;
        RECT 1744.940 7.890 1745.080 341.710 ;
        RECT 1744.940 7.750 1745.540 7.890 ;
        RECT 1745.400 2.400 1745.540 7.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 2513.070 1762.760 2513.350 1763.040 ;
      LAYER met3 ;
        RECT 2506.000 1763.050 2510.000 1763.200 ;
        RECT 2513.045 1763.050 2513.375 1763.065 ;
        RECT 2506.000 1762.750 2513.375 1763.050 ;
        RECT 2506.000 1762.600 2510.000 1762.750 ;
        RECT 2513.045 1762.735 2513.375 1762.750 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1020.810 74.700 1021.130 74.760 ;
        RECT 1759.570 74.700 1759.890 74.760 ;
        RECT 1020.810 74.560 1759.890 74.700 ;
        RECT 1020.810 74.500 1021.130 74.560 ;
        RECT 1759.570 74.500 1759.890 74.560 ;
        RECT 1759.570 62.120 1759.890 62.180 ;
        RECT 1762.790 62.120 1763.110 62.180 ;
        RECT 1759.570 61.980 1763.110 62.120 ;
        RECT 1759.570 61.920 1759.890 61.980 ;
        RECT 1762.790 61.920 1763.110 61.980 ;
      LAYER via ;
        RECT 1020.840 74.500 1021.100 74.760 ;
        RECT 1759.600 74.500 1759.860 74.760 ;
        RECT 1759.600 61.920 1759.860 62.180 ;
        RECT 1762.820 61.920 1763.080 62.180 ;
      LAYER met2 ;
        RECT 1017.290 510.410 1017.570 514.000 ;
        RECT 1017.290 510.270 1021.040 510.410 ;
        RECT 1017.290 510.000 1017.570 510.270 ;
        RECT 1020.900 74.790 1021.040 510.270 ;
        RECT 1020.840 74.470 1021.100 74.790 ;
        RECT 1759.600 74.470 1759.860 74.790 ;
        RECT 1759.660 62.210 1759.800 74.470 ;
        RECT 1759.600 61.890 1759.860 62.210 ;
        RECT 1762.820 61.890 1763.080 62.210 ;
        RECT 1762.880 2.400 1763.020 61.890 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1780.730 20.300 1781.050 20.360 ;
        RECT 1786.710 20.300 1787.030 20.360 ;
        RECT 1780.730 20.160 1787.030 20.300 ;
        RECT 1780.730 20.100 1781.050 20.160 ;
        RECT 1786.710 20.100 1787.030 20.160 ;
      LAYER via ;
        RECT 1780.760 20.100 1781.020 20.360 ;
        RECT 1786.740 20.100 1787.000 20.360 ;
      LAYER met2 ;
        RECT 2025.610 3006.690 2025.890 3010.000 ;
        RECT 2027.310 3006.690 2027.590 3006.805 ;
        RECT 2025.610 3006.550 2027.590 3006.690 ;
        RECT 2025.610 3006.000 2025.890 3006.550 ;
        RECT 2027.310 3006.435 2027.590 3006.550 ;
        RECT 2464.310 510.155 2464.590 510.525 ;
        RECT 2464.380 480.605 2464.520 510.155 ;
        RECT 1786.730 480.235 1787.010 480.605 ;
        RECT 2464.310 480.235 2464.590 480.605 ;
        RECT 1786.800 20.390 1786.940 480.235 ;
        RECT 1780.760 20.070 1781.020 20.390 ;
        RECT 1786.740 20.070 1787.000 20.390 ;
        RECT 1780.820 2.400 1780.960 20.070 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
      LAYER via2 ;
        RECT 2027.310 3006.480 2027.590 3006.760 ;
        RECT 2464.310 510.200 2464.590 510.480 ;
        RECT 1786.730 480.280 1787.010 480.560 ;
        RECT 2464.310 480.280 2464.590 480.560 ;
      LAYER met3 ;
        RECT 2027.285 3006.770 2027.615 3006.785 ;
        RECT 2045.430 3006.770 2045.810 3006.780 ;
        RECT 2027.285 3006.470 2045.810 3006.770 ;
        RECT 2027.285 3006.455 2027.615 3006.470 ;
        RECT 2045.430 3006.460 2045.810 3006.470 ;
        RECT 2045.430 3002.690 2045.810 3002.700 ;
        RECT 2471.390 3002.690 2471.770 3002.700 ;
        RECT 2045.430 3002.390 2471.770 3002.690 ;
        RECT 2045.430 3002.380 2045.810 3002.390 ;
        RECT 2471.390 3002.380 2471.770 3002.390 ;
        RECT 2468.630 512.530 2469.010 512.540 ;
        RECT 2464.990 512.230 2469.010 512.530 ;
        RECT 2464.990 511.860 2465.290 512.230 ;
        RECT 2468.630 512.220 2469.010 512.230 ;
        RECT 2464.950 511.540 2465.330 511.860 ;
        RECT 2464.285 510.490 2464.615 510.505 ;
        RECT 2464.950 510.490 2465.330 510.500 ;
        RECT 2464.285 510.190 2465.330 510.490 ;
        RECT 2464.285 510.175 2464.615 510.190 ;
        RECT 2464.950 510.180 2465.330 510.190 ;
        RECT 1786.705 480.570 1787.035 480.585 ;
        RECT 2464.285 480.570 2464.615 480.585 ;
        RECT 1786.705 480.270 2464.615 480.570 ;
        RECT 1786.705 480.255 1787.035 480.270 ;
        RECT 2464.285 480.255 2464.615 480.270 ;
      LAYER via3 ;
        RECT 2045.460 3006.460 2045.780 3006.780 ;
        RECT 2045.460 3002.380 2045.780 3002.700 ;
        RECT 2471.420 3002.380 2471.740 3002.700 ;
        RECT 2468.660 512.220 2468.980 512.540 ;
        RECT 2464.980 511.540 2465.300 511.860 ;
        RECT 2464.980 510.180 2465.300 510.500 ;
      LAYER met4 ;
        RECT 2045.455 3006.455 2045.785 3006.785 ;
        RECT 2045.470 3002.705 2045.770 3006.455 ;
        RECT 2045.455 3002.375 2045.785 3002.705 ;
        RECT 2471.415 3002.375 2471.745 3002.705 ;
        RECT 2471.430 2973.450 2471.730 3002.375 ;
        RECT 2471.430 2973.150 2472.650 2973.450 ;
        RECT 2472.350 2946.250 2472.650 2973.150 ;
        RECT 2471.430 2945.950 2472.650 2946.250 ;
        RECT 2471.430 2925.850 2471.730 2945.950 ;
        RECT 2471.430 2925.550 2472.650 2925.850 ;
        RECT 2472.350 2912.250 2472.650 2925.550 ;
        RECT 2470.510 2911.950 2472.650 2912.250 ;
        RECT 2470.510 2840.850 2470.810 2911.950 ;
        RECT 2469.590 2840.550 2470.810 2840.850 ;
        RECT 2469.590 2820.450 2469.890 2840.550 ;
        RECT 2469.590 2820.150 2470.810 2820.450 ;
        RECT 2470.510 2817.050 2470.810 2820.150 ;
        RECT 2470.510 2816.750 2472.650 2817.050 ;
        RECT 2472.350 2766.050 2472.650 2816.750 ;
        RECT 2471.430 2765.750 2472.650 2766.050 ;
        RECT 2471.430 2606.250 2471.730 2765.750 ;
        RECT 2470.510 2605.950 2471.730 2606.250 ;
        RECT 2470.510 2524.650 2470.810 2605.950 ;
        RECT 2469.590 2524.350 2470.810 2524.650 ;
        RECT 2469.590 2402.250 2469.890 2524.350 ;
        RECT 2469.590 2401.950 2470.810 2402.250 ;
        RECT 2470.510 2378.450 2470.810 2401.950 ;
        RECT 2470.510 2378.150 2472.650 2378.450 ;
        RECT 2472.350 2368.250 2472.650 2378.150 ;
        RECT 2471.430 2367.950 2472.650 2368.250 ;
        RECT 2471.430 2354.650 2471.730 2367.950 ;
        RECT 2471.430 2354.350 2473.570 2354.650 ;
        RECT 2473.270 2276.450 2473.570 2354.350 ;
        RECT 2472.350 2276.150 2473.570 2276.450 ;
        RECT 2472.350 2252.650 2472.650 2276.150 ;
        RECT 2470.510 2252.350 2472.650 2252.650 ;
        RECT 2470.510 2249.250 2470.810 2252.350 ;
        RECT 2470.510 2248.950 2473.570 2249.250 ;
        RECT 2473.270 2239.050 2473.570 2248.950 ;
        RECT 2470.510 2238.750 2473.570 2239.050 ;
        RECT 2470.510 2225.450 2470.810 2238.750 ;
        RECT 2469.590 2225.150 2470.810 2225.450 ;
        RECT 2469.590 2205.050 2469.890 2225.150 ;
        RECT 2469.590 2204.750 2473.570 2205.050 ;
        RECT 2473.270 2177.850 2473.570 2204.750 ;
        RECT 2471.430 2177.550 2473.570 2177.850 ;
        RECT 2471.430 2143.850 2471.730 2177.550 ;
        RECT 2470.510 2143.550 2471.730 2143.850 ;
        RECT 2470.510 2126.850 2470.810 2143.550 ;
        RECT 2470.510 2126.550 2473.570 2126.850 ;
        RECT 2473.270 2055.450 2473.570 2126.550 ;
        RECT 2472.350 2055.150 2473.570 2055.450 ;
        RECT 2472.350 2011.250 2472.650 2055.150 ;
        RECT 2471.430 2010.950 2472.650 2011.250 ;
        RECT 2471.430 1987.450 2471.730 2010.950 ;
        RECT 2469.590 1987.150 2471.730 1987.450 ;
        RECT 2469.590 1963.650 2469.890 1987.150 ;
        RECT 2469.590 1963.350 2471.730 1963.650 ;
        RECT 2471.430 1929.650 2471.730 1963.350 ;
        RECT 2470.510 1929.350 2471.730 1929.650 ;
        RECT 2470.510 1868.450 2470.810 1929.350 ;
        RECT 2470.510 1868.150 2471.730 1868.450 ;
        RECT 2471.430 1827.650 2471.730 1868.150 ;
        RECT 2468.670 1827.350 2471.730 1827.650 ;
        RECT 2468.670 1800.890 2468.970 1827.350 ;
        RECT 2468.230 1799.710 2469.410 1800.890 ;
        RECT 2471.910 1799.710 2473.090 1800.890 ;
        RECT 2472.350 1763.050 2472.650 1799.710 ;
        RECT 2472.350 1762.750 2473.570 1763.050 ;
        RECT 2473.270 1712.490 2473.570 1762.750 ;
        RECT 2469.150 1711.310 2470.330 1712.490 ;
        RECT 2472.830 1711.310 2474.010 1712.490 ;
        RECT 2469.590 1698.450 2469.890 1711.310 ;
        RECT 2469.590 1698.150 2473.570 1698.450 ;
        RECT 2473.270 1674.650 2473.570 1698.150 ;
        RECT 2469.590 1674.350 2473.570 1674.650 ;
        RECT 2469.590 1667.850 2469.890 1674.350 ;
        RECT 2469.590 1667.550 2470.810 1667.850 ;
        RECT 2470.510 1630.450 2470.810 1667.550 ;
        RECT 2468.670 1630.150 2470.810 1630.450 ;
        RECT 2468.670 1599.850 2468.970 1630.150 ;
        RECT 2468.670 1599.550 2473.570 1599.850 ;
        RECT 2473.270 1477.450 2473.570 1599.550 ;
        RECT 2471.430 1477.150 2473.570 1477.450 ;
        RECT 2471.430 1423.050 2471.730 1477.150 ;
        RECT 2468.670 1422.750 2471.730 1423.050 ;
        RECT 2468.670 1331.690 2468.970 1422.750 ;
        RECT 2468.230 1330.510 2469.410 1331.690 ;
        RECT 2473.750 1330.510 2474.930 1331.690 ;
        RECT 2474.190 1327.850 2474.490 1330.510 ;
        RECT 2474.190 1327.550 2476.330 1327.850 ;
        RECT 2476.030 1266.650 2476.330 1327.550 ;
        RECT 2474.190 1266.350 2476.330 1266.650 ;
        RECT 2474.190 1263.690 2474.490 1266.350 ;
        RECT 2469.150 1262.510 2470.330 1263.690 ;
        RECT 2473.750 1262.510 2474.930 1263.690 ;
        RECT 2469.590 1242.850 2469.890 1262.510 ;
        RECT 2469.590 1242.550 2473.570 1242.850 ;
        RECT 2473.270 1205.450 2473.570 1242.550 ;
        RECT 2469.590 1205.150 2473.570 1205.450 ;
        RECT 2469.590 1181.650 2469.890 1205.150 ;
        RECT 2469.590 1181.350 2470.810 1181.650 ;
        RECT 2470.510 1147.650 2470.810 1181.350 ;
        RECT 2470.510 1147.350 2471.730 1147.650 ;
        RECT 2471.430 1130.650 2471.730 1147.350 ;
        RECT 2470.510 1130.350 2471.730 1130.650 ;
        RECT 2470.510 1072.850 2470.810 1130.350 ;
        RECT 2470.510 1072.550 2473.570 1072.850 ;
        RECT 2473.270 896.050 2473.570 1072.550 ;
        RECT 2470.510 895.750 2473.570 896.050 ;
        RECT 2470.510 889.250 2470.810 895.750 ;
        RECT 2469.590 888.950 2470.810 889.250 ;
        RECT 2469.590 804.250 2469.890 888.950 ;
        RECT 2468.670 803.950 2469.890 804.250 ;
        RECT 2468.670 800.850 2468.970 803.950 ;
        RECT 2467.750 800.550 2468.970 800.850 ;
        RECT 2467.750 766.850 2468.050 800.550 ;
        RECT 2465.910 766.550 2468.050 766.850 ;
        RECT 2465.910 630.850 2466.210 766.550 ;
        RECT 2465.910 630.550 2468.050 630.850 ;
        RECT 2467.750 586.650 2468.050 630.550 ;
        RECT 2467.750 586.350 2468.970 586.650 ;
        RECT 2468.670 512.545 2468.970 586.350 ;
        RECT 2468.655 512.215 2468.985 512.545 ;
        RECT 2464.975 511.535 2465.305 511.865 ;
        RECT 2464.990 510.505 2465.290 511.535 ;
        RECT 2464.975 510.175 2465.305 510.505 ;
      LAYER met5 ;
        RECT 2468.020 1799.500 2473.300 1801.100 ;
        RECT 2468.940 1711.100 2474.220 1712.700 ;
        RECT 2468.020 1330.300 2475.140 1331.900 ;
        RECT 2468.940 1262.300 2475.140 1263.900 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 397.510 210.360 397.830 210.420 ;
        RECT 1794.070 210.360 1794.390 210.420 ;
        RECT 397.510 210.220 1794.390 210.360 ;
        RECT 397.510 210.160 397.830 210.220 ;
        RECT 1794.070 210.160 1794.390 210.220 ;
        RECT 1794.070 2.960 1794.390 3.020 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1794.070 2.820 1798.990 2.960 ;
        RECT 1794.070 2.760 1794.390 2.820 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 397.540 210.160 397.800 210.420 ;
        RECT 1794.100 210.160 1794.360 210.420 ;
        RECT 1794.100 2.760 1794.360 3.020 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 397.530 714.155 397.810 714.525 ;
        RECT 397.600 210.450 397.740 714.155 ;
        RECT 397.540 210.130 397.800 210.450 ;
        RECT 1794.100 210.130 1794.360 210.450 ;
        RECT 1794.160 3.050 1794.300 210.130 ;
        RECT 1794.100 2.730 1794.360 3.050 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 397.530 714.200 397.810 714.480 ;
      LAYER met3 ;
        RECT 397.505 714.490 397.835 714.505 ;
        RECT 410.000 714.490 414.000 714.640 ;
        RECT 397.505 714.190 414.000 714.490 ;
        RECT 397.505 714.175 397.835 714.190 ;
        RECT 410.000 714.040 414.000 714.190 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1820.750 355.540 1821.070 355.600 ;
        RECT 1856.170 355.540 1856.490 355.600 ;
        RECT 1820.750 355.400 1856.490 355.540 ;
        RECT 1820.750 355.340 1821.070 355.400 ;
        RECT 1856.170 355.340 1856.490 355.400 ;
        RECT 1816.610 16.900 1816.930 16.960 ;
        RECT 1820.750 16.900 1821.070 16.960 ;
        RECT 1816.610 16.760 1821.070 16.900 ;
        RECT 1816.610 16.700 1816.930 16.760 ;
        RECT 1820.750 16.700 1821.070 16.760 ;
      LAYER via ;
        RECT 1820.780 355.340 1821.040 355.600 ;
        RECT 1856.200 355.340 1856.460 355.600 ;
        RECT 1816.640 16.700 1816.900 16.960 ;
        RECT 1820.780 16.700 1821.040 16.960 ;
      LAYER met2 ;
        RECT 1858.170 510.410 1858.450 514.000 ;
        RECT 1856.260 510.270 1858.450 510.410 ;
        RECT 1856.260 355.630 1856.400 510.270 ;
        RECT 1858.170 510.000 1858.450 510.270 ;
        RECT 1820.780 355.310 1821.040 355.630 ;
        RECT 1856.200 355.310 1856.460 355.630 ;
        RECT 1820.840 16.990 1820.980 355.310 ;
        RECT 1816.640 16.670 1816.900 16.990 ;
        RECT 1820.780 16.670 1821.040 16.990 ;
        RECT 1816.700 2.400 1816.840 16.670 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 502.420 1153.610 502.480 ;
        RECT 1158.810 502.420 1159.130 502.480 ;
        RECT 1153.290 502.280 1159.130 502.420 ;
        RECT 1153.290 502.220 1153.610 502.280 ;
        RECT 1158.810 502.220 1159.130 502.280 ;
        RECT 1158.810 86.940 1159.130 87.000 ;
        RECT 1828.570 86.940 1828.890 87.000 ;
        RECT 1158.810 86.800 1828.890 86.940 ;
        RECT 1158.810 86.740 1159.130 86.800 ;
        RECT 1828.570 86.740 1828.890 86.800 ;
        RECT 1828.570 16.900 1828.890 16.960 ;
        RECT 1834.550 16.900 1834.870 16.960 ;
        RECT 1828.570 16.760 1834.870 16.900 ;
        RECT 1828.570 16.700 1828.890 16.760 ;
        RECT 1834.550 16.700 1834.870 16.760 ;
      LAYER via ;
        RECT 1153.320 502.220 1153.580 502.480 ;
        RECT 1158.840 502.220 1159.100 502.480 ;
        RECT 1158.840 86.740 1159.100 87.000 ;
        RECT 1828.600 86.740 1828.860 87.000 ;
        RECT 1828.600 16.700 1828.860 16.960 ;
        RECT 1834.580 16.700 1834.840 16.960 ;
      LAYER met2 ;
        RECT 1153.450 510.340 1153.730 514.000 ;
        RECT 1153.380 510.000 1153.730 510.340 ;
        RECT 1153.380 502.510 1153.520 510.000 ;
        RECT 1153.320 502.190 1153.580 502.510 ;
        RECT 1158.840 502.190 1159.100 502.510 ;
        RECT 1158.900 87.030 1159.040 502.190 ;
        RECT 1158.840 86.710 1159.100 87.030 ;
        RECT 1828.600 86.710 1828.860 87.030 ;
        RECT 1828.660 16.990 1828.800 86.710 ;
        RECT 1828.600 16.670 1828.860 16.990 ;
        RECT 1834.580 16.670 1834.840 16.990 ;
        RECT 1834.640 2.400 1834.780 16.670 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 334.800 1856.030 334.860 ;
        RECT 1891.130 334.800 1891.450 334.860 ;
        RECT 1855.710 334.660 1891.450 334.800 ;
        RECT 1855.710 334.600 1856.030 334.660 ;
        RECT 1891.130 334.600 1891.450 334.660 ;
        RECT 1852.030 16.900 1852.350 16.960 ;
        RECT 1855.710 16.900 1856.030 16.960 ;
        RECT 1852.030 16.760 1856.030 16.900 ;
        RECT 1852.030 16.700 1852.350 16.760 ;
        RECT 1855.710 16.700 1856.030 16.760 ;
      LAYER via ;
        RECT 1855.740 334.600 1856.000 334.860 ;
        RECT 1891.160 334.600 1891.420 334.860 ;
        RECT 1852.060 16.700 1852.320 16.960 ;
        RECT 1855.740 16.700 1856.000 16.960 ;
      LAYER met2 ;
        RECT 1894.970 510.410 1895.250 514.000 ;
        RECT 1891.220 510.270 1895.250 510.410 ;
        RECT 1891.220 334.890 1891.360 510.270 ;
        RECT 1894.970 510.000 1895.250 510.270 ;
        RECT 1855.740 334.570 1856.000 334.890 ;
        RECT 1891.160 334.570 1891.420 334.890 ;
        RECT 1855.800 16.990 1855.940 334.570 ;
        RECT 1852.060 16.670 1852.320 16.990 ;
        RECT 1855.740 16.670 1856.000 16.990 ;
        RECT 1852.120 2.400 1852.260 16.670 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1875.950 355.200 1876.270 355.260 ;
        RECT 2090.770 355.200 2091.090 355.260 ;
        RECT 1875.950 355.060 2091.090 355.200 ;
        RECT 1875.950 355.000 1876.270 355.060 ;
        RECT 2090.770 355.000 2091.090 355.060 ;
        RECT 1869.970 16.900 1870.290 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1869.970 16.760 1876.270 16.900 ;
        RECT 1869.970 16.700 1870.290 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1875.980 355.000 1876.240 355.260 ;
        RECT 2090.800 355.000 2091.060 355.260 ;
        RECT 1870.000 16.700 1870.260 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 2092.770 510.410 2093.050 514.000 ;
        RECT 2090.860 510.270 2093.050 510.410 ;
        RECT 2090.860 355.290 2091.000 510.270 ;
        RECT 2092.770 510.000 2093.050 510.270 ;
        RECT 1875.980 354.970 1876.240 355.290 ;
        RECT 2090.800 354.970 2091.060 355.290 ;
        RECT 1876.040 16.990 1876.180 354.970 ;
        RECT 1870.000 16.670 1870.260 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1870.060 2.400 1870.200 16.670 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 475.785 2999.905 476.875 3000.075 ;
        RECT 476.705 2999.225 476.875 2999.905 ;
        RECT 565.945 2999.225 566.115 3000.415 ;
        RECT 613.785 2999.565 613.955 3000.415 ;
        RECT 716.825 2999.735 716.995 3000.075 ;
        RECT 621.145 2999.565 621.775 2999.735 ;
        RECT 716.825 2999.565 717.455 2999.735 ;
        RECT 717.745 2999.565 717.915 3000.415 ;
        RECT 730.165 2999.565 730.335 3000.415 ;
        RECT 789.505 2999.565 790.135 2999.735 ;
        RECT 800.545 2999.225 800.715 3000.755 ;
        RECT 848.845 2999.905 849.015 3001.095 ;
        RECT 897.145 2999.905 897.315 3000.755 ;
        RECT 944.985 2999.565 945.155 3000.755 ;
        RECT 979.025 2999.565 979.655 2999.735 ;
        RECT 1014.445 2999.565 1014.615 3000.415 ;
        RECT 1062.285 2999.565 1062.455 3000.415 ;
        RECT 1075.625 2999.565 1077.175 2999.735 ;
        RECT 1111.045 2999.565 1111.215 3000.415 ;
        RECT 1158.885 2999.565 1159.055 3000.415 ;
        RECT 1172.225 2999.565 1173.775 2999.735 ;
        RECT 1207.645 2999.565 1207.815 3000.415 ;
        RECT 1255.485 2999.565 1255.655 3000.415 ;
        RECT 1268.825 2999.565 1270.375 2999.735 ;
        RECT 1304.245 2999.565 1304.415 3000.415 ;
        RECT 1352.085 2999.565 1352.255 3000.415 ;
        RECT 1352.545 2999.565 1352.715 3000.755 ;
        RECT 1400.385 2999.905 1400.555 3000.755 ;
        RECT 1418.785 2999.905 1418.955 3006.535 ;
      LAYER mcon ;
        RECT 1418.785 3006.365 1418.955 3006.535 ;
        RECT 848.845 3000.925 849.015 3001.095 ;
        RECT 800.545 3000.585 800.715 3000.755 ;
        RECT 565.945 3000.245 566.115 3000.415 ;
        RECT 613.785 3000.245 613.955 3000.415 ;
        RECT 717.745 3000.245 717.915 3000.415 ;
        RECT 716.825 2999.905 716.995 3000.075 ;
        RECT 621.605 2999.565 621.775 2999.735 ;
        RECT 717.285 2999.565 717.455 2999.735 ;
        RECT 730.165 3000.245 730.335 3000.415 ;
        RECT 789.965 2999.565 790.135 2999.735 ;
        RECT 897.145 3000.585 897.315 3000.755 ;
        RECT 944.985 3000.585 945.155 3000.755 ;
        RECT 1352.545 3000.585 1352.715 3000.755 ;
        RECT 1014.445 3000.245 1014.615 3000.415 ;
        RECT 979.485 2999.565 979.655 2999.735 ;
        RECT 1062.285 3000.245 1062.455 3000.415 ;
        RECT 1111.045 3000.245 1111.215 3000.415 ;
        RECT 1077.005 2999.565 1077.175 2999.735 ;
        RECT 1158.885 3000.245 1159.055 3000.415 ;
        RECT 1207.645 3000.245 1207.815 3000.415 ;
        RECT 1173.605 2999.565 1173.775 2999.735 ;
        RECT 1255.485 3000.245 1255.655 3000.415 ;
        RECT 1304.245 3000.245 1304.415 3000.415 ;
        RECT 1270.205 2999.565 1270.375 2999.735 ;
        RECT 1352.085 3000.245 1352.255 3000.415 ;
        RECT 1400.385 3000.585 1400.555 3000.755 ;
      LAYER met1 ;
        RECT 1418.710 3006.520 1419.030 3006.580 ;
        RECT 1418.515 3006.380 1419.030 3006.520 ;
        RECT 1418.710 3006.320 1419.030 3006.380 ;
        RECT 848.785 3001.080 849.075 3001.125 ;
        RECT 848.400 3000.940 849.075 3001.080 ;
        RECT 800.485 3000.740 800.775 3000.785 ;
        RECT 848.400 3000.740 848.540 3000.940 ;
        RECT 848.785 3000.895 849.075 3000.940 ;
        RECT 800.485 3000.600 848.540 3000.740 ;
        RECT 897.085 3000.740 897.375 3000.785 ;
        RECT 944.925 3000.740 945.215 3000.785 ;
        RECT 897.085 3000.600 945.215 3000.740 ;
        RECT 800.485 3000.555 800.775 3000.600 ;
        RECT 897.085 3000.555 897.375 3000.600 ;
        RECT 944.925 3000.555 945.215 3000.600 ;
        RECT 1352.485 3000.740 1352.775 3000.785 ;
        RECT 1400.325 3000.740 1400.615 3000.785 ;
        RECT 1352.485 3000.600 1400.615 3000.740 ;
        RECT 1352.485 3000.555 1352.775 3000.600 ;
        RECT 1400.325 3000.555 1400.615 3000.600 ;
        RECT 565.885 3000.400 566.175 3000.445 ;
        RECT 613.725 3000.400 614.015 3000.445 ;
        RECT 565.885 3000.260 614.015 3000.400 ;
        RECT 565.885 3000.215 566.175 3000.260 ;
        RECT 613.725 3000.215 614.015 3000.260 ;
        RECT 717.685 3000.400 717.975 3000.445 ;
        RECT 730.105 3000.400 730.395 3000.445 ;
        RECT 717.685 3000.260 730.395 3000.400 ;
        RECT 717.685 3000.215 717.975 3000.260 ;
        RECT 730.105 3000.215 730.395 3000.260 ;
        RECT 1014.385 3000.400 1014.675 3000.445 ;
        RECT 1062.225 3000.400 1062.515 3000.445 ;
        RECT 1014.385 3000.260 1062.515 3000.400 ;
        RECT 1014.385 3000.215 1014.675 3000.260 ;
        RECT 1062.225 3000.215 1062.515 3000.260 ;
        RECT 1110.985 3000.400 1111.275 3000.445 ;
        RECT 1158.825 3000.400 1159.115 3000.445 ;
        RECT 1110.985 3000.260 1159.115 3000.400 ;
        RECT 1110.985 3000.215 1111.275 3000.260 ;
        RECT 1158.825 3000.215 1159.115 3000.260 ;
        RECT 1207.585 3000.400 1207.875 3000.445 ;
        RECT 1255.425 3000.400 1255.715 3000.445 ;
        RECT 1207.585 3000.260 1255.715 3000.400 ;
        RECT 1207.585 3000.215 1207.875 3000.260 ;
        RECT 1255.425 3000.215 1255.715 3000.260 ;
        RECT 1304.185 3000.400 1304.475 3000.445 ;
        RECT 1352.025 3000.400 1352.315 3000.445 ;
        RECT 1304.185 3000.260 1352.315 3000.400 ;
        RECT 1304.185 3000.215 1304.475 3000.260 ;
        RECT 1352.025 3000.215 1352.315 3000.260 ;
        RECT 475.725 3000.060 476.015 3000.105 ;
        RECT 716.765 3000.060 717.055 3000.105 ;
        RECT 458.780 2999.920 476.015 3000.060 ;
        RECT 458.780 2999.380 458.920 2999.920 ;
        RECT 475.725 2999.875 476.015 2999.920 ;
        RECT 693.380 2999.920 717.055 3000.060 ;
        RECT 613.725 2999.720 614.015 2999.765 ;
        RECT 621.085 2999.720 621.375 2999.765 ;
        RECT 613.725 2999.580 621.375 2999.720 ;
        RECT 613.725 2999.535 614.015 2999.580 ;
        RECT 621.085 2999.535 621.375 2999.580 ;
        RECT 621.545 2999.720 621.835 2999.765 ;
        RECT 693.380 2999.720 693.520 2999.920 ;
        RECT 716.765 2999.875 717.055 2999.920 ;
        RECT 848.785 3000.060 849.075 3000.105 ;
        RECT 897.085 3000.060 897.375 3000.105 ;
        RECT 848.785 2999.920 897.375 3000.060 ;
        RECT 848.785 2999.875 849.075 2999.920 ;
        RECT 897.085 2999.875 897.375 2999.920 ;
        RECT 1400.325 3000.060 1400.615 3000.105 ;
        RECT 1418.725 3000.060 1419.015 3000.105 ;
        RECT 1400.325 2999.920 1419.015 3000.060 ;
        RECT 1400.325 2999.875 1400.615 2999.920 ;
        RECT 1418.725 2999.875 1419.015 2999.920 ;
        RECT 621.545 2999.580 693.520 2999.720 ;
        RECT 717.225 2999.720 717.515 2999.765 ;
        RECT 717.685 2999.720 717.975 2999.765 ;
        RECT 717.225 2999.580 717.975 2999.720 ;
        RECT 621.545 2999.535 621.835 2999.580 ;
        RECT 717.225 2999.535 717.515 2999.580 ;
        RECT 717.685 2999.535 717.975 2999.580 ;
        RECT 730.105 2999.720 730.395 2999.765 ;
        RECT 789.445 2999.720 789.735 2999.765 ;
        RECT 730.105 2999.580 789.735 2999.720 ;
        RECT 730.105 2999.535 730.395 2999.580 ;
        RECT 789.445 2999.535 789.735 2999.580 ;
        RECT 789.905 2999.535 790.195 2999.765 ;
        RECT 944.925 2999.535 945.215 2999.765 ;
        RECT 978.965 2999.720 979.255 2999.765 ;
        RECT 978.580 2999.580 979.255 2999.720 ;
        RECT 415.080 2999.240 458.920 2999.380 ;
        RECT 476.645 2999.380 476.935 2999.425 ;
        RECT 565.885 2999.380 566.175 2999.425 ;
        RECT 476.645 2999.240 566.175 2999.380 ;
        RECT 789.980 2999.380 790.120 2999.535 ;
        RECT 800.485 2999.380 800.775 2999.425 ;
        RECT 789.980 2999.240 800.775 2999.380 ;
        RECT 945.000 2999.380 945.140 2999.535 ;
        RECT 978.580 2999.380 978.720 2999.580 ;
        RECT 978.965 2999.535 979.255 2999.580 ;
        RECT 979.425 2999.535 979.715 2999.765 ;
        RECT 1014.385 2999.720 1014.675 2999.765 ;
        RECT 990.080 2999.580 1014.675 2999.720 ;
        RECT 945.000 2999.240 978.720 2999.380 ;
        RECT 979.500 2999.380 979.640 2999.535 ;
        RECT 990.080 2999.380 990.220 2999.580 ;
        RECT 1014.385 2999.535 1014.675 2999.580 ;
        RECT 1062.225 2999.535 1062.515 2999.765 ;
        RECT 1075.565 2999.535 1075.855 2999.765 ;
        RECT 1076.945 2999.720 1077.235 2999.765 ;
        RECT 1110.985 2999.720 1111.275 2999.765 ;
        RECT 1076.945 2999.580 1111.275 2999.720 ;
        RECT 1076.945 2999.535 1077.235 2999.580 ;
        RECT 1110.985 2999.535 1111.275 2999.580 ;
        RECT 1158.825 2999.535 1159.115 2999.765 ;
        RECT 1172.165 2999.535 1172.455 2999.765 ;
        RECT 1173.545 2999.720 1173.835 2999.765 ;
        RECT 1207.585 2999.720 1207.875 2999.765 ;
        RECT 1173.545 2999.580 1207.875 2999.720 ;
        RECT 1173.545 2999.535 1173.835 2999.580 ;
        RECT 1207.585 2999.535 1207.875 2999.580 ;
        RECT 1255.425 2999.535 1255.715 2999.765 ;
        RECT 1268.765 2999.535 1269.055 2999.765 ;
        RECT 1270.145 2999.720 1270.435 2999.765 ;
        RECT 1304.185 2999.720 1304.475 2999.765 ;
        RECT 1270.145 2999.580 1304.475 2999.720 ;
        RECT 1270.145 2999.535 1270.435 2999.580 ;
        RECT 1304.185 2999.535 1304.475 2999.580 ;
        RECT 1352.025 2999.535 1352.315 2999.765 ;
        RECT 1352.485 2999.535 1352.775 2999.765 ;
        RECT 979.500 2999.240 990.220 2999.380 ;
        RECT 1062.300 2999.380 1062.440 2999.535 ;
        RECT 1075.640 2999.380 1075.780 2999.535 ;
        RECT 1062.300 2999.240 1075.780 2999.380 ;
        RECT 1158.900 2999.380 1159.040 2999.535 ;
        RECT 1172.240 2999.380 1172.380 2999.535 ;
        RECT 1158.900 2999.240 1172.380 2999.380 ;
        RECT 1255.500 2999.380 1255.640 2999.535 ;
        RECT 1268.840 2999.380 1268.980 2999.535 ;
        RECT 1255.500 2999.240 1268.980 2999.380 ;
        RECT 1352.100 2999.380 1352.240 2999.535 ;
        RECT 1352.560 2999.380 1352.700 2999.535 ;
        RECT 1352.100 2999.240 1352.700 2999.380 ;
        RECT 378.190 2999.040 378.510 2999.100 ;
        RECT 415.080 2999.040 415.220 2999.240 ;
        RECT 476.645 2999.195 476.935 2999.240 ;
        RECT 565.885 2999.195 566.175 2999.240 ;
        RECT 800.485 2999.195 800.775 2999.240 ;
        RECT 378.190 2998.900 415.220 2999.040 ;
        RECT 378.190 2998.840 378.510 2998.900 ;
        RECT 378.190 495.620 378.510 495.680 ;
        RECT 745.270 495.620 745.590 495.680 ;
        RECT 378.190 495.480 745.590 495.620 ;
        RECT 378.190 495.420 378.510 495.480 ;
        RECT 745.270 495.420 745.590 495.480 ;
      LAYER via ;
        RECT 1418.740 3006.320 1419.000 3006.580 ;
        RECT 378.220 2998.840 378.480 2999.100 ;
        RECT 378.220 495.420 378.480 495.680 ;
        RECT 745.300 495.420 745.560 495.680 ;
      LAYER met2 ;
        RECT 1420.250 3006.690 1420.530 3010.000 ;
        RECT 1418.800 3006.610 1420.530 3006.690 ;
        RECT 1418.740 3006.550 1420.530 3006.610 ;
        RECT 1418.740 3006.290 1419.000 3006.550 ;
        RECT 1420.250 3006.000 1420.530 3006.550 ;
        RECT 378.220 2998.810 378.480 2999.130 ;
        RECT 378.280 495.710 378.420 2998.810 ;
        RECT 378.220 495.390 378.480 495.710 ;
        RECT 745.300 495.390 745.560 495.710 ;
        RECT 745.360 17.410 745.500 495.390 ;
        RECT 745.360 17.270 746.420 17.410 ;
        RECT 746.280 2.400 746.420 17.270 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 533.700 413.470 533.760 ;
        RECT 414.530 533.700 414.850 533.760 ;
        RECT 413.150 533.560 414.850 533.700 ;
        RECT 413.150 533.500 413.470 533.560 ;
        RECT 414.530 533.500 414.850 533.560 ;
        RECT 414.990 524.180 415.310 524.240 ;
        RECT 414.620 524.040 415.310 524.180 ;
        RECT 414.620 523.900 414.760 524.040 ;
        RECT 414.990 523.980 415.310 524.040 ;
        RECT 414.530 523.640 414.850 523.900 ;
        RECT 415.450 472.840 415.770 472.900 ;
        RECT 417.290 472.840 417.610 472.900 ;
        RECT 415.450 472.700 417.610 472.840 ;
        RECT 415.450 472.640 415.770 472.700 ;
        RECT 417.290 472.640 417.610 472.700 ;
        RECT 418.210 352.280 418.530 352.540 ;
        RECT 418.300 351.860 418.440 352.280 ;
        RECT 418.210 351.600 418.530 351.860 ;
        RECT 418.210 286.180 418.530 286.240 ;
        RECT 1883.770 286.180 1884.090 286.240 ;
        RECT 418.210 286.040 1884.090 286.180 ;
        RECT 418.210 285.980 418.530 286.040 ;
        RECT 1883.770 285.980 1884.090 286.040 ;
        RECT 1883.770 2.960 1884.090 3.020 ;
        RECT 1887.910 2.960 1888.230 3.020 ;
        RECT 1883.770 2.820 1888.230 2.960 ;
        RECT 1883.770 2.760 1884.090 2.820 ;
        RECT 1887.910 2.760 1888.230 2.820 ;
      LAYER via ;
        RECT 413.180 533.500 413.440 533.760 ;
        RECT 414.560 533.500 414.820 533.760 ;
        RECT 415.020 523.980 415.280 524.240 ;
        RECT 414.560 523.640 414.820 523.900 ;
        RECT 415.480 472.640 415.740 472.900 ;
        RECT 417.320 472.640 417.580 472.900 ;
        RECT 418.240 352.280 418.500 352.540 ;
        RECT 418.240 351.600 418.500 351.860 ;
        RECT 418.240 285.980 418.500 286.240 ;
        RECT 1883.800 285.980 1884.060 286.240 ;
        RECT 1883.800 2.760 1884.060 3.020 ;
        RECT 1887.940 2.760 1888.200 3.020 ;
      LAYER met2 ;
        RECT 413.180 533.645 413.440 533.790 ;
        RECT 413.170 533.275 413.450 533.645 ;
        RECT 414.560 533.530 414.820 533.790 ;
        RECT 414.560 533.470 415.220 533.530 ;
        RECT 414.620 533.390 415.220 533.470 ;
        RECT 415.080 524.270 415.220 533.390 ;
        RECT 415.020 523.950 415.280 524.270 ;
        RECT 414.560 523.610 414.820 523.930 ;
        RECT 414.620 498.170 414.760 523.610 ;
        RECT 414.620 498.030 415.680 498.170 ;
        RECT 415.540 472.930 415.680 498.030 ;
        RECT 415.480 472.610 415.740 472.930 ;
        RECT 417.320 472.610 417.580 472.930 ;
        RECT 417.380 425.410 417.520 472.610 ;
        RECT 417.380 425.270 418.440 425.410 ;
        RECT 418.300 352.570 418.440 425.270 ;
        RECT 418.240 352.250 418.500 352.570 ;
        RECT 418.240 351.570 418.500 351.890 ;
        RECT 418.300 286.270 418.440 351.570 ;
        RECT 418.240 285.950 418.500 286.270 ;
        RECT 1883.800 285.950 1884.060 286.270 ;
        RECT 1883.860 3.050 1884.000 285.950 ;
        RECT 1883.800 2.730 1884.060 3.050 ;
        RECT 1887.940 2.730 1888.200 3.050 ;
        RECT 1888.000 2.400 1888.140 2.730 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
      LAYER via2 ;
        RECT 413.170 533.320 413.450 533.600 ;
      LAYER met3 ;
        RECT 413.145 533.610 413.475 533.625 ;
        RECT 413.145 533.295 413.690 533.610 ;
        RECT 413.390 532.400 413.690 533.295 ;
        RECT 410.000 531.800 414.000 532.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2519.970 1799.435 2520.250 1799.805 ;
        RECT 2520.040 756.005 2520.180 1799.435 ;
        RECT 2519.970 755.635 2520.250 756.005 ;
        RECT 2509.850 634.595 2510.130 634.965 ;
        RECT 2509.920 596.885 2510.060 634.595 ;
        RECT 2509.850 596.515 2510.130 596.885 ;
        RECT 1905.870 17.155 1906.150 17.525 ;
        RECT 1905.940 2.400 1906.080 17.155 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 2519.970 1799.480 2520.250 1799.760 ;
        RECT 2519.970 755.680 2520.250 755.960 ;
        RECT 2509.850 634.640 2510.130 634.920 ;
        RECT 2509.850 596.560 2510.130 596.840 ;
        RECT 1905.870 17.200 1906.150 17.480 ;
      LAYER met3 ;
        RECT 2506.000 1799.770 2510.000 1799.920 ;
        RECT 2519.945 1799.770 2520.275 1799.785 ;
        RECT 2506.000 1799.470 2520.275 1799.770 ;
        RECT 2506.000 1799.320 2510.000 1799.470 ;
        RECT 2519.945 1799.455 2520.275 1799.470 ;
        RECT 2507.270 755.970 2507.650 755.980 ;
        RECT 2519.945 755.970 2520.275 755.985 ;
        RECT 2507.270 755.670 2520.275 755.970 ;
        RECT 2507.270 755.660 2507.650 755.670 ;
        RECT 2519.945 755.655 2520.275 755.670 ;
        RECT 2507.270 634.930 2507.650 634.940 ;
        RECT 2509.825 634.930 2510.155 634.945 ;
        RECT 2507.270 634.630 2510.155 634.930 ;
        RECT 2507.270 634.620 2507.650 634.630 ;
        RECT 2509.825 634.615 2510.155 634.630 ;
        RECT 2507.270 596.850 2507.650 596.860 ;
        RECT 2509.825 596.850 2510.155 596.865 ;
        RECT 2507.270 596.550 2510.155 596.850 ;
        RECT 2507.270 596.540 2507.650 596.550 ;
        RECT 2509.825 596.535 2510.155 596.550 ;
        RECT 1905.845 17.490 1906.175 17.505 ;
        RECT 2507.270 17.490 2507.650 17.500 ;
        RECT 1905.845 17.190 2507.650 17.490 ;
        RECT 1905.845 17.175 1906.175 17.190 ;
        RECT 2507.270 17.180 2507.650 17.190 ;
      LAYER via3 ;
        RECT 2507.300 755.660 2507.620 755.980 ;
        RECT 2507.300 634.620 2507.620 634.940 ;
        RECT 2507.300 596.540 2507.620 596.860 ;
        RECT 2507.300 17.180 2507.620 17.500 ;
      LAYER met4 ;
        RECT 2507.295 755.655 2507.625 755.985 ;
        RECT 2507.310 634.945 2507.610 755.655 ;
        RECT 2507.295 634.615 2507.625 634.945 ;
        RECT 2507.295 596.535 2507.625 596.865 ;
        RECT 2507.310 17.505 2507.610 596.535 ;
        RECT 2507.295 17.175 2507.625 17.505 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 80.480 1925.030 80.540 ;
        RECT 2297.770 80.480 2298.090 80.540 ;
        RECT 1924.710 80.340 2298.090 80.480 ;
        RECT 1924.710 80.280 1925.030 80.340 ;
        RECT 2297.770 80.280 2298.090 80.340 ;
      LAYER via ;
        RECT 1924.740 80.280 1925.000 80.540 ;
        RECT 2297.800 80.280 2298.060 80.540 ;
      LAYER met2 ;
        RECT 2302.530 510.410 2302.810 514.000 ;
        RECT 2297.860 510.270 2302.810 510.410 ;
        RECT 2297.860 80.570 2298.000 510.270 ;
        RECT 2302.530 510.000 2302.810 510.270 ;
        RECT 1924.740 80.250 1925.000 80.570 ;
        RECT 2297.800 80.250 2298.060 80.570 ;
        RECT 1924.800 17.410 1924.940 80.250 ;
        RECT 1923.420 17.270 1924.940 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2522.710 717.980 2523.030 718.040 ;
        RECT 2554.910 717.980 2555.230 718.040 ;
        RECT 2522.710 717.840 2555.230 717.980 ;
        RECT 2522.710 717.780 2523.030 717.840 ;
        RECT 2554.910 717.780 2555.230 717.840 ;
        RECT 1945.410 481.340 1945.730 481.400 ;
        RECT 2554.910 481.340 2555.230 481.400 ;
        RECT 1945.410 481.200 2555.230 481.340 ;
        RECT 1945.410 481.140 1945.730 481.200 ;
        RECT 2554.910 481.140 2555.230 481.200 ;
        RECT 1941.270 16.900 1941.590 16.960 ;
        RECT 1945.410 16.900 1945.730 16.960 ;
        RECT 1941.270 16.760 1945.730 16.900 ;
        RECT 1941.270 16.700 1941.590 16.760 ;
        RECT 1945.410 16.700 1945.730 16.760 ;
      LAYER via ;
        RECT 2522.740 717.780 2523.000 718.040 ;
        RECT 2554.940 717.780 2555.200 718.040 ;
        RECT 1945.440 481.140 1945.700 481.400 ;
        RECT 2554.940 481.140 2555.200 481.400 ;
        RECT 1941.300 16.700 1941.560 16.960 ;
        RECT 1945.440 16.700 1945.700 16.960 ;
      LAYER met2 ;
        RECT 2522.730 722.315 2523.010 722.685 ;
        RECT 2522.800 718.070 2522.940 722.315 ;
        RECT 2522.740 717.750 2523.000 718.070 ;
        RECT 2554.940 717.750 2555.200 718.070 ;
        RECT 2555.000 481.430 2555.140 717.750 ;
        RECT 1945.440 481.110 1945.700 481.430 ;
        RECT 2554.940 481.110 2555.200 481.430 ;
        RECT 1945.500 16.990 1945.640 481.110 ;
        RECT 1941.300 16.670 1941.560 16.990 ;
        RECT 1945.440 16.670 1945.700 16.990 ;
        RECT 1941.360 2.400 1941.500 16.670 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
      LAYER via2 ;
        RECT 2522.730 722.360 2523.010 722.640 ;
      LAYER met3 ;
        RECT 2506.000 722.650 2510.000 722.800 ;
        RECT 2522.705 722.650 2523.035 722.665 ;
        RECT 2506.000 722.350 2523.035 722.650 ;
        RECT 2506.000 722.200 2510.000 722.350 ;
        RECT 2522.705 722.335 2523.035 722.350 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1958.825 48.365 1958.995 96.475 ;
      LAYER mcon ;
        RECT 1958.825 96.305 1958.995 96.475 ;
      LAYER met1 ;
        RECT 1958.750 265.440 1959.070 265.500 ;
        RECT 2435.770 265.440 2436.090 265.500 ;
        RECT 1958.750 265.300 2436.090 265.440 ;
        RECT 1958.750 265.240 1959.070 265.300 ;
        RECT 2435.770 265.240 2436.090 265.300 ;
        RECT 1958.750 96.460 1959.070 96.520 ;
        RECT 1958.555 96.320 1959.070 96.460 ;
        RECT 1958.750 96.260 1959.070 96.320 ;
        RECT 1958.765 48.520 1959.055 48.565 ;
        RECT 1959.210 48.520 1959.530 48.580 ;
        RECT 1958.765 48.380 1959.530 48.520 ;
        RECT 1958.765 48.335 1959.055 48.380 ;
        RECT 1959.210 48.320 1959.530 48.380 ;
      LAYER via ;
        RECT 1958.780 265.240 1959.040 265.500 ;
        RECT 2435.800 265.240 2436.060 265.500 ;
        RECT 1958.780 96.260 1959.040 96.520 ;
        RECT 1959.240 48.320 1959.500 48.580 ;
      LAYER met2 ;
        RECT 2438.690 510.410 2438.970 514.000 ;
        RECT 2435.860 510.270 2438.970 510.410 ;
        RECT 2435.860 265.530 2436.000 510.270 ;
        RECT 2438.690 510.000 2438.970 510.270 ;
        RECT 1958.780 265.210 1959.040 265.530 ;
        RECT 2435.800 265.210 2436.060 265.530 ;
        RECT 1958.840 96.550 1958.980 265.210 ;
        RECT 1958.780 96.230 1959.040 96.550 ;
        RECT 1959.240 48.290 1959.500 48.610 ;
        RECT 1959.300 2.400 1959.440 48.290 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1099.030 3030.235 1099.310 3030.605 ;
        RECT 1099.100 3010.000 1099.240 3030.235 ;
        RECT 1099.100 3009.340 1099.450 3010.000 ;
        RECT 1099.170 3006.000 1099.450 3009.340 ;
        RECT 1977.170 45.035 1977.450 45.405 ;
        RECT 1977.240 2.400 1977.380 45.035 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
      LAYER via2 ;
        RECT 1099.030 3030.280 1099.310 3030.560 ;
        RECT 1977.170 45.080 1977.450 45.360 ;
      LAYER met3 ;
        RECT 1099.005 3030.570 1099.335 3030.585 ;
        RECT 2497.150 3030.570 2497.530 3030.580 ;
        RECT 1099.005 3030.270 2497.530 3030.570 ;
        RECT 1099.005 3030.255 1099.335 3030.270 ;
        RECT 2497.150 3030.260 2497.530 3030.270 ;
        RECT 1977.145 45.370 1977.475 45.385 ;
        RECT 2487.030 45.370 2487.410 45.380 ;
        RECT 1977.145 45.070 2487.410 45.370 ;
        RECT 1977.145 45.055 1977.475 45.070 ;
        RECT 2487.030 45.060 2487.410 45.070 ;
      LAYER via3 ;
        RECT 2497.180 3030.260 2497.500 3030.580 ;
        RECT 2487.060 45.060 2487.380 45.380 ;
      LAYER met4 ;
        RECT 2497.175 3030.255 2497.505 3030.585 ;
        RECT 2497.190 1195.250 2497.490 3030.255 ;
        RECT 2497.190 1194.950 2499.330 1195.250 ;
        RECT 2499.030 1185.050 2499.330 1194.950 ;
        RECT 2497.190 1184.750 2499.330 1185.050 ;
        RECT 2497.190 1096.650 2497.490 1184.750 ;
        RECT 2497.190 1096.350 2499.330 1096.650 ;
        RECT 2499.030 1089.850 2499.330 1096.350 ;
        RECT 2497.190 1089.550 2499.330 1089.850 ;
        RECT 2497.190 780.890 2497.490 1089.550 ;
        RECT 2486.630 779.710 2487.810 780.890 ;
        RECT 2496.750 779.710 2497.930 780.890 ;
        RECT 2487.070 45.385 2487.370 779.710 ;
        RECT 2487.055 45.055 2487.385 45.385 ;
      LAYER met5 ;
        RECT 2486.420 779.500 2498.140 781.100 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 20.300 1995.410 20.360 ;
        RECT 2000.610 20.300 2000.930 20.360 ;
        RECT 1995.090 20.160 2000.930 20.300 ;
        RECT 1995.090 20.100 1995.410 20.160 ;
        RECT 2000.610 20.100 2000.930 20.160 ;
      LAYER via ;
        RECT 1995.120 20.100 1995.380 20.360 ;
        RECT 2000.640 20.100 2000.900 20.360 ;
      LAYER met2 ;
        RECT 2431.650 3006.690 2431.930 3006.805 ;
        RECT 2433.170 3006.690 2433.450 3010.000 ;
        RECT 2431.650 3006.550 2433.450 3006.690 ;
        RECT 2431.650 3006.435 2431.930 3006.550 ;
        RECT 2433.170 3006.000 2433.450 3006.550 ;
        RECT 2000.630 251.755 2000.910 252.125 ;
        RECT 2000.700 20.390 2000.840 251.755 ;
        RECT 1995.120 20.070 1995.380 20.390 ;
        RECT 2000.640 20.070 2000.900 20.390 ;
        RECT 1995.180 2.400 1995.320 20.070 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
      LAYER via2 ;
        RECT 2431.650 3006.480 2431.930 3006.760 ;
        RECT 2000.630 251.800 2000.910 252.080 ;
      LAYER met3 ;
        RECT 2430.910 3006.770 2431.290 3006.780 ;
        RECT 2431.625 3006.770 2431.955 3006.785 ;
        RECT 2430.910 3006.470 2431.955 3006.770 ;
        RECT 2430.910 3006.460 2431.290 3006.470 ;
        RECT 2431.625 3006.455 2431.955 3006.470 ;
        RECT 2000.605 252.090 2000.935 252.105 ;
        RECT 2430.910 252.090 2431.290 252.100 ;
        RECT 2000.605 251.790 2431.290 252.090 ;
        RECT 2000.605 251.775 2000.935 251.790 ;
        RECT 2430.910 251.780 2431.290 251.790 ;
      LAYER via3 ;
        RECT 2430.940 3006.460 2431.260 3006.780 ;
        RECT 2430.940 251.780 2431.260 252.100 ;
      LAYER met4 ;
        RECT 2430.935 3006.455 2431.265 3006.785 ;
        RECT 2430.950 252.105 2431.250 3006.455 ;
        RECT 2430.935 251.775 2431.265 252.105 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1326.250 498.340 1326.570 498.400 ;
        RECT 1331.310 498.340 1331.630 498.400 ;
        RECT 1326.250 498.200 1331.630 498.340 ;
        RECT 1326.250 498.140 1326.570 498.200 ;
        RECT 1331.310 498.140 1331.630 498.200 ;
        RECT 1331.310 134.880 1331.630 134.940 ;
        RECT 2007.970 134.880 2008.290 134.940 ;
        RECT 1331.310 134.740 2008.290 134.880 ;
        RECT 1331.310 134.680 1331.630 134.740 ;
        RECT 2007.970 134.680 2008.290 134.740 ;
        RECT 2007.970 2.960 2008.290 3.020 ;
        RECT 2012.570 2.960 2012.890 3.020 ;
        RECT 2007.970 2.820 2012.890 2.960 ;
        RECT 2007.970 2.760 2008.290 2.820 ;
        RECT 2012.570 2.760 2012.890 2.820 ;
      LAYER via ;
        RECT 1326.280 498.140 1326.540 498.400 ;
        RECT 1331.340 498.140 1331.600 498.400 ;
        RECT 1331.340 134.680 1331.600 134.940 ;
        RECT 2008.000 134.680 2008.260 134.940 ;
        RECT 2008.000 2.760 2008.260 3.020 ;
        RECT 2012.600 2.760 2012.860 3.020 ;
      LAYER met2 ;
        RECT 1326.410 510.340 1326.690 514.000 ;
        RECT 1326.340 510.000 1326.690 510.340 ;
        RECT 1326.340 498.430 1326.480 510.000 ;
        RECT 1326.280 498.110 1326.540 498.430 ;
        RECT 1331.340 498.110 1331.600 498.430 ;
        RECT 1331.400 134.970 1331.540 498.110 ;
        RECT 1331.340 134.650 1331.600 134.970 ;
        RECT 2008.000 134.650 2008.260 134.970 ;
        RECT 2008.060 3.050 2008.200 134.650 ;
        RECT 2008.000 2.730 2008.260 3.050 ;
        RECT 2012.600 2.730 2012.860 3.050 ;
        RECT 2012.660 2.400 2012.800 2.730 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2030.510 33.220 2030.830 33.280 ;
        RECT 2173.570 33.220 2173.890 33.280 ;
        RECT 2030.510 33.080 2173.890 33.220 ;
        RECT 2030.510 33.020 2030.830 33.080 ;
        RECT 2173.570 33.020 2173.890 33.080 ;
      LAYER via ;
        RECT 2030.540 33.020 2030.800 33.280 ;
        RECT 2173.600 33.020 2173.860 33.280 ;
      LAYER met2 ;
        RECT 2179.250 510.410 2179.530 514.000 ;
        RECT 2173.660 510.270 2179.530 510.410 ;
        RECT 2173.660 33.310 2173.800 510.270 ;
        RECT 2179.250 510.000 2179.530 510.270 ;
        RECT 2030.540 32.990 2030.800 33.310 ;
        RECT 2173.600 32.990 2173.860 33.310 ;
        RECT 2030.600 2.400 2030.740 32.990 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 498.250 500.720 498.570 500.780 ;
        RECT 503.310 500.720 503.630 500.780 ;
        RECT 498.250 500.580 503.630 500.720 ;
        RECT 498.250 500.520 498.570 500.580 ;
        RECT 503.310 500.520 503.630 500.580 ;
        RECT 503.310 128.080 503.630 128.140 ;
        RECT 2042.470 128.080 2042.790 128.140 ;
        RECT 503.310 127.940 2042.790 128.080 ;
        RECT 503.310 127.880 503.630 127.940 ;
        RECT 2042.470 127.880 2042.790 127.940 ;
        RECT 2042.470 38.320 2042.790 38.380 ;
        RECT 2048.450 38.320 2048.770 38.380 ;
        RECT 2042.470 38.180 2048.770 38.320 ;
        RECT 2042.470 38.120 2042.790 38.180 ;
        RECT 2048.450 38.120 2048.770 38.180 ;
      LAYER via ;
        RECT 498.280 500.520 498.540 500.780 ;
        RECT 503.340 500.520 503.600 500.780 ;
        RECT 503.340 127.880 503.600 128.140 ;
        RECT 2042.500 127.880 2042.760 128.140 ;
        RECT 2042.500 38.120 2042.760 38.380 ;
        RECT 2048.480 38.120 2048.740 38.380 ;
      LAYER met2 ;
        RECT 498.410 510.340 498.690 514.000 ;
        RECT 498.340 510.000 498.690 510.340 ;
        RECT 498.340 500.810 498.480 510.000 ;
        RECT 498.280 500.490 498.540 500.810 ;
        RECT 503.340 500.490 503.600 500.810 ;
        RECT 503.400 128.170 503.540 500.490 ;
        RECT 503.340 127.850 503.600 128.170 ;
        RECT 2042.500 127.850 2042.760 128.170 ;
        RECT 2042.560 38.410 2042.700 127.850 ;
        RECT 2042.500 38.090 2042.760 38.410 ;
        RECT 2048.480 38.090 2048.740 38.410 ;
        RECT 2048.540 2.400 2048.680 38.090 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1214.720 2520.730 1214.780 ;
        RECT 2535.130 1214.720 2535.450 1214.780 ;
        RECT 2520.410 1214.580 2535.450 1214.720 ;
        RECT 2520.410 1214.520 2520.730 1214.580 ;
        RECT 2535.130 1214.520 2535.450 1214.580 ;
        RECT 765.510 245.040 765.830 245.100 ;
        RECT 2535.130 245.040 2535.450 245.100 ;
        RECT 765.510 244.900 2535.450 245.040 ;
        RECT 765.510 244.840 765.830 244.900 ;
        RECT 2535.130 244.840 2535.450 244.900 ;
      LAYER via ;
        RECT 2520.440 1214.520 2520.700 1214.780 ;
        RECT 2535.160 1214.520 2535.420 1214.780 ;
        RECT 765.540 244.840 765.800 245.100 ;
        RECT 2535.160 244.840 2535.420 245.100 ;
      LAYER met2 ;
        RECT 2520.430 1215.995 2520.710 1216.365 ;
        RECT 2520.500 1214.810 2520.640 1215.995 ;
        RECT 2520.440 1214.490 2520.700 1214.810 ;
        RECT 2535.160 1214.490 2535.420 1214.810 ;
        RECT 2535.220 245.130 2535.360 1214.490 ;
        RECT 765.540 244.810 765.800 245.130 ;
        RECT 2535.160 244.810 2535.420 245.130 ;
        RECT 765.600 17.410 765.740 244.810 ;
        RECT 763.760 17.270 765.740 17.410 ;
        RECT 763.760 2.400 763.900 17.270 ;
        RECT 763.550 -4.800 764.110 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1216.040 2520.710 1216.320 ;
      LAYER met3 ;
        RECT 2506.000 1216.330 2510.000 1216.480 ;
        RECT 2520.405 1216.330 2520.735 1216.345 ;
        RECT 2506.000 1216.030 2520.735 1216.330 ;
        RECT 2506.000 1215.880 2510.000 1216.030 ;
        RECT 2520.405 1216.015 2520.735 1216.030 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 363.470 966.180 363.790 966.240 ;
        RECT 393.370 966.180 393.690 966.240 ;
        RECT 363.470 966.040 393.690 966.180 ;
        RECT 363.470 965.980 363.790 966.040 ;
        RECT 393.370 965.980 393.690 966.040 ;
        RECT 363.470 74.020 363.790 74.080 ;
        RECT 2063.170 74.020 2063.490 74.080 ;
        RECT 363.470 73.880 2063.490 74.020 ;
        RECT 363.470 73.820 363.790 73.880 ;
        RECT 2063.170 73.820 2063.490 73.880 ;
        RECT 2063.170 62.120 2063.490 62.180 ;
        RECT 2066.390 62.120 2066.710 62.180 ;
        RECT 2063.170 61.980 2066.710 62.120 ;
        RECT 2063.170 61.920 2063.490 61.980 ;
        RECT 2066.390 61.920 2066.710 61.980 ;
      LAYER via ;
        RECT 363.500 965.980 363.760 966.240 ;
        RECT 393.400 965.980 393.660 966.240 ;
        RECT 363.500 73.820 363.760 74.080 ;
        RECT 2063.200 73.820 2063.460 74.080 ;
        RECT 2063.200 61.920 2063.460 62.180 ;
        RECT 2066.420 61.920 2066.680 62.180 ;
      LAYER met2 ;
        RECT 393.390 969.835 393.670 970.205 ;
        RECT 393.460 966.270 393.600 969.835 ;
        RECT 363.500 965.950 363.760 966.270 ;
        RECT 393.400 965.950 393.660 966.270 ;
        RECT 363.560 74.110 363.700 965.950 ;
        RECT 363.500 73.790 363.760 74.110 ;
        RECT 2063.200 73.790 2063.460 74.110 ;
        RECT 2063.260 62.210 2063.400 73.790 ;
        RECT 2063.200 61.890 2063.460 62.210 ;
        RECT 2066.420 61.890 2066.680 62.210 ;
        RECT 2066.480 2.400 2066.620 61.890 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
      LAYER via2 ;
        RECT 393.390 969.880 393.670 970.160 ;
      LAYER met3 ;
        RECT 393.365 970.170 393.695 970.185 ;
        RECT 410.000 970.170 414.000 970.320 ;
        RECT 393.365 969.870 414.000 970.170 ;
        RECT 393.365 969.855 393.695 969.870 ;
        RECT 410.000 969.720 414.000 969.870 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 32.880 1145.330 32.940 ;
        RECT 2084.330 32.880 2084.650 32.940 ;
        RECT 1145.010 32.740 2084.650 32.880 ;
        RECT 1145.010 32.680 1145.330 32.740 ;
        RECT 2084.330 32.680 2084.650 32.740 ;
      LAYER via ;
        RECT 1145.040 32.680 1145.300 32.940 ;
        RECT 2084.360 32.680 2084.620 32.940 ;
      LAYER met2 ;
        RECT 1141.490 510.410 1141.770 514.000 ;
        RECT 1141.490 510.270 1145.240 510.410 ;
        RECT 1141.490 510.000 1141.770 510.270 ;
        RECT 1145.100 32.970 1145.240 510.270 ;
        RECT 1145.040 32.650 1145.300 32.970 ;
        RECT 2084.360 32.650 2084.620 32.970 ;
        RECT 2084.420 2.400 2084.560 32.650 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.450 280.060 1772.770 280.120 ;
        RECT 2097.670 280.060 2097.990 280.120 ;
        RECT 1772.450 279.920 2097.990 280.060 ;
        RECT 1772.450 279.860 1772.770 279.920 ;
        RECT 2097.670 279.860 2097.990 279.920 ;
      LAYER via ;
        RECT 1772.480 279.860 1772.740 280.120 ;
        RECT 2097.700 279.860 2097.960 280.120 ;
      LAYER met2 ;
        RECT 1771.690 510.410 1771.970 514.000 ;
        RECT 1771.690 510.270 1772.680 510.410 ;
        RECT 1771.690 510.000 1771.970 510.270 ;
        RECT 1772.540 280.150 1772.680 510.270 ;
        RECT 1772.480 279.830 1772.740 280.150 ;
        RECT 2097.700 279.830 2097.960 280.150 ;
        RECT 2097.760 17.410 2097.900 279.830 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2099.050 3024.880 2099.370 3024.940 ;
        RECT 2567.790 3024.880 2568.110 3024.940 ;
        RECT 2099.050 3024.740 2568.110 3024.880 ;
        RECT 2099.050 3024.680 2099.370 3024.740 ;
        RECT 2567.790 3024.680 2568.110 3024.740 ;
        RECT 2119.750 32.540 2120.070 32.600 ;
        RECT 2567.790 32.540 2568.110 32.600 ;
        RECT 2119.750 32.400 2568.110 32.540 ;
        RECT 2119.750 32.340 2120.070 32.400 ;
        RECT 2567.790 32.340 2568.110 32.400 ;
      LAYER via ;
        RECT 2099.080 3024.680 2099.340 3024.940 ;
        RECT 2567.820 3024.680 2568.080 3024.940 ;
        RECT 2119.780 32.340 2120.040 32.600 ;
        RECT 2567.820 32.340 2568.080 32.600 ;
      LAYER met2 ;
        RECT 2099.080 3024.650 2099.340 3024.970 ;
        RECT 2567.820 3024.650 2568.080 3024.970 ;
        RECT 2099.140 3010.000 2099.280 3024.650 ;
        RECT 2099.140 3009.340 2099.490 3010.000 ;
        RECT 2099.210 3006.000 2099.490 3009.340 ;
        RECT 2567.880 32.630 2568.020 3024.650 ;
        RECT 2119.780 32.310 2120.040 32.630 ;
        RECT 2567.820 32.310 2568.080 32.630 ;
        RECT 2119.840 2.400 2119.980 32.310 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2132.190 334.035 2132.470 334.405 ;
        RECT 2132.260 16.730 2132.400 334.035 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
      LAYER via2 ;
        RECT 2132.190 334.080 2132.470 334.360 ;
      LAYER met3 ;
        RECT 390.350 1828.330 390.730 1828.340 ;
        RECT 410.000 1828.330 414.000 1828.480 ;
        RECT 390.350 1828.030 414.000 1828.330 ;
        RECT 390.350 1828.020 390.730 1828.030 ;
        RECT 410.000 1827.880 414.000 1828.030 ;
        RECT 390.350 334.370 390.730 334.380 ;
        RECT 2132.165 334.370 2132.495 334.385 ;
        RECT 390.350 334.070 2132.495 334.370 ;
        RECT 390.350 334.060 390.730 334.070 ;
        RECT 2132.165 334.055 2132.495 334.070 ;
      LAYER via3 ;
        RECT 390.380 1828.020 390.700 1828.340 ;
        RECT 390.380 334.060 390.700 334.380 ;
      LAYER met4 ;
        RECT 390.375 1828.015 390.705 1828.345 ;
        RECT 390.390 334.385 390.690 1828.015 ;
        RECT 390.375 334.055 390.705 334.385 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2519.490 537.780 2519.810 537.840 ;
        RECT 2521.790 537.780 2522.110 537.840 ;
        RECT 2519.490 537.640 2522.110 537.780 ;
        RECT 2519.490 537.580 2519.810 537.640 ;
        RECT 2521.790 537.580 2522.110 537.640 ;
        RECT 2197.490 507.860 2197.810 507.920 ;
        RECT 2521.790 507.860 2522.110 507.920 ;
        RECT 2197.490 507.720 2522.110 507.860 ;
        RECT 2197.490 507.660 2197.810 507.720 ;
        RECT 2521.790 507.660 2522.110 507.720 ;
        RECT 2155.630 19.280 2155.950 19.340 ;
        RECT 2197.490 19.280 2197.810 19.340 ;
        RECT 2155.630 19.140 2197.810 19.280 ;
        RECT 2155.630 19.080 2155.950 19.140 ;
        RECT 2197.490 19.080 2197.810 19.140 ;
      LAYER via ;
        RECT 2519.520 537.580 2519.780 537.840 ;
        RECT 2521.820 537.580 2522.080 537.840 ;
        RECT 2197.520 507.660 2197.780 507.920 ;
        RECT 2521.820 507.660 2522.080 507.920 ;
        RECT 2155.660 19.080 2155.920 19.340 ;
        RECT 2197.520 19.080 2197.780 19.340 ;
      LAYER met2 ;
        RECT 2519.510 1855.195 2519.790 1855.565 ;
        RECT 2519.580 537.870 2519.720 1855.195 ;
        RECT 2519.520 537.550 2519.780 537.870 ;
        RECT 2521.820 537.550 2522.080 537.870 ;
        RECT 2521.880 507.950 2522.020 537.550 ;
        RECT 2197.520 507.630 2197.780 507.950 ;
        RECT 2521.820 507.630 2522.080 507.950 ;
        RECT 2197.580 19.370 2197.720 507.630 ;
        RECT 2155.660 19.050 2155.920 19.370 ;
        RECT 2197.520 19.050 2197.780 19.370 ;
        RECT 2155.720 2.400 2155.860 19.050 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
      LAYER via2 ;
        RECT 2519.510 1855.240 2519.790 1855.520 ;
      LAYER met3 ;
        RECT 2506.000 1855.530 2510.000 1855.680 ;
        RECT 2519.485 1855.530 2519.815 1855.545 ;
        RECT 2506.000 1855.230 2519.815 1855.530 ;
        RECT 2506.000 1855.080 2510.000 1855.230 ;
        RECT 2519.485 1855.215 2519.815 1855.230 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1795.450 502.760 1795.770 502.820 ;
        RECT 1800.510 502.760 1800.830 502.820 ;
        RECT 1795.450 502.620 1800.830 502.760 ;
        RECT 1795.450 502.560 1795.770 502.620 ;
        RECT 1800.510 502.560 1800.830 502.620 ;
        RECT 1800.510 328.340 1800.830 328.400 ;
        RECT 2166.670 328.340 2166.990 328.400 ;
        RECT 1800.510 328.200 2166.990 328.340 ;
        RECT 1800.510 328.140 1800.830 328.200 ;
        RECT 2166.670 328.140 2166.990 328.200 ;
        RECT 2166.670 16.900 2166.990 16.960 ;
        RECT 2173.110 16.900 2173.430 16.960 ;
        RECT 2166.670 16.760 2173.430 16.900 ;
        RECT 2166.670 16.700 2166.990 16.760 ;
        RECT 2173.110 16.700 2173.430 16.760 ;
      LAYER via ;
        RECT 1795.480 502.560 1795.740 502.820 ;
        RECT 1800.540 502.560 1800.800 502.820 ;
        RECT 1800.540 328.140 1800.800 328.400 ;
        RECT 2166.700 328.140 2166.960 328.400 ;
        RECT 2166.700 16.700 2166.960 16.960 ;
        RECT 2173.140 16.700 2173.400 16.960 ;
      LAYER met2 ;
        RECT 1795.610 510.340 1795.890 514.000 ;
        RECT 1795.540 510.000 1795.890 510.340 ;
        RECT 1795.540 502.850 1795.680 510.000 ;
        RECT 1795.480 502.530 1795.740 502.850 ;
        RECT 1800.540 502.530 1800.800 502.850 ;
        RECT 1800.600 328.430 1800.740 502.530 ;
        RECT 1800.540 328.110 1800.800 328.430 ;
        RECT 2166.700 328.110 2166.960 328.430 ;
        RECT 2166.760 16.990 2166.900 328.110 ;
        RECT 2166.700 16.670 2166.960 16.990 ;
        RECT 2173.140 16.670 2173.400 16.990 ;
        RECT 2173.200 2.400 2173.340 16.670 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2187.850 355.115 2188.130 355.485 ;
        RECT 2187.920 16.730 2188.060 355.115 ;
        RECT 2187.920 16.590 2191.280 16.730 ;
        RECT 2191.140 2.400 2191.280 16.590 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
      LAYER via2 ;
        RECT 2187.850 355.160 2188.130 355.440 ;
      LAYER met3 ;
        RECT 397.710 2449.850 398.090 2449.860 ;
        RECT 410.000 2449.850 414.000 2450.000 ;
        RECT 397.710 2449.550 414.000 2449.850 ;
        RECT 397.710 2449.540 398.090 2449.550 ;
        RECT 410.000 2449.400 414.000 2449.550 ;
        RECT 397.710 355.450 398.090 355.460 ;
        RECT 2187.825 355.450 2188.155 355.465 ;
        RECT 397.710 355.150 2188.155 355.450 ;
        RECT 397.710 355.140 398.090 355.150 ;
        RECT 2187.825 355.135 2188.155 355.150 ;
      LAYER via3 ;
        RECT 397.740 2449.540 398.060 2449.860 ;
        RECT 397.740 355.140 398.060 355.460 ;
      LAYER met4 ;
        RECT 397.735 2449.535 398.065 2449.865 ;
        RECT 397.750 355.465 398.050 2449.535 ;
        RECT 397.735 355.135 398.065 355.465 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1959.210 203.900 1959.530 203.960 ;
        RECT 2208.070 203.900 2208.390 203.960 ;
        RECT 1959.210 203.760 2208.390 203.900 ;
        RECT 1959.210 203.700 1959.530 203.760 ;
        RECT 2208.070 203.700 2208.390 203.760 ;
      LAYER via ;
        RECT 1959.240 203.700 1959.500 203.960 ;
        RECT 2208.100 203.700 2208.360 203.960 ;
      LAYER met2 ;
        RECT 1956.610 510.410 1956.890 514.000 ;
        RECT 1956.610 510.270 1959.440 510.410 ;
        RECT 1956.610 510.000 1956.890 510.270 ;
        RECT 1959.300 203.990 1959.440 510.270 ;
        RECT 1959.240 203.670 1959.500 203.990 ;
        RECT 2208.100 203.670 2208.360 203.990 ;
        RECT 2208.160 16.730 2208.300 203.670 ;
        RECT 2208.160 16.590 2209.220 16.730 ;
        RECT 2209.080 2.400 2209.220 16.590 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 397.050 458.900 397.370 458.960 ;
        RECT 2221.870 458.900 2222.190 458.960 ;
        RECT 397.050 458.760 2222.190 458.900 ;
        RECT 397.050 458.700 397.370 458.760 ;
        RECT 2221.870 458.700 2222.190 458.760 ;
      LAYER via ;
        RECT 397.080 458.700 397.340 458.960 ;
        RECT 2221.900 458.700 2222.160 458.960 ;
      LAYER met2 ;
        RECT 397.070 623.035 397.350 623.405 ;
        RECT 397.140 458.990 397.280 623.035 ;
        RECT 397.080 458.670 397.340 458.990 ;
        RECT 2221.900 458.670 2222.160 458.990 ;
        RECT 2221.960 16.730 2222.100 458.670 ;
        RECT 2221.960 16.590 2227.160 16.730 ;
        RECT 2227.020 2.400 2227.160 16.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
      LAYER via2 ;
        RECT 397.070 623.080 397.350 623.360 ;
      LAYER met3 ;
        RECT 397.045 623.370 397.375 623.385 ;
        RECT 410.000 623.370 414.000 623.520 ;
        RECT 397.045 623.070 414.000 623.370 ;
        RECT 397.045 623.055 397.375 623.070 ;
        RECT 410.000 622.920 414.000 623.070 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 385.090 2794.700 385.410 2794.760 ;
        RECT 397.970 2794.700 398.290 2794.760 ;
        RECT 385.090 2794.560 398.290 2794.700 ;
        RECT 385.090 2794.500 385.410 2794.560 ;
        RECT 397.970 2794.500 398.290 2794.560 ;
        RECT 385.090 424.560 385.410 424.620 ;
        RECT 779.770 424.560 780.090 424.620 ;
        RECT 385.090 424.420 780.090 424.560 ;
        RECT 385.090 424.360 385.410 424.420 ;
        RECT 779.770 424.360 780.090 424.420 ;
      LAYER via ;
        RECT 385.120 2794.500 385.380 2794.760 ;
        RECT 398.000 2794.500 398.260 2794.760 ;
        RECT 385.120 424.360 385.380 424.620 ;
        RECT 779.800 424.360 780.060 424.620 ;
      LAYER met2 ;
        RECT 397.990 2796.315 398.270 2796.685 ;
        RECT 398.060 2794.790 398.200 2796.315 ;
        RECT 385.120 2794.470 385.380 2794.790 ;
        RECT 398.000 2794.470 398.260 2794.790 ;
        RECT 385.180 424.650 385.320 2794.470 ;
        RECT 385.120 424.330 385.380 424.650 ;
        RECT 779.800 424.330 780.060 424.650 ;
        RECT 779.860 17.410 780.000 424.330 ;
        RECT 779.860 17.270 781.840 17.410 ;
        RECT 781.700 2.400 781.840 17.270 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 397.990 2796.360 398.270 2796.640 ;
      LAYER met3 ;
        RECT 397.965 2796.650 398.295 2796.665 ;
        RECT 410.000 2796.650 414.000 2796.800 ;
        RECT 397.965 2796.350 414.000 2796.650 ;
        RECT 397.965 2796.335 398.295 2796.350 ;
        RECT 410.000 2796.200 414.000 2796.350 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2242.570 62.120 2242.890 62.180 ;
        RECT 2244.870 62.120 2245.190 62.180 ;
        RECT 2242.570 61.980 2245.190 62.120 ;
        RECT 2242.570 61.920 2242.890 61.980 ;
        RECT 2244.870 61.920 2245.190 61.980 ;
      LAYER via ;
        RECT 2242.600 61.920 2242.860 62.180 ;
        RECT 2244.900 61.920 2245.160 62.180 ;
      LAYER met2 ;
        RECT 2242.590 430.595 2242.870 430.965 ;
        RECT 2242.660 62.210 2242.800 430.595 ;
        RECT 2242.600 61.890 2242.860 62.210 ;
        RECT 2244.900 61.890 2245.160 62.210 ;
        RECT 2244.960 2.400 2245.100 61.890 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
      LAYER via2 ;
        RECT 2242.590 430.640 2242.870 430.920 ;
      LAYER met3 ;
        RECT 406.910 2906.810 407.290 2906.820 ;
        RECT 410.000 2906.810 414.000 2906.960 ;
        RECT 406.910 2906.510 414.000 2906.810 ;
        RECT 406.910 2906.500 407.290 2906.510 ;
        RECT 410.000 2906.360 414.000 2906.510 ;
        RECT 406.910 430.930 407.290 430.940 ;
        RECT 2242.565 430.930 2242.895 430.945 ;
        RECT 406.910 430.630 2242.895 430.930 ;
        RECT 406.910 430.620 407.290 430.630 ;
        RECT 2242.565 430.615 2242.895 430.630 ;
      LAYER via3 ;
        RECT 406.940 2906.500 407.260 2906.820 ;
        RECT 406.940 430.620 407.260 430.940 ;
      LAYER met4 ;
        RECT 406.935 2906.495 407.265 2906.825 ;
        RECT 406.950 430.945 407.250 2906.495 ;
        RECT 406.935 430.615 407.265 430.945 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 396.130 417.420 396.450 417.480 ;
        RECT 2256.370 417.420 2256.690 417.480 ;
        RECT 396.130 417.280 2256.690 417.420 ;
        RECT 396.130 417.220 396.450 417.280 ;
        RECT 2256.370 417.220 2256.690 417.280 ;
        RECT 2256.370 37.980 2256.690 38.040 ;
        RECT 2262.350 37.980 2262.670 38.040 ;
        RECT 2256.370 37.840 2262.670 37.980 ;
        RECT 2256.370 37.780 2256.690 37.840 ;
        RECT 2262.350 37.780 2262.670 37.840 ;
      LAYER via ;
        RECT 396.160 417.220 396.420 417.480 ;
        RECT 2256.400 417.220 2256.660 417.480 ;
        RECT 2256.400 37.780 2256.660 38.040 ;
        RECT 2262.380 37.780 2262.640 38.040 ;
      LAYER met2 ;
        RECT 396.150 933.115 396.430 933.485 ;
        RECT 396.220 417.510 396.360 933.115 ;
        RECT 396.160 417.190 396.420 417.510 ;
        RECT 2256.400 417.190 2256.660 417.510 ;
        RECT 2256.460 38.070 2256.600 417.190 ;
        RECT 2256.400 37.750 2256.660 38.070 ;
        RECT 2262.380 37.750 2262.640 38.070 ;
        RECT 2262.440 2.400 2262.580 37.750 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
      LAYER via2 ;
        RECT 396.150 933.160 396.430 933.440 ;
      LAYER met3 ;
        RECT 396.125 933.450 396.455 933.465 ;
        RECT 410.000 933.450 414.000 933.600 ;
        RECT 396.125 933.150 414.000 933.450 ;
        RECT 396.125 933.135 396.455 933.150 ;
        RECT 410.000 933.000 414.000 933.150 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2562.805 481.525 2562.975 482.715 ;
      LAYER mcon ;
        RECT 2562.805 482.545 2562.975 482.715 ;
      LAYER met1 ;
        RECT 2520.410 1690.720 2520.730 1690.780 ;
        RECT 2596.310 1690.720 2596.630 1690.780 ;
        RECT 2520.410 1690.580 2596.630 1690.720 ;
        RECT 2520.410 1690.520 2520.730 1690.580 ;
        RECT 2596.310 1690.520 2596.630 1690.580 ;
        RECT 2283.050 482.700 2283.370 482.760 ;
        RECT 2562.745 482.700 2563.035 482.745 ;
        RECT 2283.050 482.560 2563.035 482.700 ;
        RECT 2283.050 482.500 2283.370 482.560 ;
        RECT 2562.745 482.515 2563.035 482.560 ;
        RECT 2562.745 481.680 2563.035 481.725 ;
        RECT 2596.310 481.680 2596.630 481.740 ;
        RECT 2562.745 481.540 2596.630 481.680 ;
        RECT 2562.745 481.495 2563.035 481.540 ;
        RECT 2596.310 481.480 2596.630 481.540 ;
        RECT 2280.290 20.300 2280.610 20.360 ;
        RECT 2283.050 20.300 2283.370 20.360 ;
        RECT 2280.290 20.160 2283.370 20.300 ;
        RECT 2280.290 20.100 2280.610 20.160 ;
        RECT 2283.050 20.100 2283.370 20.160 ;
      LAYER via ;
        RECT 2520.440 1690.520 2520.700 1690.780 ;
        RECT 2596.340 1690.520 2596.600 1690.780 ;
        RECT 2283.080 482.500 2283.340 482.760 ;
        RECT 2596.340 481.480 2596.600 481.740 ;
        RECT 2280.320 20.100 2280.580 20.360 ;
        RECT 2283.080 20.100 2283.340 20.360 ;
      LAYER met2 ;
        RECT 2520.430 1690.635 2520.710 1691.005 ;
        RECT 2520.440 1690.490 2520.700 1690.635 ;
        RECT 2596.340 1690.490 2596.600 1690.810 ;
        RECT 2283.080 482.470 2283.340 482.790 ;
        RECT 2283.140 20.390 2283.280 482.470 ;
        RECT 2596.400 481.770 2596.540 1690.490 ;
        RECT 2596.340 481.450 2596.600 481.770 ;
        RECT 2280.320 20.070 2280.580 20.390 ;
        RECT 2283.080 20.070 2283.340 20.390 ;
        RECT 2280.380 2.400 2280.520 20.070 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1690.680 2520.710 1690.960 ;
      LAYER met3 ;
        RECT 2506.000 1690.970 2510.000 1691.120 ;
        RECT 2520.405 1690.970 2520.735 1690.985 ;
        RECT 2506.000 1690.670 2520.735 1690.970 ;
        RECT 2506.000 1690.520 2510.000 1690.670 ;
        RECT 2520.405 1690.655 2520.735 1690.670 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1149.610 3009.240 1149.930 3009.300 ;
        RECT 2553.070 3009.240 2553.390 3009.300 ;
        RECT 1149.610 3009.100 2553.390 3009.240 ;
        RECT 1149.610 3009.040 1149.930 3009.100 ;
        RECT 2553.070 3009.040 2553.390 3009.100 ;
        RECT 2298.230 33.220 2298.550 33.280 ;
        RECT 2553.070 33.220 2553.390 33.280 ;
        RECT 2298.230 33.080 2553.390 33.220 ;
        RECT 2298.230 33.020 2298.550 33.080 ;
        RECT 2553.070 33.020 2553.390 33.080 ;
      LAYER via ;
        RECT 1149.640 3009.040 1149.900 3009.300 ;
        RECT 2553.100 3009.040 2553.360 3009.300 ;
        RECT 2298.260 33.020 2298.520 33.280 ;
        RECT 2553.100 33.020 2553.360 33.280 ;
      LAYER met2 ;
        RECT 1147.930 3009.410 1148.210 3010.000 ;
        RECT 1147.930 3009.330 1149.840 3009.410 ;
        RECT 1147.930 3009.270 1149.900 3009.330 ;
        RECT 1147.930 3006.000 1148.210 3009.270 ;
        RECT 1149.640 3009.010 1149.900 3009.270 ;
        RECT 2553.100 3009.010 2553.360 3009.330 ;
        RECT 2553.160 33.310 2553.300 3009.010 ;
        RECT 2298.260 32.990 2298.520 33.310 ;
        RECT 2553.100 32.990 2553.360 33.310 ;
        RECT 2298.320 2.400 2298.460 32.990 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 487.460 2318.330 487.520 ;
        RECT 2526.850 487.460 2527.170 487.520 ;
        RECT 2318.010 487.320 2527.170 487.460 ;
        RECT 2318.010 487.260 2318.330 487.320 ;
        RECT 2526.850 487.260 2527.170 487.320 ;
      LAYER via ;
        RECT 2318.040 487.260 2318.300 487.520 ;
        RECT 2526.880 487.260 2527.140 487.520 ;
      LAYER met2 ;
        RECT 2526.870 1653.915 2527.150 1654.285 ;
        RECT 2526.940 487.550 2527.080 1653.915 ;
        RECT 2318.040 487.230 2318.300 487.550 ;
        RECT 2526.880 487.230 2527.140 487.550 ;
        RECT 2318.100 17.410 2318.240 487.230 ;
        RECT 2316.260 17.270 2318.240 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 2526.870 1653.960 2527.150 1654.240 ;
      LAYER met3 ;
        RECT 2506.000 1654.250 2510.000 1654.400 ;
        RECT 2526.845 1654.250 2527.175 1654.265 ;
        RECT 2506.000 1653.950 2527.175 1654.250 ;
        RECT 2506.000 1653.800 2510.000 1653.950 ;
        RECT 2526.845 1653.935 2527.175 1653.950 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2338.710 300.460 2339.030 300.520 ;
        RECT 2470.270 300.460 2470.590 300.520 ;
        RECT 2338.710 300.320 2470.590 300.460 ;
        RECT 2338.710 300.260 2339.030 300.320 ;
        RECT 2470.270 300.260 2470.590 300.320 ;
        RECT 2334.110 20.300 2334.430 20.360 ;
        RECT 2338.710 20.300 2339.030 20.360 ;
        RECT 2334.110 20.160 2339.030 20.300 ;
        RECT 2334.110 20.100 2334.430 20.160 ;
        RECT 2338.710 20.100 2339.030 20.160 ;
      LAYER via ;
        RECT 2338.740 300.260 2339.000 300.520 ;
        RECT 2470.300 300.260 2470.560 300.520 ;
        RECT 2334.140 20.100 2334.400 20.360 ;
        RECT 2338.740 20.100 2339.000 20.360 ;
      LAYER met2 ;
        RECT 2475.490 510.410 2475.770 514.000 ;
        RECT 2470.360 510.270 2475.770 510.410 ;
        RECT 2470.360 300.550 2470.500 510.270 ;
        RECT 2475.490 510.000 2475.770 510.270 ;
        RECT 2338.740 300.230 2339.000 300.550 ;
        RECT 2470.300 300.230 2470.560 300.550 ;
        RECT 2338.800 20.390 2338.940 300.230 ;
        RECT 2334.140 20.070 2334.400 20.390 ;
        RECT 2338.740 20.070 2339.000 20.390 ;
        RECT 2334.200 2.400 2334.340 20.070 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 703.410 3022.500 703.730 3022.560 ;
        RECT 2518.570 3022.500 2518.890 3022.560 ;
        RECT 703.410 3022.360 2518.890 3022.500 ;
        RECT 703.410 3022.300 703.730 3022.360 ;
        RECT 2518.570 3022.300 2518.890 3022.360 ;
        RECT 2351.590 19.960 2351.910 20.020 ;
        RECT 2470.730 19.960 2471.050 20.020 ;
        RECT 2351.590 19.820 2471.050 19.960 ;
        RECT 2351.590 19.760 2351.910 19.820 ;
        RECT 2470.730 19.760 2471.050 19.820 ;
      LAYER via ;
        RECT 703.440 3022.300 703.700 3022.560 ;
        RECT 2518.600 3022.300 2518.860 3022.560 ;
        RECT 2351.620 19.760 2351.880 20.020 ;
        RECT 2470.760 19.760 2471.020 20.020 ;
      LAYER met2 ;
        RECT 703.440 3022.270 703.700 3022.590 ;
        RECT 2518.600 3022.270 2518.860 3022.590 ;
        RECT 703.500 3010.000 703.640 3022.270 ;
        RECT 703.500 3009.340 703.850 3010.000 ;
        RECT 703.570 3006.000 703.850 3009.340 ;
        RECT 2518.660 870.245 2518.800 3022.270 ;
        RECT 2518.590 869.875 2518.870 870.245 ;
        RECT 2470.750 509.475 2471.030 509.845 ;
        RECT 2470.820 20.050 2470.960 509.475 ;
        RECT 2351.620 19.730 2351.880 20.050 ;
        RECT 2470.760 19.730 2471.020 20.050 ;
        RECT 2351.680 2.400 2351.820 19.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
      LAYER via2 ;
        RECT 2518.590 869.920 2518.870 870.200 ;
        RECT 2470.750 509.520 2471.030 509.800 ;
      LAYER met3 ;
        RECT 2518.565 870.220 2518.895 870.225 ;
        RECT 2518.310 870.210 2518.895 870.220 ;
        RECT 2518.110 869.910 2518.895 870.210 ;
        RECT 2518.310 869.900 2518.895 869.910 ;
        RECT 2518.565 869.895 2518.895 869.900 ;
        RECT 2475.990 511.170 2476.370 511.180 ;
        RECT 2470.510 510.870 2476.370 511.170 ;
        RECT 2470.510 509.825 2470.810 510.870 ;
        RECT 2475.990 510.860 2476.370 510.870 ;
        RECT 2470.510 509.510 2471.055 509.825 ;
        RECT 2470.725 509.495 2471.055 509.510 ;
      LAYER via3 ;
        RECT 2518.340 869.900 2518.660 870.220 ;
        RECT 2476.020 510.860 2476.340 511.180 ;
      LAYER met4 ;
        RECT 2518.335 869.895 2518.665 870.225 ;
        RECT 2518.350 868.850 2518.650 869.895 ;
        RECT 2517.430 868.550 2518.650 868.850 ;
        RECT 2517.430 865.890 2517.730 868.550 ;
        RECT 2475.590 864.710 2476.770 865.890 ;
        RECT 2516.990 864.710 2518.170 865.890 ;
        RECT 2476.030 824.650 2476.330 864.710 ;
        RECT 2473.270 824.350 2476.330 824.650 ;
        RECT 2473.270 651.250 2473.570 824.350 ;
        RECT 2473.270 650.950 2474.490 651.250 ;
        RECT 2474.190 634.930 2474.490 650.950 ;
        RECT 2473.270 634.630 2474.490 634.930 ;
        RECT 2473.270 634.250 2473.570 634.630 ;
        RECT 2473.270 633.950 2474.490 634.250 ;
        RECT 2474.190 617.690 2474.490 633.950 ;
        RECT 2465.470 616.510 2466.650 617.690 ;
        RECT 2473.750 616.510 2474.930 617.690 ;
        RECT 2465.910 600.690 2466.210 616.510 ;
        RECT 2465.470 599.510 2466.650 600.690 ;
        RECT 2475.590 599.510 2476.770 600.690 ;
        RECT 2476.030 545.850 2476.330 599.510 ;
        RECT 2476.030 545.550 2476.560 545.850 ;
        RECT 2476.260 542.450 2476.560 545.550 ;
        RECT 2476.030 542.150 2476.560 542.450 ;
        RECT 2476.030 511.185 2476.330 542.150 ;
        RECT 2476.015 510.855 2476.345 511.185 ;
      LAYER met5 ;
        RECT 2475.380 864.500 2518.380 866.100 ;
        RECT 2465.260 616.300 2475.140 617.900 ;
        RECT 2465.260 599.300 2476.980 600.900 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 475.710 107.000 476.030 107.060 ;
        RECT 2366.770 107.000 2367.090 107.060 ;
        RECT 475.710 106.860 2367.090 107.000 ;
        RECT 475.710 106.800 476.030 106.860 ;
        RECT 2366.770 106.800 2367.090 106.860 ;
        RECT 2366.770 62.120 2367.090 62.180 ;
        RECT 2369.530 62.120 2369.850 62.180 ;
        RECT 2366.770 61.980 2369.850 62.120 ;
        RECT 2366.770 61.920 2367.090 61.980 ;
        RECT 2369.530 61.920 2369.850 61.980 ;
      LAYER via ;
        RECT 475.740 106.800 476.000 107.060 ;
        RECT 2366.800 106.800 2367.060 107.060 ;
        RECT 2366.800 61.920 2367.060 62.180 ;
        RECT 2369.560 61.920 2369.820 62.180 ;
      LAYER met2 ;
        RECT 474.490 510.410 474.770 514.000 ;
        RECT 474.490 510.270 475.940 510.410 ;
        RECT 474.490 510.000 474.770 510.270 ;
        RECT 475.800 107.090 475.940 510.270 ;
        RECT 475.740 106.770 476.000 107.090 ;
        RECT 2366.800 106.770 2367.060 107.090 ;
        RECT 2366.860 62.210 2367.000 106.770 ;
        RECT 2366.800 61.890 2367.060 62.210 ;
        RECT 2369.560 61.890 2369.820 62.210 ;
        RECT 2369.620 2.400 2369.760 61.890 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2482.305 16.745 2482.475 19.635 ;
      LAYER mcon ;
        RECT 2482.305 19.465 2482.475 19.635 ;
      LAYER met1 ;
        RECT 2371.370 3011.280 2371.690 3011.340 ;
        RECT 2539.270 3011.280 2539.590 3011.340 ;
        RECT 2371.370 3011.140 2539.590 3011.280 ;
        RECT 2371.370 3011.080 2371.690 3011.140 ;
        RECT 2539.270 3011.080 2539.590 3011.140 ;
        RECT 2387.470 19.620 2387.790 19.680 ;
        RECT 2482.245 19.620 2482.535 19.665 ;
        RECT 2387.470 19.480 2482.535 19.620 ;
        RECT 2387.470 19.420 2387.790 19.480 ;
        RECT 2482.245 19.435 2482.535 19.480 ;
        RECT 2482.245 16.900 2482.535 16.945 ;
        RECT 2539.270 16.900 2539.590 16.960 ;
        RECT 2482.245 16.760 2539.590 16.900 ;
        RECT 2482.245 16.715 2482.535 16.760 ;
        RECT 2539.270 16.700 2539.590 16.760 ;
      LAYER via ;
        RECT 2371.400 3011.080 2371.660 3011.340 ;
        RECT 2539.300 3011.080 2539.560 3011.340 ;
        RECT 2387.500 19.420 2387.760 19.680 ;
        RECT 2539.300 16.700 2539.560 16.960 ;
      LAYER met2 ;
        RECT 2371.400 3011.050 2371.660 3011.370 ;
        RECT 2539.300 3011.050 2539.560 3011.370 ;
        RECT 2371.460 3010.000 2371.600 3011.050 ;
        RECT 2371.460 3009.340 2371.810 3010.000 ;
        RECT 2371.530 3006.000 2371.810 3009.340 ;
        RECT 2387.500 19.390 2387.760 19.710 ;
        RECT 2387.560 2.400 2387.700 19.390 ;
        RECT 2539.360 16.990 2539.500 3011.050 ;
        RECT 2539.300 16.670 2539.560 16.990 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2521.865 2980.865 2522.035 3008.915 ;
        RECT 2521.865 2656.505 2522.035 2670.955 ;
        RECT 2522.325 2621.485 2522.495 2656.335 ;
        RECT 2521.865 2559.945 2522.035 2574.055 ;
        RECT 2521.865 2173.705 2522.035 2221.815 ;
        RECT 2521.865 2077.145 2522.035 2125.255 ;
      LAYER mcon ;
        RECT 2521.865 3008.745 2522.035 3008.915 ;
        RECT 2521.865 2670.785 2522.035 2670.955 ;
        RECT 2522.325 2656.165 2522.495 2656.335 ;
        RECT 2521.865 2573.885 2522.035 2574.055 ;
        RECT 2521.865 2221.645 2522.035 2221.815 ;
        RECT 2521.865 2125.085 2522.035 2125.255 ;
      LAYER met1 ;
        RECT 2297.770 3008.900 2298.090 3008.960 ;
        RECT 2521.805 3008.900 2522.095 3008.945 ;
        RECT 2297.770 3008.760 2522.095 3008.900 ;
        RECT 2297.770 3008.700 2298.090 3008.760 ;
        RECT 2521.805 3008.715 2522.095 3008.760 ;
        RECT 2521.790 2981.020 2522.110 2981.080 ;
        RECT 2521.595 2980.880 2522.110 2981.020 ;
        RECT 2521.790 2980.820 2522.110 2980.880 ;
        RECT 2521.790 2891.260 2522.110 2891.320 ;
        RECT 2522.250 2891.260 2522.570 2891.320 ;
        RECT 2521.790 2891.120 2522.570 2891.260 ;
        RECT 2521.790 2891.060 2522.110 2891.120 ;
        RECT 2522.250 2891.060 2522.570 2891.120 ;
        RECT 2521.790 2864.060 2522.110 2864.120 ;
        RECT 2521.420 2863.920 2522.110 2864.060 ;
        RECT 2521.420 2863.440 2521.560 2863.920 ;
        RECT 2521.790 2863.860 2522.110 2863.920 ;
        RECT 2521.330 2863.180 2521.650 2863.440 ;
        RECT 2521.790 2814.760 2522.110 2814.820 ;
        RECT 2522.710 2814.760 2523.030 2814.820 ;
        RECT 2521.790 2814.620 2523.030 2814.760 ;
        RECT 2521.790 2814.560 2522.110 2814.620 ;
        RECT 2522.710 2814.560 2523.030 2814.620 ;
        RECT 2521.805 2670.940 2522.095 2670.985 ;
        RECT 2522.250 2670.940 2522.570 2671.000 ;
        RECT 2521.805 2670.800 2522.570 2670.940 ;
        RECT 2521.805 2670.755 2522.095 2670.800 ;
        RECT 2522.250 2670.740 2522.570 2670.800 ;
        RECT 2521.790 2656.660 2522.110 2656.720 ;
        RECT 2521.595 2656.520 2522.110 2656.660 ;
        RECT 2521.790 2656.460 2522.110 2656.520 ;
        RECT 2522.250 2656.320 2522.570 2656.380 ;
        RECT 2522.055 2656.180 2522.570 2656.320 ;
        RECT 2522.250 2656.120 2522.570 2656.180 ;
        RECT 2522.250 2621.640 2522.570 2621.700 ;
        RECT 2522.055 2621.500 2522.570 2621.640 ;
        RECT 2522.250 2621.440 2522.570 2621.500 ;
        RECT 2521.790 2574.040 2522.110 2574.100 ;
        RECT 2521.595 2573.900 2522.110 2574.040 ;
        RECT 2521.790 2573.840 2522.110 2573.900 ;
        RECT 2521.790 2560.100 2522.110 2560.160 ;
        RECT 2521.595 2559.960 2522.110 2560.100 ;
        RECT 2521.790 2559.900 2522.110 2559.960 ;
        RECT 2521.790 2525.560 2522.110 2525.820 ;
        RECT 2521.880 2525.080 2522.020 2525.560 ;
        RECT 2522.250 2525.080 2522.570 2525.140 ;
        RECT 2521.880 2524.940 2522.570 2525.080 ;
        RECT 2522.250 2524.880 2522.570 2524.940 ;
        RECT 2520.870 2487.680 2521.190 2487.740 ;
        RECT 2521.790 2487.680 2522.110 2487.740 ;
        RECT 2520.870 2487.540 2522.110 2487.680 ;
        RECT 2520.870 2487.480 2521.190 2487.540 ;
        RECT 2521.790 2487.480 2522.110 2487.540 ;
        RECT 2521.790 2429.000 2522.110 2429.260 ;
        RECT 2521.880 2428.520 2522.020 2429.000 ;
        RECT 2522.250 2428.520 2522.570 2428.580 ;
        RECT 2521.880 2428.380 2522.570 2428.520 ;
        RECT 2522.250 2428.320 2522.570 2428.380 ;
        RECT 2522.250 2414.920 2522.570 2414.980 ;
        RECT 2523.170 2414.920 2523.490 2414.980 ;
        RECT 2522.250 2414.780 2523.490 2414.920 ;
        RECT 2522.250 2414.720 2522.570 2414.780 ;
        RECT 2523.170 2414.720 2523.490 2414.780 ;
        RECT 2521.790 2332.100 2522.110 2332.360 ;
        RECT 2521.880 2331.960 2522.020 2332.100 ;
        RECT 2522.250 2331.960 2522.570 2332.020 ;
        RECT 2521.880 2331.820 2522.570 2331.960 ;
        RECT 2522.250 2331.760 2522.570 2331.820 ;
        RECT 2520.870 2318.360 2521.190 2318.420 ;
        RECT 2522.250 2318.360 2522.570 2318.420 ;
        RECT 2520.870 2318.220 2522.570 2318.360 ;
        RECT 2520.870 2318.160 2521.190 2318.220 ;
        RECT 2522.250 2318.160 2522.570 2318.220 ;
        RECT 2521.805 2221.800 2522.095 2221.845 ;
        RECT 2522.250 2221.800 2522.570 2221.860 ;
        RECT 2521.805 2221.660 2522.570 2221.800 ;
        RECT 2521.805 2221.615 2522.095 2221.660 ;
        RECT 2522.250 2221.600 2522.570 2221.660 ;
        RECT 2521.790 2173.860 2522.110 2173.920 ;
        RECT 2521.595 2173.720 2522.110 2173.860 ;
        RECT 2521.790 2173.660 2522.110 2173.720 ;
        RECT 2521.790 2138.980 2522.110 2139.240 ;
        RECT 2521.880 2138.840 2522.020 2138.980 ;
        RECT 2522.250 2138.840 2522.570 2138.900 ;
        RECT 2521.880 2138.700 2522.570 2138.840 ;
        RECT 2522.250 2138.640 2522.570 2138.700 ;
        RECT 2521.805 2125.240 2522.095 2125.285 ;
        RECT 2522.250 2125.240 2522.570 2125.300 ;
        RECT 2521.805 2125.100 2522.570 2125.240 ;
        RECT 2521.805 2125.055 2522.095 2125.100 ;
        RECT 2522.250 2125.040 2522.570 2125.100 ;
        RECT 2521.790 2077.300 2522.110 2077.360 ;
        RECT 2521.595 2077.160 2522.110 2077.300 ;
        RECT 2521.790 2077.100 2522.110 2077.160 ;
        RECT 2521.790 2042.420 2522.110 2042.680 ;
        RECT 2521.880 2041.940 2522.020 2042.420 ;
        RECT 2522.250 2041.940 2522.570 2042.000 ;
        RECT 2521.880 2041.800 2522.570 2041.940 ;
        RECT 2522.250 2041.740 2522.570 2041.800 ;
        RECT 2522.250 2004.540 2522.570 2004.600 ;
        RECT 2523.170 2004.540 2523.490 2004.600 ;
        RECT 2522.250 2004.400 2523.490 2004.540 ;
        RECT 2522.250 2004.340 2522.570 2004.400 ;
        RECT 2523.170 2004.340 2523.490 2004.400 ;
        RECT 2521.790 1966.460 2522.110 1966.520 ;
        RECT 2522.250 1966.460 2522.570 1966.520 ;
        RECT 2521.790 1966.320 2522.570 1966.460 ;
        RECT 2521.790 1966.260 2522.110 1966.320 ;
        RECT 2522.250 1966.260 2522.570 1966.320 ;
        RECT 2522.250 1835.220 2522.570 1835.280 ;
        RECT 2521.880 1835.080 2522.570 1835.220 ;
        RECT 2521.880 1834.940 2522.020 1835.080 ;
        RECT 2522.250 1835.020 2522.570 1835.080 ;
        RECT 2521.790 1834.680 2522.110 1834.940 ;
        RECT 2521.790 1573.420 2522.110 1573.480 ;
        RECT 2522.250 1573.420 2522.570 1573.480 ;
        RECT 2521.790 1573.280 2522.570 1573.420 ;
        RECT 2521.790 1573.220 2522.110 1573.280 ;
        RECT 2522.250 1573.220 2522.570 1573.280 ;
        RECT 2521.790 969.240 2522.110 969.300 ;
        RECT 2576.070 969.240 2576.390 969.300 ;
        RECT 2521.790 969.100 2576.390 969.240 ;
        RECT 2521.790 969.040 2522.110 969.100 ;
        RECT 2576.070 969.040 2576.390 969.100 ;
        RECT 2405.410 33.560 2405.730 33.620 ;
        RECT 2576.070 33.560 2576.390 33.620 ;
        RECT 2405.410 33.420 2576.390 33.560 ;
        RECT 2405.410 33.360 2405.730 33.420 ;
        RECT 2576.070 33.360 2576.390 33.420 ;
      LAYER via ;
        RECT 2297.800 3008.700 2298.060 3008.960 ;
        RECT 2521.820 2980.820 2522.080 2981.080 ;
        RECT 2521.820 2891.060 2522.080 2891.320 ;
        RECT 2522.280 2891.060 2522.540 2891.320 ;
        RECT 2521.820 2863.860 2522.080 2864.120 ;
        RECT 2521.360 2863.180 2521.620 2863.440 ;
        RECT 2521.820 2814.560 2522.080 2814.820 ;
        RECT 2522.740 2814.560 2523.000 2814.820 ;
        RECT 2522.280 2670.740 2522.540 2671.000 ;
        RECT 2521.820 2656.460 2522.080 2656.720 ;
        RECT 2522.280 2656.120 2522.540 2656.380 ;
        RECT 2522.280 2621.440 2522.540 2621.700 ;
        RECT 2521.820 2573.840 2522.080 2574.100 ;
        RECT 2521.820 2559.900 2522.080 2560.160 ;
        RECT 2521.820 2525.560 2522.080 2525.820 ;
        RECT 2522.280 2524.880 2522.540 2525.140 ;
        RECT 2520.900 2487.480 2521.160 2487.740 ;
        RECT 2521.820 2487.480 2522.080 2487.740 ;
        RECT 2521.820 2429.000 2522.080 2429.260 ;
        RECT 2522.280 2428.320 2522.540 2428.580 ;
        RECT 2522.280 2414.720 2522.540 2414.980 ;
        RECT 2523.200 2414.720 2523.460 2414.980 ;
        RECT 2521.820 2332.100 2522.080 2332.360 ;
        RECT 2522.280 2331.760 2522.540 2332.020 ;
        RECT 2520.900 2318.160 2521.160 2318.420 ;
        RECT 2522.280 2318.160 2522.540 2318.420 ;
        RECT 2522.280 2221.600 2522.540 2221.860 ;
        RECT 2521.820 2173.660 2522.080 2173.920 ;
        RECT 2521.820 2138.980 2522.080 2139.240 ;
        RECT 2522.280 2138.640 2522.540 2138.900 ;
        RECT 2522.280 2125.040 2522.540 2125.300 ;
        RECT 2521.820 2077.100 2522.080 2077.360 ;
        RECT 2521.820 2042.420 2522.080 2042.680 ;
        RECT 2522.280 2041.740 2522.540 2042.000 ;
        RECT 2522.280 2004.340 2522.540 2004.600 ;
        RECT 2523.200 2004.340 2523.460 2004.600 ;
        RECT 2521.820 1966.260 2522.080 1966.520 ;
        RECT 2522.280 1966.260 2522.540 1966.520 ;
        RECT 2522.280 1835.020 2522.540 1835.280 ;
        RECT 2521.820 1834.680 2522.080 1834.940 ;
        RECT 2521.820 1573.220 2522.080 1573.480 ;
        RECT 2522.280 1573.220 2522.540 1573.480 ;
        RECT 2521.820 969.040 2522.080 969.300 ;
        RECT 2576.100 969.040 2576.360 969.300 ;
        RECT 2405.440 33.360 2405.700 33.620 ;
        RECT 2576.100 33.360 2576.360 33.620 ;
      LAYER met2 ;
        RECT 2297.010 3008.730 2297.290 3010.000 ;
        RECT 2297.800 3008.730 2298.060 3008.990 ;
        RECT 2297.010 3008.670 2298.060 3008.730 ;
        RECT 2297.010 3008.590 2298.000 3008.670 ;
        RECT 2297.010 3006.000 2297.290 3008.590 ;
        RECT 2521.820 2980.790 2522.080 2981.110 ;
        RECT 2521.880 2963.850 2522.020 2980.790 ;
        RECT 2521.880 2963.710 2522.480 2963.850 ;
        RECT 2522.340 2891.350 2522.480 2963.710 ;
        RECT 2521.820 2891.030 2522.080 2891.350 ;
        RECT 2522.280 2891.030 2522.540 2891.350 ;
        RECT 2521.880 2864.150 2522.020 2891.030 ;
        RECT 2521.820 2863.830 2522.080 2864.150 ;
        RECT 2521.360 2863.150 2521.620 2863.470 ;
        RECT 2521.420 2849.610 2521.560 2863.150 ;
        RECT 2521.810 2849.610 2522.090 2849.725 ;
        RECT 2521.420 2849.470 2522.090 2849.610 ;
        RECT 2521.810 2849.355 2522.090 2849.470 ;
        RECT 2522.730 2849.355 2523.010 2849.725 ;
        RECT 2522.800 2814.850 2522.940 2849.355 ;
        RECT 2521.820 2814.530 2522.080 2814.850 ;
        RECT 2522.740 2814.530 2523.000 2814.850 ;
        RECT 2521.880 2719.050 2522.020 2814.530 ;
        RECT 2521.880 2718.910 2522.480 2719.050 ;
        RECT 2522.340 2671.030 2522.480 2718.910 ;
        RECT 2522.280 2670.710 2522.540 2671.030 ;
        RECT 2521.880 2656.750 2522.020 2656.905 ;
        RECT 2521.820 2656.490 2522.080 2656.750 ;
        RECT 2521.820 2656.430 2522.480 2656.490 ;
        RECT 2521.880 2656.410 2522.480 2656.430 ;
        RECT 2521.880 2656.350 2522.540 2656.410 ;
        RECT 2522.280 2656.090 2522.540 2656.350 ;
        RECT 2522.280 2621.410 2522.540 2621.730 ;
        RECT 2522.340 2608.210 2522.480 2621.410 ;
        RECT 2521.880 2608.070 2522.480 2608.210 ;
        RECT 2521.880 2574.130 2522.020 2608.070 ;
        RECT 2521.820 2573.810 2522.080 2574.130 ;
        RECT 2521.820 2559.870 2522.080 2560.190 ;
        RECT 2521.880 2525.850 2522.020 2559.870 ;
        RECT 2521.820 2525.530 2522.080 2525.850 ;
        RECT 2522.280 2524.850 2522.540 2525.170 ;
        RECT 2522.340 2511.650 2522.480 2524.850 ;
        RECT 2521.880 2511.510 2522.480 2511.650 ;
        RECT 2521.880 2487.770 2522.020 2511.510 ;
        RECT 2520.900 2487.450 2521.160 2487.770 ;
        RECT 2521.820 2487.450 2522.080 2487.770 ;
        RECT 2520.960 2463.485 2521.100 2487.450 ;
        RECT 2520.890 2463.115 2521.170 2463.485 ;
        RECT 2521.810 2463.115 2522.090 2463.485 ;
        RECT 2521.880 2429.290 2522.020 2463.115 ;
        RECT 2521.820 2428.970 2522.080 2429.290 ;
        RECT 2522.280 2428.290 2522.540 2428.610 ;
        RECT 2522.340 2415.010 2522.480 2428.290 ;
        RECT 2522.280 2414.690 2522.540 2415.010 ;
        RECT 2523.200 2414.690 2523.460 2415.010 ;
        RECT 2523.260 2366.925 2523.400 2414.690 ;
        RECT 2522.270 2366.810 2522.550 2366.925 ;
        RECT 2521.880 2366.670 2522.550 2366.810 ;
        RECT 2521.880 2332.390 2522.020 2366.670 ;
        RECT 2522.270 2366.555 2522.550 2366.670 ;
        RECT 2523.190 2366.555 2523.470 2366.925 ;
        RECT 2521.820 2332.070 2522.080 2332.390 ;
        RECT 2522.280 2331.730 2522.540 2332.050 ;
        RECT 2522.340 2318.450 2522.480 2331.730 ;
        RECT 2520.900 2318.130 2521.160 2318.450 ;
        RECT 2522.280 2318.130 2522.540 2318.450 ;
        RECT 2520.960 2270.365 2521.100 2318.130 ;
        RECT 2520.890 2269.995 2521.170 2270.365 ;
        RECT 2521.810 2269.995 2522.090 2270.365 ;
        RECT 2521.880 2234.890 2522.020 2269.995 ;
        RECT 2521.880 2234.750 2522.480 2234.890 ;
        RECT 2522.340 2221.890 2522.480 2234.750 ;
        RECT 2522.280 2221.570 2522.540 2221.890 ;
        RECT 2521.820 2173.630 2522.080 2173.950 ;
        RECT 2521.880 2139.270 2522.020 2173.630 ;
        RECT 2521.820 2138.950 2522.080 2139.270 ;
        RECT 2522.280 2138.610 2522.540 2138.930 ;
        RECT 2522.340 2125.330 2522.480 2138.610 ;
        RECT 2522.280 2125.010 2522.540 2125.330 ;
        RECT 2521.820 2077.070 2522.080 2077.390 ;
        RECT 2521.880 2042.710 2522.020 2077.070 ;
        RECT 2521.820 2042.390 2522.080 2042.710 ;
        RECT 2522.280 2041.710 2522.540 2042.030 ;
        RECT 2522.340 2004.630 2522.480 2041.710 ;
        RECT 2522.280 2004.310 2522.540 2004.630 ;
        RECT 2523.200 2004.310 2523.460 2004.630 ;
        RECT 2523.260 1980.685 2523.400 2004.310 ;
        RECT 2522.270 1980.570 2522.550 1980.685 ;
        RECT 2521.880 1980.430 2522.550 1980.570 ;
        RECT 2521.880 1966.550 2522.020 1980.430 ;
        RECT 2522.270 1980.315 2522.550 1980.430 ;
        RECT 2523.190 1980.315 2523.470 1980.685 ;
        RECT 2521.820 1966.230 2522.080 1966.550 ;
        RECT 2522.280 1966.230 2522.540 1966.550 ;
        RECT 2522.340 1835.310 2522.480 1966.230 ;
        RECT 2522.280 1834.990 2522.540 1835.310 ;
        RECT 2521.820 1834.650 2522.080 1834.970 ;
        RECT 2521.880 1725.400 2522.020 1834.650 ;
        RECT 2521.880 1725.260 2522.480 1725.400 ;
        RECT 2522.340 1629.010 2522.480 1725.260 ;
        RECT 2522.340 1628.870 2522.940 1629.010 ;
        RECT 2522.800 1628.330 2522.940 1628.870 ;
        RECT 2522.340 1628.190 2522.940 1628.330 ;
        RECT 2522.340 1573.510 2522.480 1628.190 ;
        RECT 2521.820 1573.190 2522.080 1573.510 ;
        RECT 2522.280 1573.190 2522.540 1573.510 ;
        RECT 2521.880 1535.170 2522.020 1573.190 ;
        RECT 2521.880 1535.030 2522.480 1535.170 ;
        RECT 2522.340 1466.490 2522.480 1535.030 ;
        RECT 2521.880 1466.350 2522.480 1466.490 ;
        RECT 2521.880 969.330 2522.020 1466.350 ;
        RECT 2521.820 969.010 2522.080 969.330 ;
        RECT 2576.100 969.010 2576.360 969.330 ;
        RECT 2576.160 33.650 2576.300 969.010 ;
        RECT 2405.440 33.330 2405.700 33.650 ;
        RECT 2576.100 33.330 2576.360 33.650 ;
        RECT 2405.500 2.400 2405.640 33.330 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
      LAYER via2 ;
        RECT 2521.810 2849.400 2522.090 2849.680 ;
        RECT 2522.730 2849.400 2523.010 2849.680 ;
        RECT 2520.890 2463.160 2521.170 2463.440 ;
        RECT 2521.810 2463.160 2522.090 2463.440 ;
        RECT 2522.270 2366.600 2522.550 2366.880 ;
        RECT 2523.190 2366.600 2523.470 2366.880 ;
        RECT 2520.890 2270.040 2521.170 2270.320 ;
        RECT 2521.810 2270.040 2522.090 2270.320 ;
        RECT 2522.270 1980.360 2522.550 1980.640 ;
        RECT 2523.190 1980.360 2523.470 1980.640 ;
      LAYER met3 ;
        RECT 2521.785 2849.690 2522.115 2849.705 ;
        RECT 2522.705 2849.690 2523.035 2849.705 ;
        RECT 2521.785 2849.390 2523.035 2849.690 ;
        RECT 2521.785 2849.375 2522.115 2849.390 ;
        RECT 2522.705 2849.375 2523.035 2849.390 ;
        RECT 2520.865 2463.450 2521.195 2463.465 ;
        RECT 2521.785 2463.450 2522.115 2463.465 ;
        RECT 2520.865 2463.150 2522.115 2463.450 ;
        RECT 2520.865 2463.135 2521.195 2463.150 ;
        RECT 2521.785 2463.135 2522.115 2463.150 ;
        RECT 2522.245 2366.890 2522.575 2366.905 ;
        RECT 2523.165 2366.890 2523.495 2366.905 ;
        RECT 2522.245 2366.590 2523.495 2366.890 ;
        RECT 2522.245 2366.575 2522.575 2366.590 ;
        RECT 2523.165 2366.575 2523.495 2366.590 ;
        RECT 2520.865 2270.330 2521.195 2270.345 ;
        RECT 2521.785 2270.330 2522.115 2270.345 ;
        RECT 2520.865 2270.030 2522.115 2270.330 ;
        RECT 2520.865 2270.015 2521.195 2270.030 ;
        RECT 2521.785 2270.015 2522.115 2270.030 ;
        RECT 2522.245 1980.650 2522.575 1980.665 ;
        RECT 2523.165 1980.650 2523.495 1980.665 ;
        RECT 2522.245 1980.350 2523.495 1980.650 ;
        RECT 2522.245 1980.335 2522.575 1980.350 ;
        RECT 2523.165 1980.335 2523.495 1980.350 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 302.750 3015.700 303.070 3015.760 ;
        RECT 443.970 3015.700 444.290 3015.760 ;
        RECT 302.750 3015.560 444.290 3015.700 ;
        RECT 302.750 3015.500 303.070 3015.560 ;
        RECT 443.970 3015.500 444.290 3015.560 ;
        RECT 302.750 33.900 303.070 33.960 ;
        RECT 799.550 33.900 799.870 33.960 ;
        RECT 302.750 33.760 799.870 33.900 ;
        RECT 302.750 33.700 303.070 33.760 ;
        RECT 799.550 33.700 799.870 33.760 ;
      LAYER via ;
        RECT 302.780 3015.500 303.040 3015.760 ;
        RECT 444.000 3015.500 444.260 3015.760 ;
        RECT 302.780 33.700 303.040 33.960 ;
        RECT 799.580 33.700 799.840 33.960 ;
      LAYER met2 ;
        RECT 302.780 3015.470 303.040 3015.790 ;
        RECT 444.000 3015.470 444.260 3015.790 ;
        RECT 302.840 33.990 302.980 3015.470 ;
        RECT 444.060 3010.000 444.200 3015.470 ;
        RECT 444.060 3009.340 444.410 3010.000 ;
        RECT 444.130 3006.000 444.410 3009.340 ;
        RECT 302.780 33.670 303.040 33.990 ;
        RECT 799.580 33.670 799.840 33.990 ;
        RECT 799.640 2.400 799.780 33.670 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 404.870 507.520 405.190 507.580 ;
        RECT 641.770 507.520 642.090 507.580 ;
        RECT 404.870 507.380 642.090 507.520 ;
        RECT 404.870 507.320 405.190 507.380 ;
        RECT 641.770 507.320 642.090 507.380 ;
        RECT 641.770 2.960 642.090 3.020 ;
        RECT 644.990 2.960 645.310 3.020 ;
        RECT 641.770 2.820 645.310 2.960 ;
        RECT 641.770 2.760 642.090 2.820 ;
        RECT 644.990 2.760 645.310 2.820 ;
      LAYER via ;
        RECT 404.900 507.320 405.160 507.580 ;
        RECT 641.800 507.320 642.060 507.580 ;
        RECT 641.800 2.760 642.060 3.020 ;
        RECT 645.020 2.760 645.280 3.020 ;
      LAYER met2 ;
        RECT 404.890 2412.795 405.170 2413.165 ;
        RECT 404.960 507.610 405.100 2412.795 ;
        RECT 404.900 507.290 405.160 507.610 ;
        RECT 641.800 507.290 642.060 507.610 ;
        RECT 641.860 3.050 642.000 507.290 ;
        RECT 641.800 2.730 642.060 3.050 ;
        RECT 645.020 2.730 645.280 3.050 ;
        RECT 645.080 2.400 645.220 2.730 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 404.890 2412.840 405.170 2413.120 ;
      LAYER met3 ;
        RECT 404.865 2413.130 405.195 2413.145 ;
        RECT 410.000 2413.130 414.000 2413.280 ;
        RECT 404.865 2412.830 414.000 2413.130 ;
        RECT 404.865 2412.815 405.195 2412.830 ;
        RECT 410.000 2412.680 414.000 2412.830 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2366.980 2519.810 2367.040 ;
        RECT 2616.550 2366.980 2616.870 2367.040 ;
        RECT 2519.490 2366.840 2616.870 2366.980 ;
        RECT 2519.490 2366.780 2519.810 2366.840 ;
        RECT 2616.550 2366.780 2616.870 2366.840 ;
        RECT 2434.850 496.300 2435.170 496.360 ;
        RECT 2616.550 496.300 2616.870 496.360 ;
        RECT 2434.850 496.160 2616.870 496.300 ;
        RECT 2434.850 496.100 2435.170 496.160 ;
        RECT 2616.550 496.100 2616.870 496.160 ;
        RECT 2428.870 20.300 2429.190 20.360 ;
        RECT 2434.850 20.300 2435.170 20.360 ;
        RECT 2428.870 20.160 2435.170 20.300 ;
        RECT 2428.870 20.100 2429.190 20.160 ;
        RECT 2434.850 20.100 2435.170 20.160 ;
      LAYER via ;
        RECT 2519.520 2366.780 2519.780 2367.040 ;
        RECT 2616.580 2366.780 2616.840 2367.040 ;
        RECT 2434.880 496.100 2435.140 496.360 ;
        RECT 2616.580 496.100 2616.840 496.360 ;
        RECT 2428.900 20.100 2429.160 20.360 ;
        RECT 2434.880 20.100 2435.140 20.360 ;
      LAYER met2 ;
        RECT 2519.520 2366.925 2519.780 2367.070 ;
        RECT 2519.510 2366.555 2519.790 2366.925 ;
        RECT 2616.580 2366.750 2616.840 2367.070 ;
        RECT 2616.640 496.390 2616.780 2366.750 ;
        RECT 2434.880 496.070 2435.140 496.390 ;
        RECT 2616.580 496.070 2616.840 496.390 ;
        RECT 2434.940 20.390 2435.080 496.070 ;
        RECT 2428.900 20.070 2429.160 20.390 ;
        RECT 2434.880 20.070 2435.140 20.390 ;
        RECT 2428.960 2.400 2429.100 20.070 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2366.600 2519.790 2366.880 ;
      LAYER met3 ;
        RECT 2506.000 2366.890 2510.000 2367.040 ;
        RECT 2519.485 2366.890 2519.815 2366.905 ;
        RECT 2506.000 2366.590 2519.815 2366.890 ;
        RECT 2506.000 2366.440 2510.000 2366.590 ;
        RECT 2519.485 2366.575 2519.815 2366.590 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.950 3010.515 1445.230 3010.885 ;
        RECT 1445.020 3010.000 1445.160 3010.515 ;
        RECT 1445.020 3009.340 1445.370 3010.000 ;
        RECT 1445.090 3006.000 1445.370 3009.340 ;
        RECT 2446.830 19.875 2447.110 20.245 ;
        RECT 2446.900 2.400 2447.040 19.875 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
      LAYER via2 ;
        RECT 1444.950 3010.560 1445.230 3010.840 ;
        RECT 2446.830 19.920 2447.110 20.200 ;
      LAYER met3 ;
        RECT 1444.925 3010.850 1445.255 3010.865 ;
        RECT 2442.870 3010.850 2443.250 3010.860 ;
        RECT 1444.925 3010.550 2443.250 3010.850 ;
        RECT 1444.925 3010.535 1445.255 3010.550 ;
        RECT 2442.870 3010.540 2443.250 3010.550 ;
        RECT 2442.870 20.210 2443.250 20.220 ;
        RECT 2446.805 20.210 2447.135 20.225 ;
        RECT 2442.870 19.910 2447.135 20.210 ;
        RECT 2442.870 19.900 2443.250 19.910 ;
        RECT 2446.805 19.895 2447.135 19.910 ;
      LAYER via3 ;
        RECT 2442.900 3010.540 2443.220 3010.860 ;
        RECT 2442.900 19.900 2443.220 20.220 ;
      LAYER met4 ;
        RECT 2442.895 3010.535 2443.225 3010.865 ;
        RECT 2442.910 1878.650 2443.210 3010.535 ;
        RECT 2441.990 1878.350 2443.210 1878.650 ;
        RECT 2441.990 1868.450 2442.290 1878.350 ;
        RECT 2441.990 1868.150 2445.050 1868.450 ;
        RECT 2444.750 1841.250 2445.050 1868.150 ;
        RECT 2442.910 1840.950 2445.050 1841.250 ;
        RECT 2442.910 977.650 2443.210 1840.950 ;
        RECT 2442.910 977.350 2445.050 977.650 ;
        RECT 2444.750 970.850 2445.050 977.350 ;
        RECT 2442.910 970.550 2445.050 970.850 ;
        RECT 2442.910 20.225 2443.210 970.550 ;
        RECT 2442.895 19.895 2443.225 20.225 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.510 210.700 1179.830 210.760 ;
        RECT 2463.370 210.700 2463.690 210.760 ;
        RECT 1179.510 210.560 2463.690 210.700 ;
        RECT 1179.510 210.500 1179.830 210.560 ;
        RECT 2463.370 210.500 2463.690 210.560 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2463.370 2.820 2465.070 2.960 ;
        RECT 2463.370 2.760 2463.690 2.820 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
      LAYER via ;
        RECT 1179.540 210.500 1179.800 210.760 ;
        RECT 2463.400 210.500 2463.660 210.760 ;
        RECT 2463.400 2.760 2463.660 3.020 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
      LAYER met2 ;
        RECT 1178.290 510.410 1178.570 514.000 ;
        RECT 1178.290 510.270 1179.740 510.410 ;
        RECT 1178.290 510.000 1178.570 510.270 ;
        RECT 1179.600 210.790 1179.740 510.270 ;
        RECT 1179.540 210.470 1179.800 210.790 ;
        RECT 2463.400 210.470 2463.660 210.790 ;
        RECT 2463.460 3.050 2463.600 210.470 ;
        RECT 2463.400 2.730 2463.660 3.050 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.150 168.880 1241.470 168.940 ;
        RECT 2477.170 168.880 2477.490 168.940 ;
        RECT 1241.150 168.740 2477.490 168.880 ;
        RECT 1241.150 168.680 1241.470 168.740 ;
        RECT 2477.170 168.680 2477.490 168.740 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1241.180 168.680 1241.440 168.940 ;
        RECT 2477.200 168.680 2477.460 168.940 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1239.930 510.410 1240.210 514.000 ;
        RECT 1239.930 510.270 1241.380 510.410 ;
        RECT 1239.930 510.000 1240.210 510.270 ;
        RECT 1241.240 168.970 1241.380 510.270 ;
        RECT 1241.180 168.650 1241.440 168.970 ;
        RECT 2477.200 168.650 2477.460 168.970 ;
        RECT 2477.260 3.050 2477.400 168.650 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1904.580 2519.810 1904.640 ;
        RECT 2595.850 1904.580 2596.170 1904.640 ;
        RECT 2519.490 1904.440 2596.170 1904.580 ;
        RECT 2519.490 1904.380 2519.810 1904.440 ;
        RECT 2595.850 1904.380 2596.170 1904.440 ;
        RECT 2504.310 507.180 2504.630 507.240 ;
        RECT 2595.850 507.180 2596.170 507.240 ;
        RECT 2504.310 507.040 2596.170 507.180 ;
        RECT 2504.310 506.980 2504.630 507.040 ;
        RECT 2595.850 506.980 2596.170 507.040 ;
        RECT 2500.630 19.620 2500.950 19.680 ;
        RECT 2504.310 19.620 2504.630 19.680 ;
        RECT 2500.630 19.480 2504.630 19.620 ;
        RECT 2500.630 19.420 2500.950 19.480 ;
        RECT 2504.310 19.420 2504.630 19.480 ;
      LAYER via ;
        RECT 2519.520 1904.380 2519.780 1904.640 ;
        RECT 2595.880 1904.380 2596.140 1904.640 ;
        RECT 2504.340 506.980 2504.600 507.240 ;
        RECT 2595.880 506.980 2596.140 507.240 ;
        RECT 2500.660 19.420 2500.920 19.680 ;
        RECT 2504.340 19.420 2504.600 19.680 ;
      LAYER met2 ;
        RECT 2519.510 1909.595 2519.790 1909.965 ;
        RECT 2519.580 1904.670 2519.720 1909.595 ;
        RECT 2519.520 1904.350 2519.780 1904.670 ;
        RECT 2595.880 1904.350 2596.140 1904.670 ;
        RECT 2595.940 507.270 2596.080 1904.350 ;
        RECT 2504.340 506.950 2504.600 507.270 ;
        RECT 2595.880 506.950 2596.140 507.270 ;
        RECT 2504.400 19.710 2504.540 506.950 ;
        RECT 2500.660 19.390 2500.920 19.710 ;
        RECT 2504.340 19.390 2504.600 19.710 ;
        RECT 2500.720 2.400 2500.860 19.390 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 2519.510 1909.640 2519.790 1909.920 ;
      LAYER met3 ;
        RECT 2506.000 1909.930 2510.000 1910.080 ;
        RECT 2519.485 1909.930 2519.815 1909.945 ;
        RECT 2506.000 1909.630 2519.815 1909.930 ;
        RECT 2506.000 1909.480 2510.000 1909.630 ;
        RECT 2519.485 1909.615 2519.815 1909.630 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2512.130 23.360 2512.450 23.420 ;
        RECT 2518.110 23.360 2518.430 23.420 ;
        RECT 2512.130 23.220 2518.430 23.360 ;
        RECT 2512.130 23.160 2512.450 23.220 ;
        RECT 2518.110 23.160 2518.430 23.220 ;
      LAYER via ;
        RECT 2512.160 23.160 2512.420 23.420 ;
        RECT 2518.140 23.160 2518.400 23.420 ;
      LAYER met2 ;
        RECT 2512.150 1562.795 2512.430 1563.165 ;
        RECT 2512.220 23.450 2512.360 1562.795 ;
        RECT 2512.160 23.130 2512.420 23.450 ;
        RECT 2518.140 23.130 2518.400 23.450 ;
        RECT 2518.200 2.400 2518.340 23.130 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
      LAYER via2 ;
        RECT 2512.150 1562.840 2512.430 1563.120 ;
      LAYER met3 ;
        RECT 2506.000 1563.130 2510.000 1563.280 ;
        RECT 2512.125 1563.130 2512.455 1563.145 ;
        RECT 2506.000 1562.830 2512.455 1563.130 ;
        RECT 2506.000 1562.680 2510.000 1562.830 ;
        RECT 2512.125 1562.815 2512.455 1562.830 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.510 300.120 489.830 300.180 ;
        RECT 2521.790 300.120 2522.110 300.180 ;
        RECT 489.510 299.980 2522.110 300.120 ;
        RECT 489.510 299.920 489.830 299.980 ;
        RECT 2521.790 299.920 2522.110 299.980 ;
        RECT 2521.790 15.200 2522.110 15.260 ;
        RECT 2536.050 15.200 2536.370 15.260 ;
        RECT 2521.790 15.060 2536.370 15.200 ;
        RECT 2521.790 15.000 2522.110 15.060 ;
        RECT 2536.050 15.000 2536.370 15.060 ;
      LAYER via ;
        RECT 489.540 299.920 489.800 300.180 ;
        RECT 2521.820 299.920 2522.080 300.180 ;
        RECT 2521.820 15.000 2522.080 15.260 ;
        RECT 2536.080 15.000 2536.340 15.260 ;
      LAYER met2 ;
        RECT 486.450 510.410 486.730 514.000 ;
        RECT 486.450 510.270 489.740 510.410 ;
        RECT 486.450 510.000 486.730 510.270 ;
        RECT 489.600 300.210 489.740 510.270 ;
        RECT 489.540 299.890 489.800 300.210 ;
        RECT 2521.820 299.890 2522.080 300.210 ;
        RECT 2521.880 15.290 2522.020 299.890 ;
        RECT 2521.820 14.970 2522.080 15.290 ;
        RECT 2536.080 14.970 2536.340 15.290 ;
        RECT 2536.140 2.400 2536.280 14.970 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 46.140 1366.130 46.200 ;
        RECT 2553.990 46.140 2554.310 46.200 ;
        RECT 1365.810 46.000 2554.310 46.140 ;
        RECT 1365.810 45.940 1366.130 46.000 ;
        RECT 2553.990 45.940 2554.310 46.000 ;
      LAYER via ;
        RECT 1365.840 45.940 1366.100 46.200 ;
        RECT 2554.020 45.940 2554.280 46.200 ;
      LAYER met2 ;
        RECT 1363.210 510.410 1363.490 514.000 ;
        RECT 1363.210 510.270 1366.040 510.410 ;
        RECT 1363.210 510.000 1363.490 510.270 ;
        RECT 1365.900 46.230 1366.040 510.270 ;
        RECT 1365.840 45.910 1366.100 46.230 ;
        RECT 2554.020 45.910 2554.280 46.230 ;
        RECT 2554.080 2.400 2554.220 45.910 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2470.340 2519.810 2470.400 ;
        RECT 2568.250 2470.340 2568.570 2470.400 ;
        RECT 2519.490 2470.200 2568.570 2470.340 ;
        RECT 2519.490 2470.140 2519.810 2470.200 ;
        RECT 2568.250 2470.140 2568.570 2470.200 ;
        RECT 2568.250 2.960 2568.570 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2568.250 2.820 2572.250 2.960 ;
        RECT 2568.250 2.760 2568.570 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 2519.520 2470.140 2519.780 2470.400 ;
        RECT 2568.280 2470.140 2568.540 2470.400 ;
        RECT 2568.280 2.760 2568.540 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 2519.510 2475.355 2519.790 2475.725 ;
        RECT 2519.580 2470.430 2519.720 2475.355 ;
        RECT 2519.520 2470.110 2519.780 2470.430 ;
        RECT 2568.280 2470.110 2568.540 2470.430 ;
        RECT 2568.340 3.050 2568.480 2470.110 ;
        RECT 2568.280 2.730 2568.540 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2475.400 2519.790 2475.680 ;
      LAYER met3 ;
        RECT 2506.000 2475.690 2510.000 2475.840 ;
        RECT 2519.485 2475.690 2519.815 2475.705 ;
        RECT 2506.000 2475.390 2519.815 2475.690 ;
        RECT 2506.000 2475.240 2510.000 2475.390 ;
        RECT 2519.485 2475.375 2519.815 2475.390 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.770 3009.410 1334.050 3010.000 ;
        RECT 1335.470 3009.410 1335.750 3009.525 ;
        RECT 1333.770 3009.270 1335.750 3009.410 ;
        RECT 1333.770 3006.000 1334.050 3009.270 ;
        RECT 1335.470 3009.155 1335.750 3009.270 ;
        RECT 2587.590 3009.155 2587.870 3009.525 ;
        RECT 2587.660 17.410 2587.800 3009.155 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
      LAYER via2 ;
        RECT 1335.470 3009.200 1335.750 3009.480 ;
        RECT 2587.590 3009.200 2587.870 3009.480 ;
      LAYER met3 ;
        RECT 1335.445 3009.490 1335.775 3009.505 ;
        RECT 2587.565 3009.490 2587.895 3009.505 ;
        RECT 1335.445 3009.190 2587.895 3009.490 ;
        RECT 1335.445 3009.175 1335.775 3009.190 ;
        RECT 2587.565 3009.175 2587.895 3009.190 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2104.840 2519.810 2104.900 ;
        RECT 2533.290 2104.840 2533.610 2104.900 ;
        RECT 2519.490 2104.700 2533.610 2104.840 ;
        RECT 2519.490 2104.640 2519.810 2104.700 ;
        RECT 2533.290 2104.640 2533.610 2104.700 ;
        RECT 827.610 314.060 827.930 314.120 ;
        RECT 2533.290 314.060 2533.610 314.120 ;
        RECT 827.610 313.920 2533.610 314.060 ;
        RECT 827.610 313.860 827.930 313.920 ;
        RECT 2533.290 313.860 2533.610 313.920 ;
        RECT 823.470 15.200 823.790 15.260 ;
        RECT 827.610 15.200 827.930 15.260 ;
        RECT 823.470 15.060 827.930 15.200 ;
        RECT 823.470 15.000 823.790 15.060 ;
        RECT 827.610 15.000 827.930 15.060 ;
      LAYER via ;
        RECT 2519.520 2104.640 2519.780 2104.900 ;
        RECT 2533.320 2104.640 2533.580 2104.900 ;
        RECT 827.640 313.860 827.900 314.120 ;
        RECT 2533.320 313.860 2533.580 314.120 ;
        RECT 823.500 15.000 823.760 15.260 ;
        RECT 827.640 15.000 827.900 15.260 ;
      LAYER met2 ;
        RECT 2519.510 2110.875 2519.790 2111.245 ;
        RECT 2519.580 2104.930 2519.720 2110.875 ;
        RECT 2519.520 2104.610 2519.780 2104.930 ;
        RECT 2533.320 2104.610 2533.580 2104.930 ;
        RECT 2533.380 314.150 2533.520 2104.610 ;
        RECT 827.640 313.830 827.900 314.150 ;
        RECT 2533.320 313.830 2533.580 314.150 ;
        RECT 827.700 15.290 827.840 313.830 ;
        RECT 823.500 14.970 823.760 15.290 ;
        RECT 827.640 14.970 827.900 15.290 ;
        RECT 823.560 2.400 823.700 14.970 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2110.920 2519.790 2111.200 ;
      LAYER met3 ;
        RECT 2506.000 2111.210 2510.000 2111.360 ;
        RECT 2519.485 2111.210 2519.815 2111.225 ;
        RECT 2506.000 2110.910 2519.815 2111.210 ;
        RECT 2506.000 2110.760 2510.000 2110.910 ;
        RECT 2519.485 2110.895 2519.815 2110.910 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.410 3010.260 1347.730 3010.320 ;
        RECT 2409.090 3010.260 2409.410 3010.320 ;
        RECT 1347.410 3010.120 2409.410 3010.260 ;
        RECT 1347.410 3010.060 1347.730 3010.120 ;
        RECT 2409.090 3010.060 2409.410 3010.120 ;
        RECT 2601.370 17.920 2601.690 17.980 ;
        RECT 2607.350 17.920 2607.670 17.980 ;
        RECT 2601.370 17.780 2607.670 17.920 ;
        RECT 2601.370 17.720 2601.690 17.780 ;
        RECT 2607.350 17.720 2607.670 17.780 ;
      LAYER via ;
        RECT 1347.440 3010.060 1347.700 3010.320 ;
        RECT 2409.120 3010.060 2409.380 3010.320 ;
        RECT 2601.400 17.720 2601.660 17.980 ;
        RECT 2607.380 17.720 2607.640 17.980 ;
      LAYER met2 ;
        RECT 1347.440 3010.030 1347.700 3010.350 ;
        RECT 2409.120 3010.205 2409.380 3010.350 ;
        RECT 1345.730 3009.410 1346.010 3010.000 ;
        RECT 1347.500 3009.410 1347.640 3010.030 ;
        RECT 2409.110 3009.835 2409.390 3010.205 ;
        RECT 2601.390 3009.835 2601.670 3010.205 ;
        RECT 1345.730 3009.270 1347.640 3009.410 ;
        RECT 1345.730 3006.000 1346.010 3009.270 ;
        RECT 2601.460 18.010 2601.600 3009.835 ;
        RECT 2601.400 17.690 2601.660 18.010 ;
        RECT 2607.380 17.690 2607.640 18.010 ;
        RECT 2607.440 2.400 2607.580 17.690 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
      LAYER via2 ;
        RECT 2409.110 3009.880 2409.390 3010.160 ;
        RECT 2601.390 3009.880 2601.670 3010.160 ;
      LAYER met3 ;
        RECT 2409.085 3010.170 2409.415 3010.185 ;
        RECT 2601.365 3010.170 2601.695 3010.185 ;
        RECT 2409.085 3009.870 2601.695 3010.170 ;
        RECT 2409.085 3009.855 2409.415 3009.870 ;
        RECT 2601.365 3009.855 2601.695 3009.870 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1889.290 3010.940 1889.610 3011.000 ;
        RECT 2622.070 3010.940 2622.390 3011.000 ;
        RECT 1889.290 3010.800 2622.390 3010.940 ;
        RECT 1889.290 3010.740 1889.610 3010.800 ;
        RECT 2622.070 3010.740 2622.390 3010.800 ;
      LAYER via ;
        RECT 1889.320 3010.740 1889.580 3011.000 ;
        RECT 2622.100 3010.740 2622.360 3011.000 ;
      LAYER met2 ;
        RECT 1889.320 3010.710 1889.580 3011.030 ;
        RECT 2622.100 3010.710 2622.360 3011.030 ;
        RECT 1889.380 3010.000 1889.520 3010.710 ;
        RECT 1889.380 3009.340 1889.730 3010.000 ;
        RECT 1889.450 3006.000 1889.730 3009.340 ;
        RECT 2622.160 16.730 2622.300 3010.710 ;
        RECT 2622.160 16.590 2625.520 16.730 ;
        RECT 2625.380 2.400 2625.520 16.590 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.970 496.980 1870.290 497.040 ;
        RECT 1876.410 496.980 1876.730 497.040 ;
        RECT 1869.970 496.840 1876.730 496.980 ;
        RECT 1869.970 496.780 1870.290 496.840 ;
        RECT 1876.410 496.780 1876.730 496.840 ;
        RECT 1876.410 74.360 1876.730 74.420 ;
        RECT 2643.230 74.360 2643.550 74.420 ;
        RECT 1876.410 74.220 2643.550 74.360 ;
        RECT 1876.410 74.160 1876.730 74.220 ;
        RECT 2643.230 74.160 2643.550 74.220 ;
      LAYER via ;
        RECT 1870.000 496.780 1870.260 497.040 ;
        RECT 1876.440 496.780 1876.700 497.040 ;
        RECT 1876.440 74.160 1876.700 74.420 ;
        RECT 2643.260 74.160 2643.520 74.420 ;
      LAYER met2 ;
        RECT 1870.130 510.340 1870.410 514.000 ;
        RECT 1870.060 510.000 1870.410 510.340 ;
        RECT 1870.060 497.070 1870.200 510.000 ;
        RECT 1870.000 496.750 1870.260 497.070 ;
        RECT 1876.440 496.750 1876.700 497.070 ;
        RECT 1876.500 74.450 1876.640 496.750 ;
        RECT 1876.440 74.130 1876.700 74.450 ;
        RECT 2643.260 74.130 2643.520 74.450 ;
        RECT 2643.320 2.400 2643.460 74.130 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 100.540 1414.430 100.600 ;
        RECT 2656.570 100.540 2656.890 100.600 ;
        RECT 1414.110 100.400 2656.890 100.540 ;
        RECT 1414.110 100.340 1414.430 100.400 ;
        RECT 2656.570 100.340 2656.890 100.400 ;
      LAYER via ;
        RECT 1414.140 100.340 1414.400 100.600 ;
        RECT 2656.600 100.340 2656.860 100.600 ;
      LAYER met2 ;
        RECT 1412.890 510.410 1413.170 514.000 ;
        RECT 1412.890 510.270 1414.340 510.410 ;
        RECT 1412.890 510.000 1413.170 510.270 ;
        RECT 1414.200 100.630 1414.340 510.270 ;
        RECT 1414.140 100.310 1414.400 100.630 ;
        RECT 2656.600 100.310 2656.860 100.630 ;
        RECT 2656.660 18.090 2656.800 100.310 ;
        RECT 2656.660 17.950 2661.400 18.090 ;
        RECT 2661.260 2.400 2661.400 17.950 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.930 29.820 1008.250 29.880 ;
        RECT 1055.310 29.820 1055.630 29.880 ;
        RECT 1007.930 29.680 1055.630 29.820 ;
        RECT 1007.930 29.620 1008.250 29.680 ;
        RECT 1055.310 29.620 1055.630 29.680 ;
        RECT 2409.090 29.820 2409.410 29.880 ;
        RECT 2456.010 29.820 2456.330 29.880 ;
        RECT 2409.090 29.680 2456.330 29.820 ;
        RECT 2409.090 29.620 2409.410 29.680 ;
        RECT 2456.010 29.620 2456.330 29.680 ;
        RECT 676.270 28.800 676.590 28.860 ;
        RECT 724.110 28.800 724.430 28.860 ;
        RECT 676.270 28.660 724.430 28.800 ;
        RECT 676.270 28.600 676.590 28.660 ;
        RECT 724.110 28.600 724.430 28.660 ;
        RECT 2190.590 28.800 2190.910 28.860 ;
        RECT 2214.510 28.800 2214.830 28.860 ;
        RECT 2190.590 28.660 2214.830 28.800 ;
        RECT 2190.590 28.600 2190.910 28.660 ;
        RECT 2214.510 28.600 2214.830 28.660 ;
        RECT 910.870 28.460 911.190 28.520 ;
        RECT 999.650 28.460 999.970 28.520 ;
        RECT 910.870 28.320 999.970 28.460 ;
        RECT 910.870 28.260 911.190 28.320 ;
        RECT 999.650 28.260 999.970 28.320 ;
      LAYER via ;
        RECT 1007.960 29.620 1008.220 29.880 ;
        RECT 1055.340 29.620 1055.600 29.880 ;
        RECT 2409.120 29.620 2409.380 29.880 ;
        RECT 2456.040 29.620 2456.300 29.880 ;
        RECT 676.300 28.600 676.560 28.860 ;
        RECT 724.140 28.600 724.400 28.860 ;
        RECT 2190.620 28.600 2190.880 28.860 ;
        RECT 2214.540 28.600 2214.800 28.860 ;
        RECT 910.900 28.260 911.160 28.520 ;
        RECT 999.680 28.260 999.940 28.520 ;
      LAYER met2 ;
        RECT 382.350 1029.675 382.630 1030.045 ;
        RECT 382.420 1027.325 382.560 1029.675 ;
        RECT 382.350 1026.955 382.630 1027.325 ;
        RECT 2076.990 32.795 2077.270 33.165 ;
        RECT 2124.830 32.795 2125.110 33.165 ;
        RECT 2077.060 30.445 2077.200 32.795 ;
        RECT 2124.900 30.445 2125.040 32.795 ;
        RECT 1103.170 30.075 1103.450 30.445 ;
        RECT 1296.830 30.075 1297.110 30.445 ;
        RECT 1973.030 30.075 1973.310 30.445 ;
        RECT 2076.990 30.075 2077.270 30.445 ;
        RECT 2124.830 30.075 2125.110 30.445 ;
        RECT 1007.960 29.765 1008.220 29.910 ;
        RECT 1055.340 29.765 1055.600 29.910 ;
        RECT 813.830 29.395 814.110 29.765 ;
        RECT 1007.950 29.395 1008.230 29.765 ;
        RECT 1055.330 29.395 1055.610 29.765 ;
        RECT 676.290 28.715 676.570 29.085 ;
        RECT 676.300 28.570 676.560 28.715 ;
        RECT 724.140 28.570 724.400 28.890 ;
        RECT 724.200 28.290 724.340 28.570 ;
        RECT 725.050 28.290 725.330 28.405 ;
        RECT 724.200 28.150 725.330 28.290 ;
        RECT 725.050 28.035 725.330 28.150 ;
        RECT 813.900 27.725 814.040 29.395 ;
        RECT 999.670 28.715 999.950 29.085 ;
        RECT 999.740 28.550 999.880 28.715 ;
        RECT 910.900 28.405 911.160 28.550 ;
        RECT 910.890 28.035 911.170 28.405 ;
        RECT 999.680 28.230 999.940 28.550 ;
        RECT 813.830 27.355 814.110 27.725 ;
        RECT 815.210 27.610 815.490 27.725 ;
        RECT 814.820 27.470 815.490 27.610 ;
        RECT 814.820 27.045 814.960 27.470 ;
        RECT 815.210 27.355 815.490 27.470 ;
        RECT 1103.240 27.045 1103.380 30.075 ;
        RECT 1296.900 28.405 1297.040 30.075 ;
        RECT 1369.510 28.715 1369.790 29.085 ;
        RECT 1414.130 28.970 1414.410 29.085 ;
        RECT 1415.050 28.970 1415.330 29.085 ;
        RECT 1414.130 28.830 1415.330 28.970 ;
        RECT 1414.130 28.715 1414.410 28.830 ;
        RECT 1415.050 28.715 1415.330 28.830 ;
        RECT 1654.250 28.970 1654.530 29.085 ;
        RECT 1654.250 28.830 1654.920 28.970 ;
        RECT 1654.250 28.715 1654.530 28.830 ;
        RECT 1296.830 28.035 1297.110 28.405 ;
        RECT 1369.580 27.725 1369.720 28.715 ;
        RECT 1654.780 28.405 1654.920 28.830 ;
        RECT 1876.430 28.715 1876.710 29.085 ;
        RECT 1654.710 28.035 1654.990 28.405 ;
        RECT 1752.230 28.290 1752.510 28.405 ;
        RECT 1753.150 28.290 1753.430 28.405 ;
        RECT 1752.230 28.150 1753.430 28.290 ;
        RECT 1752.230 28.035 1752.510 28.150 ;
        RECT 1753.150 28.035 1753.430 28.150 ;
        RECT 1876.500 27.725 1876.640 28.715 ;
        RECT 1973.100 28.405 1973.240 30.075 ;
        RECT 2409.120 29.765 2409.380 29.910 ;
        RECT 2456.040 29.765 2456.300 29.910 ;
        RECT 2342.410 29.395 2342.690 29.765 ;
        RECT 2409.110 29.395 2409.390 29.765 ;
        RECT 2456.030 29.395 2456.310 29.765 ;
        RECT 2190.610 28.715 2190.890 29.085 ;
        RECT 2214.530 28.715 2214.810 29.085 ;
        RECT 2235.230 28.970 2235.510 29.085 ;
        RECT 2235.230 28.830 2236.360 28.970 ;
        RECT 2235.230 28.715 2235.510 28.830 ;
        RECT 2190.620 28.570 2190.880 28.715 ;
        RECT 2214.540 28.570 2214.800 28.715 ;
        RECT 2236.220 28.405 2236.360 28.830 ;
        RECT 1973.030 28.035 1973.310 28.405 ;
        RECT 2236.150 28.035 2236.430 28.405 ;
        RECT 2342.480 27.725 2342.620 29.395 ;
        RECT 2573.330 28.970 2573.610 29.085 ;
        RECT 2574.250 28.970 2574.530 29.085 ;
        RECT 2573.330 28.830 2574.530 28.970 ;
        RECT 2573.330 28.715 2573.610 28.830 ;
        RECT 2574.250 28.715 2574.530 28.830 ;
        RECT 2632.210 28.715 2632.490 29.085 ;
        RECT 2632.280 27.725 2632.420 28.715 ;
        RECT 1369.510 27.355 1369.790 27.725 ;
        RECT 1876.430 27.355 1876.710 27.725 ;
        RECT 2342.410 27.355 2342.690 27.725 ;
        RECT 2632.210 27.355 2632.490 27.725 ;
        RECT 814.750 26.675 815.030 27.045 ;
        RECT 1103.170 26.675 1103.450 27.045 ;
        RECT 2678.670 19.875 2678.950 20.245 ;
        RECT 2678.740 2.400 2678.880 19.875 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
      LAYER via2 ;
        RECT 382.350 1029.720 382.630 1030.000 ;
        RECT 382.350 1027.000 382.630 1027.280 ;
        RECT 2076.990 32.840 2077.270 33.120 ;
        RECT 2124.830 32.840 2125.110 33.120 ;
        RECT 1103.170 30.120 1103.450 30.400 ;
        RECT 1296.830 30.120 1297.110 30.400 ;
        RECT 1973.030 30.120 1973.310 30.400 ;
        RECT 2076.990 30.120 2077.270 30.400 ;
        RECT 2124.830 30.120 2125.110 30.400 ;
        RECT 813.830 29.440 814.110 29.720 ;
        RECT 1007.950 29.440 1008.230 29.720 ;
        RECT 1055.330 29.440 1055.610 29.720 ;
        RECT 676.290 28.760 676.570 29.040 ;
        RECT 725.050 28.080 725.330 28.360 ;
        RECT 999.670 28.760 999.950 29.040 ;
        RECT 910.890 28.080 911.170 28.360 ;
        RECT 813.830 27.400 814.110 27.680 ;
        RECT 815.210 27.400 815.490 27.680 ;
        RECT 1369.510 28.760 1369.790 29.040 ;
        RECT 1414.130 28.760 1414.410 29.040 ;
        RECT 1415.050 28.760 1415.330 29.040 ;
        RECT 1654.250 28.760 1654.530 29.040 ;
        RECT 1296.830 28.080 1297.110 28.360 ;
        RECT 1876.430 28.760 1876.710 29.040 ;
        RECT 1654.710 28.080 1654.990 28.360 ;
        RECT 1752.230 28.080 1752.510 28.360 ;
        RECT 1753.150 28.080 1753.430 28.360 ;
        RECT 2342.410 29.440 2342.690 29.720 ;
        RECT 2409.110 29.440 2409.390 29.720 ;
        RECT 2456.030 29.440 2456.310 29.720 ;
        RECT 2190.610 28.760 2190.890 29.040 ;
        RECT 2214.530 28.760 2214.810 29.040 ;
        RECT 2235.230 28.760 2235.510 29.040 ;
        RECT 1973.030 28.080 1973.310 28.360 ;
        RECT 2236.150 28.080 2236.430 28.360 ;
        RECT 2573.330 28.760 2573.610 29.040 ;
        RECT 2574.250 28.760 2574.530 29.040 ;
        RECT 2632.210 28.760 2632.490 29.040 ;
        RECT 1369.510 27.400 1369.790 27.680 ;
        RECT 1876.430 27.400 1876.710 27.680 ;
        RECT 2342.410 27.400 2342.690 27.680 ;
        RECT 2632.210 27.400 2632.490 27.680 ;
        RECT 814.750 26.720 815.030 27.000 ;
        RECT 1103.170 26.720 1103.450 27.000 ;
        RECT 2678.670 19.920 2678.950 20.200 ;
      LAYER met3 ;
        RECT 385.750 2759.930 386.130 2759.940 ;
        RECT 410.000 2759.930 414.000 2760.080 ;
        RECT 385.750 2759.630 414.000 2759.930 ;
        RECT 385.750 2759.620 386.130 2759.630 ;
        RECT 410.000 2759.480 414.000 2759.630 ;
        RECT 382.325 1030.010 382.655 1030.025 ;
        RECT 385.750 1030.010 386.130 1030.020 ;
        RECT 382.325 1029.710 386.130 1030.010 ;
        RECT 382.325 1029.695 382.655 1029.710 ;
        RECT 385.750 1029.700 386.130 1029.710 ;
        RECT 382.325 1027.290 382.655 1027.305 ;
        RECT 385.750 1027.290 386.130 1027.300 ;
        RECT 382.325 1026.990 386.130 1027.290 ;
        RECT 382.325 1026.975 382.655 1026.990 ;
        RECT 385.750 1026.980 386.130 1026.990 ;
        RECT 2076.965 33.130 2077.295 33.145 ;
        RECT 2124.805 33.130 2125.135 33.145 ;
        RECT 2076.965 32.830 2125.135 33.130 ;
        RECT 2076.965 32.815 2077.295 32.830 ;
        RECT 2124.805 32.815 2125.135 32.830 ;
        RECT 1103.145 30.410 1103.475 30.425 ;
        RECT 1110.710 30.410 1111.090 30.420 ;
        RECT 1103.145 30.110 1111.090 30.410 ;
        RECT 1103.145 30.095 1103.475 30.110 ;
        RECT 1110.710 30.100 1111.090 30.110 ;
        RECT 1152.110 30.410 1152.490 30.420 ;
        RECT 1199.950 30.410 1200.330 30.420 ;
        RECT 1152.110 30.110 1200.330 30.410 ;
        RECT 1152.110 30.100 1152.490 30.110 ;
        RECT 1199.950 30.100 1200.330 30.110 ;
        RECT 1248.710 30.410 1249.090 30.420 ;
        RECT 1296.805 30.410 1297.135 30.425 ;
        RECT 1248.710 30.110 1297.135 30.410 ;
        RECT 1248.710 30.100 1249.090 30.110 ;
        RECT 1296.805 30.095 1297.135 30.110 ;
        RECT 1441.910 30.410 1442.290 30.420 ;
        RECT 1489.750 30.410 1490.130 30.420 ;
        RECT 1441.910 30.110 1490.130 30.410 ;
        RECT 1441.910 30.100 1442.290 30.110 ;
        RECT 1489.750 30.100 1490.130 30.110 ;
        RECT 1924.910 30.410 1925.290 30.420 ;
        RECT 1973.005 30.410 1973.335 30.425 ;
        RECT 1924.910 30.110 1973.335 30.410 ;
        RECT 1924.910 30.100 1925.290 30.110 ;
        RECT 1973.005 30.095 1973.335 30.110 ;
        RECT 2028.870 30.410 2029.250 30.420 ;
        RECT 2076.965 30.410 2077.295 30.425 ;
        RECT 2028.870 30.110 2077.295 30.410 ;
        RECT 2028.870 30.100 2029.250 30.110 ;
        RECT 2076.965 30.095 2077.295 30.110 ;
        RECT 2124.805 30.410 2125.135 30.425 ;
        RECT 2124.805 30.110 2166.290 30.410 ;
        RECT 2124.805 30.095 2125.135 30.110 ;
        RECT 765.710 29.730 766.090 29.740 ;
        RECT 813.805 29.730 814.135 29.745 ;
        RECT 1007.925 29.730 1008.255 29.745 ;
        RECT 1055.305 29.740 1055.635 29.745 ;
        RECT 1055.305 29.730 1055.890 29.740 ;
        RECT 2165.990 29.730 2166.290 30.110 ;
        RECT 2342.385 29.730 2342.715 29.745 ;
        RECT 2409.085 29.730 2409.415 29.745 ;
        RECT 765.710 29.430 814.135 29.730 ;
        RECT 765.710 29.420 766.090 29.430 ;
        RECT 813.805 29.415 814.135 29.430 ;
        RECT 1007.710 29.415 1008.255 29.730 ;
        RECT 1055.100 29.430 1055.890 29.730 ;
        RECT 1055.305 29.420 1055.890 29.430 ;
        RECT 1393.190 29.430 1400.850 29.730 ;
        RECT 2165.990 29.430 2167.210 29.730 ;
        RECT 1055.305 29.415 1055.635 29.420 ;
        RECT 385.750 29.050 386.130 29.060 ;
        RECT 676.265 29.050 676.595 29.065 ;
        RECT 385.750 28.750 676.595 29.050 ;
        RECT 385.750 28.740 386.130 28.750 ;
        RECT 676.265 28.735 676.595 28.750 ;
        RECT 999.645 29.050 999.975 29.065 ;
        RECT 1007.710 29.050 1008.010 29.415 ;
        RECT 999.645 28.750 1008.010 29.050 ;
        RECT 1199.950 29.050 1200.330 29.060 ;
        RECT 1248.710 29.050 1249.090 29.060 ;
        RECT 1199.950 28.750 1249.090 29.050 ;
        RECT 999.645 28.735 999.975 28.750 ;
        RECT 1199.950 28.740 1200.330 28.750 ;
        RECT 1248.710 28.740 1249.090 28.750 ;
        RECT 1304.830 29.050 1305.210 29.060 ;
        RECT 1345.310 29.050 1345.690 29.060 ;
        RECT 1304.830 28.750 1345.690 29.050 ;
        RECT 1304.830 28.740 1305.210 28.750 ;
        RECT 1345.310 28.740 1345.690 28.750 ;
        RECT 1369.485 29.050 1369.815 29.065 ;
        RECT 1393.190 29.050 1393.490 29.430 ;
        RECT 1369.485 28.750 1393.490 29.050 ;
        RECT 1400.550 29.050 1400.850 29.430 ;
        RECT 1414.105 29.050 1414.435 29.065 ;
        RECT 1400.550 28.750 1414.435 29.050 ;
        RECT 1369.485 28.735 1369.815 28.750 ;
        RECT 1414.105 28.735 1414.435 28.750 ;
        RECT 1415.025 29.050 1415.355 29.065 ;
        RECT 1441.910 29.050 1442.290 29.060 ;
        RECT 1415.025 28.750 1442.290 29.050 ;
        RECT 1415.025 28.735 1415.355 28.750 ;
        RECT 1441.910 28.740 1442.290 28.750 ;
        RECT 1489.750 29.050 1490.130 29.060 ;
        RECT 1538.510 29.050 1538.890 29.060 ;
        RECT 1489.750 28.750 1538.890 29.050 ;
        RECT 1489.750 28.740 1490.130 28.750 ;
        RECT 1538.510 28.740 1538.890 28.750 ;
        RECT 1586.350 29.050 1586.730 29.060 ;
        RECT 1654.225 29.050 1654.555 29.065 ;
        RECT 1800.710 29.050 1801.090 29.060 ;
        RECT 1586.350 28.750 1654.555 29.050 ;
        RECT 1586.350 28.740 1586.730 28.750 ;
        RECT 1654.225 28.735 1654.555 28.750 ;
        RECT 1707.830 28.750 1732.050 29.050 ;
        RECT 725.025 28.370 725.355 28.385 ;
        RECT 765.710 28.370 766.090 28.380 ;
        RECT 910.865 28.370 911.195 28.385 ;
        RECT 725.025 28.070 766.090 28.370 ;
        RECT 725.025 28.055 725.355 28.070 ;
        RECT 765.710 28.060 766.090 28.070 ;
        RECT 862.350 28.070 911.195 28.370 ;
        RECT 813.805 27.690 814.135 27.705 ;
        RECT 815.185 27.690 815.515 27.705 ;
        RECT 862.350 27.690 862.650 28.070 ;
        RECT 910.865 28.055 911.195 28.070 ;
        RECT 1296.805 28.370 1297.135 28.385 ;
        RECT 1303.910 28.370 1304.290 28.380 ;
        RECT 1296.805 28.070 1304.290 28.370 ;
        RECT 1296.805 28.055 1297.135 28.070 ;
        RECT 1303.910 28.060 1304.290 28.070 ;
        RECT 1654.685 28.370 1655.015 28.385 ;
        RECT 1707.830 28.370 1708.130 28.750 ;
        RECT 1654.685 28.070 1708.130 28.370 ;
        RECT 1731.750 28.370 1732.050 28.750 ;
        RECT 1786.950 28.750 1801.090 29.050 ;
        RECT 1752.205 28.370 1752.535 28.385 ;
        RECT 1731.750 28.070 1752.535 28.370 ;
        RECT 1654.685 28.055 1655.015 28.070 ;
        RECT 1752.205 28.055 1752.535 28.070 ;
        RECT 1753.125 28.370 1753.455 28.385 ;
        RECT 1786.950 28.370 1787.250 28.750 ;
        RECT 1800.710 28.740 1801.090 28.750 ;
        RECT 1801.630 29.050 1802.010 29.060 ;
        RECT 1828.310 29.050 1828.690 29.060 ;
        RECT 1801.630 28.750 1828.690 29.050 ;
        RECT 1801.630 28.740 1802.010 28.750 ;
        RECT 1828.310 28.740 1828.690 28.750 ;
        RECT 1876.405 29.050 1876.735 29.065 ;
        RECT 1924.910 29.050 1925.290 29.060 ;
        RECT 1876.405 28.750 1925.290 29.050 ;
        RECT 2166.910 29.050 2167.210 29.430 ;
        RECT 2342.385 29.430 2409.415 29.730 ;
        RECT 2342.385 29.415 2342.715 29.430 ;
        RECT 2409.085 29.415 2409.415 29.430 ;
        RECT 2456.005 29.730 2456.335 29.745 ;
        RECT 2456.005 29.430 2512.210 29.730 ;
        RECT 2456.005 29.415 2456.335 29.430 ;
        RECT 2190.585 29.050 2190.915 29.065 ;
        RECT 2166.910 28.750 2190.915 29.050 ;
        RECT 1876.405 28.735 1876.735 28.750 ;
        RECT 1924.910 28.740 1925.290 28.750 ;
        RECT 2190.585 28.735 2190.915 28.750 ;
        RECT 2214.505 29.050 2214.835 29.065 ;
        RECT 2235.205 29.050 2235.535 29.065 ;
        RECT 2283.710 29.050 2284.090 29.060 ;
        RECT 2214.505 28.750 2235.535 29.050 ;
        RECT 2214.505 28.735 2214.835 28.750 ;
        RECT 2235.205 28.735 2235.535 28.750 ;
        RECT 2269.950 28.750 2284.090 29.050 ;
        RECT 1753.125 28.070 1787.250 28.370 ;
        RECT 1973.005 28.370 1973.335 28.385 ;
        RECT 2028.870 28.370 2029.250 28.380 ;
        RECT 1973.005 28.070 2029.250 28.370 ;
        RECT 1753.125 28.055 1753.455 28.070 ;
        RECT 1973.005 28.055 1973.335 28.070 ;
        RECT 2028.870 28.060 2029.250 28.070 ;
        RECT 2236.125 28.370 2236.455 28.385 ;
        RECT 2269.950 28.370 2270.250 28.750 ;
        RECT 2283.710 28.740 2284.090 28.750 ;
        RECT 2284.630 29.050 2285.010 29.060 ;
        RECT 2511.910 29.050 2512.210 29.430 ;
        RECT 2573.305 29.050 2573.635 29.065 ;
        RECT 2284.630 28.750 2319.010 29.050 ;
        RECT 2511.910 28.750 2573.635 29.050 ;
        RECT 2284.630 28.740 2285.010 28.750 ;
        RECT 2236.125 28.070 2270.250 28.370 ;
        RECT 2236.125 28.055 2236.455 28.070 ;
        RECT 813.805 27.390 814.810 27.690 ;
        RECT 813.805 27.375 814.135 27.390 ;
        RECT 814.510 27.025 814.810 27.390 ;
        RECT 815.185 27.390 862.650 27.690 ;
        RECT 1110.710 27.690 1111.090 27.700 ;
        RECT 1152.110 27.690 1152.490 27.700 ;
        RECT 1110.710 27.390 1152.490 27.690 ;
        RECT 815.185 27.375 815.515 27.390 ;
        RECT 1110.710 27.380 1111.090 27.390 ;
        RECT 1152.110 27.380 1152.490 27.390 ;
        RECT 1345.310 27.690 1345.690 27.700 ;
        RECT 1369.485 27.690 1369.815 27.705 ;
        RECT 1345.310 27.390 1369.815 27.690 ;
        RECT 1345.310 27.380 1345.690 27.390 ;
        RECT 1369.485 27.375 1369.815 27.390 ;
        RECT 1538.510 27.690 1538.890 27.700 ;
        RECT 1586.350 27.690 1586.730 27.700 ;
        RECT 1538.510 27.390 1586.730 27.690 ;
        RECT 1538.510 27.380 1538.890 27.390 ;
        RECT 1586.350 27.380 1586.730 27.390 ;
        RECT 1828.310 27.690 1828.690 27.700 ;
        RECT 1876.405 27.690 1876.735 27.705 ;
        RECT 1828.310 27.390 1876.735 27.690 ;
        RECT 2318.710 27.690 2319.010 28.750 ;
        RECT 2573.305 28.735 2573.635 28.750 ;
        RECT 2574.225 29.050 2574.555 29.065 ;
        RECT 2632.185 29.050 2632.515 29.065 ;
        RECT 2677.470 29.050 2677.850 29.060 ;
        RECT 2574.225 28.750 2608.810 29.050 ;
        RECT 2574.225 28.735 2574.555 28.750 ;
        RECT 2342.385 27.690 2342.715 27.705 ;
        RECT 2318.710 27.390 2342.715 27.690 ;
        RECT 2608.510 27.690 2608.810 28.750 ;
        RECT 2632.185 28.750 2677.850 29.050 ;
        RECT 2632.185 28.735 2632.515 28.750 ;
        RECT 2677.470 28.740 2677.850 28.750 ;
        RECT 2632.185 27.690 2632.515 27.705 ;
        RECT 2608.510 27.390 2632.515 27.690 ;
        RECT 1828.310 27.380 1828.690 27.390 ;
        RECT 1876.405 27.375 1876.735 27.390 ;
        RECT 2342.385 27.375 2342.715 27.390 ;
        RECT 2632.185 27.375 2632.515 27.390 ;
        RECT 814.510 26.710 815.055 27.025 ;
        RECT 814.725 26.695 815.055 26.710 ;
        RECT 1055.510 27.010 1055.890 27.020 ;
        RECT 1103.145 27.010 1103.475 27.025 ;
        RECT 1055.510 26.710 1103.475 27.010 ;
        RECT 1055.510 26.700 1055.890 26.710 ;
        RECT 1103.145 26.695 1103.475 26.710 ;
        RECT 2677.470 20.210 2677.850 20.220 ;
        RECT 2678.645 20.210 2678.975 20.225 ;
        RECT 2677.470 19.910 2678.975 20.210 ;
        RECT 2677.470 19.900 2677.850 19.910 ;
        RECT 2678.645 19.895 2678.975 19.910 ;
      LAYER via3 ;
        RECT 385.780 2759.620 386.100 2759.940 ;
        RECT 385.780 1029.700 386.100 1030.020 ;
        RECT 385.780 1026.980 386.100 1027.300 ;
        RECT 1110.740 30.100 1111.060 30.420 ;
        RECT 1152.140 30.100 1152.460 30.420 ;
        RECT 1199.980 30.100 1200.300 30.420 ;
        RECT 1248.740 30.100 1249.060 30.420 ;
        RECT 1441.940 30.100 1442.260 30.420 ;
        RECT 1489.780 30.100 1490.100 30.420 ;
        RECT 1924.940 30.100 1925.260 30.420 ;
        RECT 2028.900 30.100 2029.220 30.420 ;
        RECT 765.740 29.420 766.060 29.740 ;
        RECT 1055.540 29.420 1055.860 29.740 ;
        RECT 385.780 28.740 386.100 29.060 ;
        RECT 1199.980 28.740 1200.300 29.060 ;
        RECT 1248.740 28.740 1249.060 29.060 ;
        RECT 1304.860 28.740 1305.180 29.060 ;
        RECT 1345.340 28.740 1345.660 29.060 ;
        RECT 1441.940 28.740 1442.260 29.060 ;
        RECT 1489.780 28.740 1490.100 29.060 ;
        RECT 1538.540 28.740 1538.860 29.060 ;
        RECT 1586.380 28.740 1586.700 29.060 ;
        RECT 765.740 28.060 766.060 28.380 ;
        RECT 1303.940 28.060 1304.260 28.380 ;
        RECT 1800.740 28.740 1801.060 29.060 ;
        RECT 1801.660 28.740 1801.980 29.060 ;
        RECT 1828.340 28.740 1828.660 29.060 ;
        RECT 1924.940 28.740 1925.260 29.060 ;
        RECT 2028.900 28.060 2029.220 28.380 ;
        RECT 2283.740 28.740 2284.060 29.060 ;
        RECT 2284.660 28.740 2284.980 29.060 ;
        RECT 1110.740 27.380 1111.060 27.700 ;
        RECT 1152.140 27.380 1152.460 27.700 ;
        RECT 1345.340 27.380 1345.660 27.700 ;
        RECT 1538.540 27.380 1538.860 27.700 ;
        RECT 1586.380 27.380 1586.700 27.700 ;
        RECT 1828.340 27.380 1828.660 27.700 ;
        RECT 2677.500 28.740 2677.820 29.060 ;
        RECT 1055.540 26.700 1055.860 27.020 ;
        RECT 2677.500 19.900 2677.820 20.220 ;
      LAYER met4 ;
        RECT 385.775 2759.615 386.105 2759.945 ;
        RECT 385.790 1030.025 386.090 2759.615 ;
        RECT 385.775 1029.695 386.105 1030.025 ;
        RECT 385.775 1026.975 386.105 1027.305 ;
        RECT 385.790 29.065 386.090 1026.975 ;
        RECT 1110.735 30.095 1111.065 30.425 ;
        RECT 1152.135 30.095 1152.465 30.425 ;
        RECT 1199.975 30.095 1200.305 30.425 ;
        RECT 1248.735 30.095 1249.065 30.425 ;
        RECT 1441.935 30.095 1442.265 30.425 ;
        RECT 1489.775 30.095 1490.105 30.425 ;
        RECT 1924.935 30.095 1925.265 30.425 ;
        RECT 2028.895 30.095 2029.225 30.425 ;
        RECT 765.735 29.415 766.065 29.745 ;
        RECT 1055.535 29.415 1055.865 29.745 ;
        RECT 385.775 28.735 386.105 29.065 ;
        RECT 765.750 28.385 766.050 29.415 ;
        RECT 765.735 28.055 766.065 28.385 ;
        RECT 1055.550 27.025 1055.850 29.415 ;
        RECT 1110.750 27.705 1111.050 30.095 ;
        RECT 1152.150 27.705 1152.450 30.095 ;
        RECT 1199.990 29.065 1200.290 30.095 ;
        RECT 1248.750 29.065 1249.050 30.095 ;
        RECT 1441.950 29.065 1442.250 30.095 ;
        RECT 1489.790 29.065 1490.090 30.095 ;
        RECT 1924.950 29.065 1925.250 30.095 ;
        RECT 1199.975 28.735 1200.305 29.065 ;
        RECT 1248.735 28.735 1249.065 29.065 ;
        RECT 1304.855 29.050 1305.185 29.065 ;
        RECT 1303.950 28.750 1305.185 29.050 ;
        RECT 1303.950 28.385 1304.250 28.750 ;
        RECT 1304.855 28.735 1305.185 28.750 ;
        RECT 1345.335 28.735 1345.665 29.065 ;
        RECT 1441.935 28.735 1442.265 29.065 ;
        RECT 1489.775 28.735 1490.105 29.065 ;
        RECT 1538.535 28.735 1538.865 29.065 ;
        RECT 1586.375 28.735 1586.705 29.065 ;
        RECT 1800.735 29.050 1801.065 29.065 ;
        RECT 1801.655 29.050 1801.985 29.065 ;
        RECT 1800.735 28.750 1801.985 29.050 ;
        RECT 1800.735 28.735 1801.065 28.750 ;
        RECT 1801.655 28.735 1801.985 28.750 ;
        RECT 1828.335 28.735 1828.665 29.065 ;
        RECT 1924.935 28.735 1925.265 29.065 ;
        RECT 1303.935 28.055 1304.265 28.385 ;
        RECT 1345.350 27.705 1345.650 28.735 ;
        RECT 1538.550 27.705 1538.850 28.735 ;
        RECT 1586.390 27.705 1586.690 28.735 ;
        RECT 1828.350 27.705 1828.650 28.735 ;
        RECT 2028.910 28.385 2029.210 30.095 ;
        RECT 2283.735 29.050 2284.065 29.065 ;
        RECT 2284.655 29.050 2284.985 29.065 ;
        RECT 2283.735 28.750 2284.985 29.050 ;
        RECT 2283.735 28.735 2284.065 28.750 ;
        RECT 2284.655 28.735 2284.985 28.750 ;
        RECT 2677.495 28.735 2677.825 29.065 ;
        RECT 2028.895 28.055 2029.225 28.385 ;
        RECT 1110.735 27.375 1111.065 27.705 ;
        RECT 1152.135 27.375 1152.465 27.705 ;
        RECT 1345.335 27.375 1345.665 27.705 ;
        RECT 1538.535 27.375 1538.865 27.705 ;
        RECT 1586.375 27.375 1586.705 27.705 ;
        RECT 1828.335 27.375 1828.665 27.705 ;
        RECT 1055.535 26.695 1055.865 27.025 ;
        RECT 2677.510 20.225 2677.810 28.735 ;
        RECT 2677.495 19.895 2677.825 20.225 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 390.150 217.160 390.470 217.220 ;
        RECT 2691.070 217.160 2691.390 217.220 ;
        RECT 390.150 217.020 2691.390 217.160 ;
        RECT 390.150 216.960 390.470 217.020 ;
        RECT 2691.070 216.960 2691.390 217.020 ;
      LAYER via ;
        RECT 390.180 216.960 390.440 217.220 ;
        RECT 2691.100 216.960 2691.360 217.220 ;
      LAYER met2 ;
        RECT 390.170 805.275 390.450 805.645 ;
        RECT 390.240 217.250 390.380 805.275 ;
        RECT 390.180 216.930 390.440 217.250 ;
        RECT 2691.100 216.930 2691.360 217.250 ;
        RECT 2691.160 17.410 2691.300 216.930 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 390.170 805.320 390.450 805.600 ;
      LAYER met3 ;
        RECT 390.145 805.610 390.475 805.625 ;
        RECT 410.000 805.610 414.000 805.760 ;
        RECT 390.145 805.310 414.000 805.610 ;
        RECT 390.145 805.295 390.475 805.310 ;
        RECT 410.000 805.160 414.000 805.310 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1075.165 3002.625 1075.335 3006.535 ;
      LAYER mcon ;
        RECT 1075.165 3006.365 1075.335 3006.535 ;
      LAYER met1 ;
        RECT 1075.090 3006.520 1075.410 3006.580 ;
        RECT 1074.895 3006.380 1075.410 3006.520 ;
        RECT 1075.090 3006.320 1075.410 3006.380 ;
        RECT 1075.105 3002.780 1075.395 3002.825 ;
        RECT 2590.790 3002.780 2591.110 3002.840 ;
        RECT 1075.105 3002.640 2591.110 3002.780 ;
        RECT 1075.105 3002.595 1075.395 3002.640 ;
        RECT 2590.790 3002.580 2591.110 3002.640 ;
        RECT 2590.790 17.580 2591.110 17.640 ;
        RECT 2714.530 17.580 2714.850 17.640 ;
        RECT 2590.790 17.440 2714.850 17.580 ;
        RECT 2590.790 17.380 2591.110 17.440 ;
        RECT 2714.530 17.380 2714.850 17.440 ;
      LAYER via ;
        RECT 1075.120 3006.320 1075.380 3006.580 ;
        RECT 2590.820 3002.580 2591.080 3002.840 ;
        RECT 2590.820 17.380 2591.080 17.640 ;
        RECT 2714.560 17.380 2714.820 17.640 ;
      LAYER met2 ;
        RECT 1074.330 3006.690 1074.610 3010.000 ;
        RECT 1074.330 3006.610 1075.320 3006.690 ;
        RECT 1074.330 3006.550 1075.380 3006.610 ;
        RECT 1074.330 3006.000 1074.610 3006.550 ;
        RECT 1075.120 3006.290 1075.380 3006.550 ;
        RECT 2590.820 3002.550 2591.080 3002.870 ;
        RECT 2590.880 17.670 2591.020 3002.550 ;
        RECT 2590.820 17.350 2591.080 17.670 ;
        RECT 2714.560 17.350 2714.820 17.670 ;
        RECT 2714.620 2.400 2714.760 17.350 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 3009.920 1545.530 3009.980 ;
        RECT 2714.990 3009.920 2715.310 3009.980 ;
        RECT 1545.210 3009.780 2715.310 3009.920 ;
        RECT 1545.210 3009.720 1545.530 3009.780 ;
        RECT 2714.990 3009.720 2715.310 3009.780 ;
        RECT 2714.990 16.560 2715.310 16.620 ;
        RECT 2732.470 16.560 2732.790 16.620 ;
        RECT 2714.990 16.420 2732.790 16.560 ;
        RECT 2714.990 16.360 2715.310 16.420 ;
        RECT 2732.470 16.360 2732.790 16.420 ;
      LAYER via ;
        RECT 1545.240 3009.720 1545.500 3009.980 ;
        RECT 2715.020 3009.720 2715.280 3009.980 ;
        RECT 2715.020 16.360 2715.280 16.620 ;
        RECT 2732.500 16.360 2732.760 16.620 ;
      LAYER met2 ;
        RECT 1543.530 3009.410 1543.810 3010.000 ;
        RECT 1545.240 3009.690 1545.500 3010.010 ;
        RECT 2715.020 3009.690 2715.280 3010.010 ;
        RECT 1545.300 3009.410 1545.440 3009.690 ;
        RECT 1543.530 3009.270 1545.440 3009.410 ;
        RECT 1543.530 3006.000 1543.810 3009.270 ;
        RECT 2715.080 16.650 2715.220 3009.690 ;
        RECT 2715.020 16.330 2715.280 16.650 ;
        RECT 2732.500 16.330 2732.760 16.650 ;
        RECT 2732.560 2.400 2732.700 16.330 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1228.320 2520.730 1228.380 ;
        RECT 2735.690 1228.320 2736.010 1228.380 ;
        RECT 2520.410 1228.180 2736.010 1228.320 ;
        RECT 2520.410 1228.120 2520.730 1228.180 ;
        RECT 2735.690 1228.120 2736.010 1228.180 ;
        RECT 2735.690 90.000 2736.010 90.060 ;
        RECT 2746.270 90.000 2746.590 90.060 ;
        RECT 2735.690 89.860 2746.590 90.000 ;
        RECT 2735.690 89.800 2736.010 89.860 ;
        RECT 2746.270 89.800 2746.590 89.860 ;
      LAYER via ;
        RECT 2520.440 1228.120 2520.700 1228.380 ;
        RECT 2735.720 1228.120 2735.980 1228.380 ;
        RECT 2735.720 89.800 2735.980 90.060 ;
        RECT 2746.300 89.800 2746.560 90.060 ;
      LAYER met2 ;
        RECT 2520.430 1233.675 2520.710 1234.045 ;
        RECT 2520.500 1228.410 2520.640 1233.675 ;
        RECT 2520.440 1228.090 2520.700 1228.410 ;
        RECT 2735.720 1228.090 2735.980 1228.410 ;
        RECT 2735.780 90.090 2735.920 1228.090 ;
        RECT 2735.720 89.770 2735.980 90.090 ;
        RECT 2746.300 89.770 2746.560 90.090 ;
        RECT 2746.360 17.410 2746.500 89.770 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1233.720 2520.710 1234.000 ;
      LAYER met3 ;
        RECT 2506.000 1234.010 2510.000 1234.160 ;
        RECT 2520.405 1234.010 2520.735 1234.025 ;
        RECT 2506.000 1233.710 2520.735 1234.010 ;
        RECT 2506.000 1233.560 2510.000 1233.710 ;
        RECT 2520.405 1233.695 2520.735 1233.710 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.050 362.340 420.370 362.400 ;
        RECT 2766.970 362.340 2767.290 362.400 ;
        RECT 420.050 362.200 2767.290 362.340 ;
        RECT 420.050 362.140 420.370 362.200 ;
        RECT 2766.970 362.140 2767.290 362.200 ;
      LAYER via ;
        RECT 420.080 362.140 420.340 362.400 ;
        RECT 2767.000 362.140 2767.260 362.400 ;
      LAYER met2 ;
        RECT 420.070 512.195 420.350 512.565 ;
        RECT 420.140 362.430 420.280 512.195 ;
        RECT 420.080 362.110 420.340 362.430 ;
        RECT 2767.000 362.110 2767.260 362.430 ;
        RECT 2767.060 17.410 2767.200 362.110 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
      LAYER via2 ;
        RECT 420.070 512.240 420.350 512.520 ;
      LAYER met3 ;
        RECT 410.000 1426.680 414.000 1427.280 ;
        RECT 412.470 1424.420 412.770 1426.680 ;
        RECT 412.430 1424.100 412.810 1424.420 ;
        RECT 414.270 512.530 414.650 512.540 ;
        RECT 420.045 512.530 420.375 512.545 ;
        RECT 414.270 512.230 420.375 512.530 ;
        RECT 414.270 512.220 414.650 512.230 ;
        RECT 420.045 512.215 420.375 512.230 ;
      LAYER via3 ;
        RECT 412.460 1424.100 412.780 1424.420 ;
        RECT 414.300 512.220 414.620 512.540 ;
      LAYER met4 ;
        RECT 412.455 1424.095 412.785 1424.425 ;
        RECT 412.470 1423.050 412.770 1424.095 ;
        RECT 412.470 1422.750 414.610 1423.050 ;
        RECT 414.310 512.545 414.610 1422.750 ;
        RECT 414.295 512.215 414.625 512.545 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 330.810 3032.700 331.130 3032.760 ;
        RECT 950.890 3032.700 951.210 3032.760 ;
        RECT 330.810 3032.560 951.210 3032.700 ;
        RECT 330.810 3032.500 331.130 3032.560 ;
        RECT 950.890 3032.500 951.210 3032.560 ;
        RECT 330.810 494.940 331.130 495.000 ;
        RECT 834.970 494.940 835.290 495.000 ;
        RECT 330.810 494.800 835.290 494.940 ;
        RECT 330.810 494.740 331.130 494.800 ;
        RECT 834.970 494.740 835.290 494.800 ;
        RECT 834.970 20.300 835.290 20.360 ;
        RECT 840.950 20.300 841.270 20.360 ;
        RECT 834.970 20.160 841.270 20.300 ;
        RECT 834.970 20.100 835.290 20.160 ;
        RECT 840.950 20.100 841.270 20.160 ;
      LAYER via ;
        RECT 330.840 3032.500 331.100 3032.760 ;
        RECT 950.920 3032.500 951.180 3032.760 ;
        RECT 330.840 494.740 331.100 495.000 ;
        RECT 835.000 494.740 835.260 495.000 ;
        RECT 835.000 20.100 835.260 20.360 ;
        RECT 840.980 20.100 841.240 20.360 ;
      LAYER met2 ;
        RECT 330.840 3032.470 331.100 3032.790 ;
        RECT 950.920 3032.470 951.180 3032.790 ;
        RECT 330.900 495.030 331.040 3032.470 ;
        RECT 950.980 3010.000 951.120 3032.470 ;
        RECT 950.980 3009.340 951.330 3010.000 ;
        RECT 951.050 3006.000 951.330 3009.340 ;
        RECT 330.840 494.710 331.100 495.030 ;
        RECT 835.000 494.710 835.260 495.030 ;
        RECT 835.060 20.390 835.200 494.710 ;
        RECT 835.000 20.070 835.260 20.390 ;
        RECT 840.980 20.070 841.240 20.390 ;
        RECT 841.040 2.400 841.180 20.070 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1828.645 3002.965 1828.815 3006.535 ;
      LAYER mcon ;
        RECT 1828.645 3006.365 1828.815 3006.535 ;
      LAYER met1 ;
        RECT 1828.570 3006.520 1828.890 3006.580 ;
        RECT 1828.375 3006.380 1828.890 3006.520 ;
        RECT 1828.570 3006.320 1828.890 3006.380 ;
        RECT 1828.585 3003.120 1828.875 3003.165 ;
        RECT 2780.770 3003.120 2781.090 3003.180 ;
        RECT 1828.585 3002.980 2781.090 3003.120 ;
        RECT 1828.585 3002.935 1828.875 3002.980 ;
        RECT 2780.770 3002.920 2781.090 3002.980 ;
      LAYER via ;
        RECT 1828.600 3006.320 1828.860 3006.580 ;
        RECT 2780.800 3002.920 2781.060 3003.180 ;
      LAYER met2 ;
        RECT 1827.810 3006.690 1828.090 3010.000 ;
        RECT 1827.810 3006.610 1828.800 3006.690 ;
        RECT 1827.810 3006.550 1828.860 3006.610 ;
        RECT 1827.810 3006.000 1828.090 3006.550 ;
        RECT 1828.600 3006.290 1828.860 3006.550 ;
        RECT 2780.800 3002.890 2781.060 3003.210 ;
        RECT 2780.860 17.410 2781.000 3002.890 ;
        RECT 2780.860 17.270 2786.060 17.410 ;
        RECT 2785.920 2.400 2786.060 17.270 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 343.690 952.580 344.010 952.640 ;
        RECT 393.370 952.580 393.690 952.640 ;
        RECT 343.690 952.440 393.690 952.580 ;
        RECT 343.690 952.380 344.010 952.440 ;
        RECT 393.370 952.380 393.690 952.440 ;
        RECT 343.690 72.320 344.010 72.380 ;
        RECT 2801.470 72.320 2801.790 72.380 ;
        RECT 343.690 72.180 2801.790 72.320 ;
        RECT 343.690 72.120 344.010 72.180 ;
        RECT 2801.470 72.120 2801.790 72.180 ;
      LAYER via ;
        RECT 343.720 952.380 343.980 952.640 ;
        RECT 393.400 952.380 393.660 952.640 ;
        RECT 343.720 72.120 343.980 72.380 ;
        RECT 2801.500 72.120 2801.760 72.380 ;
      LAYER met2 ;
        RECT 343.720 952.350 343.980 952.670 ;
        RECT 393.400 952.525 393.660 952.670 ;
        RECT 343.780 72.410 343.920 952.350 ;
        RECT 393.390 952.155 393.670 952.525 ;
        RECT 343.720 72.090 343.980 72.410 ;
        RECT 2801.500 72.090 2801.760 72.410 ;
        RECT 2801.560 17.410 2801.700 72.090 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 393.390 952.200 393.670 952.480 ;
      LAYER met3 ;
        RECT 393.365 952.490 393.695 952.505 ;
        RECT 410.000 952.490 414.000 952.640 ;
        RECT 393.365 952.190 414.000 952.490 ;
        RECT 393.365 952.175 393.695 952.190 ;
        RECT 410.000 952.040 414.000 952.190 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2518.570 759.120 2518.890 759.180 ;
        RECT 2763.750 759.120 2764.070 759.180 ;
        RECT 2518.570 758.980 2764.070 759.120 ;
        RECT 2518.570 758.920 2518.890 758.980 ;
        RECT 2763.750 758.920 2764.070 758.980 ;
        RECT 2763.750 37.980 2764.070 38.040 ;
        RECT 2821.710 37.980 2822.030 38.040 ;
        RECT 2763.750 37.840 2822.030 37.980 ;
        RECT 2763.750 37.780 2764.070 37.840 ;
        RECT 2821.710 37.780 2822.030 37.840 ;
      LAYER via ;
        RECT 2518.600 758.920 2518.860 759.180 ;
        RECT 2763.780 758.920 2764.040 759.180 ;
        RECT 2763.780 37.780 2764.040 38.040 ;
        RECT 2821.740 37.780 2822.000 38.040 ;
      LAYER met2 ;
        RECT 2518.590 759.035 2518.870 759.405 ;
        RECT 2518.600 758.890 2518.860 759.035 ;
        RECT 2763.780 758.890 2764.040 759.210 ;
        RECT 2763.840 38.070 2763.980 758.890 ;
        RECT 2763.780 37.750 2764.040 38.070 ;
        RECT 2821.740 37.750 2822.000 38.070 ;
        RECT 2821.800 2.400 2821.940 37.750 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 2518.590 759.080 2518.870 759.360 ;
      LAYER met3 ;
        RECT 2506.000 759.370 2510.000 759.520 ;
        RECT 2518.565 759.370 2518.895 759.385 ;
        RECT 2506.000 759.070 2518.895 759.370 ;
        RECT 2506.000 758.920 2510.000 759.070 ;
        RECT 2518.565 759.055 2518.895 759.070 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 395.670 472.500 395.990 472.560 ;
        RECT 2835.970 472.500 2836.290 472.560 ;
        RECT 395.670 472.360 2836.290 472.500 ;
        RECT 395.670 472.300 395.990 472.360 ;
        RECT 2835.970 472.300 2836.290 472.360 ;
      LAYER via ;
        RECT 395.700 472.300 395.960 472.560 ;
        RECT 2836.000 472.300 2836.260 472.560 ;
      LAYER met2 ;
        RECT 395.690 568.635 395.970 569.005 ;
        RECT 395.760 472.590 395.900 568.635 ;
        RECT 395.700 472.270 395.960 472.590 ;
        RECT 2836.000 472.270 2836.260 472.590 ;
        RECT 2836.060 16.730 2836.200 472.270 ;
        RECT 2836.060 16.590 2839.420 16.730 ;
        RECT 2839.280 2.400 2839.420 16.590 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
      LAYER via2 ;
        RECT 395.690 568.680 395.970 568.960 ;
      LAYER met3 ;
        RECT 395.665 568.970 395.995 568.985 ;
        RECT 410.000 568.970 414.000 569.120 ;
        RECT 395.665 568.670 414.000 568.970 ;
        RECT 395.665 568.655 395.995 568.670 ;
        RECT 410.000 568.520 414.000 568.670 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2522.710 517.720 2523.030 517.780 ;
        RECT 2556.750 517.720 2557.070 517.780 ;
        RECT 2522.710 517.580 2557.070 517.720 ;
        RECT 2522.710 517.520 2523.030 517.580 ;
        RECT 2556.750 517.520 2557.070 517.580 ;
        RECT 2556.750 59.400 2557.070 59.460 ;
        RECT 2856.670 59.400 2856.990 59.460 ;
        RECT 2556.750 59.260 2856.990 59.400 ;
        RECT 2556.750 59.200 2557.070 59.260 ;
        RECT 2856.670 59.200 2856.990 59.260 ;
      LAYER via ;
        RECT 2522.740 517.520 2523.000 517.780 ;
        RECT 2556.780 517.520 2557.040 517.780 ;
        RECT 2556.780 59.200 2557.040 59.460 ;
        RECT 2856.700 59.200 2856.960 59.460 ;
      LAYER met2 ;
        RECT 2522.730 521.035 2523.010 521.405 ;
        RECT 2522.800 517.810 2522.940 521.035 ;
        RECT 2522.740 517.490 2523.000 517.810 ;
        RECT 2556.780 517.490 2557.040 517.810 ;
        RECT 2556.840 59.490 2556.980 517.490 ;
        RECT 2556.780 59.170 2557.040 59.490 ;
        RECT 2856.700 59.170 2856.960 59.490 ;
        RECT 2856.760 17.410 2856.900 59.170 ;
        RECT 2856.760 17.270 2857.360 17.410 ;
        RECT 2857.220 2.400 2857.360 17.270 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 2522.730 521.080 2523.010 521.360 ;
      LAYER met3 ;
        RECT 2506.000 521.370 2510.000 521.520 ;
        RECT 2522.705 521.370 2523.035 521.385 ;
        RECT 2506.000 521.070 2523.035 521.370 ;
        RECT 2506.000 520.920 2510.000 521.070 ;
        RECT 2522.705 521.055 2523.035 521.070 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2912.000 2519.810 2912.060 ;
        RECT 2870.470 2912.000 2870.790 2912.060 ;
        RECT 2519.490 2911.860 2870.790 2912.000 ;
        RECT 2519.490 2911.800 2519.810 2911.860 ;
        RECT 2870.470 2911.800 2870.790 2911.860 ;
      LAYER via ;
        RECT 2519.520 2911.800 2519.780 2912.060 ;
        RECT 2870.500 2911.800 2870.760 2912.060 ;
      LAYER met2 ;
        RECT 2519.510 2913.275 2519.790 2913.645 ;
        RECT 2519.580 2912.090 2519.720 2913.275 ;
        RECT 2519.520 2911.770 2519.780 2912.090 ;
        RECT 2870.500 2911.770 2870.760 2912.090 ;
        RECT 2870.560 16.730 2870.700 2911.770 ;
        RECT 2870.560 16.590 2875.300 16.730 ;
        RECT 2875.160 2.400 2875.300 16.590 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2913.320 2519.790 2913.600 ;
      LAYER met3 ;
        RECT 2506.000 2913.610 2510.000 2913.760 ;
        RECT 2519.485 2913.610 2519.815 2913.625 ;
        RECT 2506.000 2913.310 2519.815 2913.610 ;
        RECT 2506.000 2913.160 2510.000 2913.310 ;
        RECT 2519.485 2913.295 2519.815 2913.310 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.870 938.640 2521.190 938.700 ;
        RECT 2770.190 938.640 2770.510 938.700 ;
        RECT 2520.870 938.500 2770.510 938.640 ;
        RECT 2520.870 938.440 2521.190 938.500 ;
        RECT 2770.190 938.440 2770.510 938.500 ;
        RECT 2770.190 24.040 2770.510 24.100 ;
        RECT 2893.010 24.040 2893.330 24.100 ;
        RECT 2770.190 23.900 2893.330 24.040 ;
        RECT 2770.190 23.840 2770.510 23.900 ;
        RECT 2893.010 23.840 2893.330 23.900 ;
      LAYER via ;
        RECT 2520.900 938.440 2521.160 938.700 ;
        RECT 2770.220 938.440 2770.480 938.700 ;
        RECT 2770.220 23.840 2770.480 24.100 ;
        RECT 2893.040 23.840 2893.300 24.100 ;
      LAYER met2 ;
        RECT 2520.890 941.275 2521.170 941.645 ;
        RECT 2520.960 938.730 2521.100 941.275 ;
        RECT 2520.900 938.410 2521.160 938.730 ;
        RECT 2770.220 938.410 2770.480 938.730 ;
        RECT 2770.280 24.130 2770.420 938.410 ;
        RECT 2770.220 23.810 2770.480 24.130 ;
        RECT 2893.040 23.810 2893.300 24.130 ;
        RECT 2893.100 2.400 2893.240 23.810 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 2520.890 941.320 2521.170 941.600 ;
      LAYER met3 ;
        RECT 2506.000 941.610 2510.000 941.760 ;
        RECT 2520.865 941.610 2521.195 941.625 ;
        RECT 2506.000 941.310 2521.195 941.610 ;
        RECT 2506.000 941.160 2510.000 941.310 ;
        RECT 2520.865 941.295 2521.195 941.310 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 141.340 724.430 141.400 ;
        RECT 2905.430 141.340 2905.750 141.400 ;
        RECT 724.110 141.200 2905.750 141.340 ;
        RECT 724.110 141.140 724.430 141.200 ;
        RECT 2905.430 141.140 2905.750 141.200 ;
        RECT 2905.430 2.960 2905.750 3.020 ;
        RECT 2910.950 2.960 2911.270 3.020 ;
        RECT 2905.430 2.820 2911.270 2.960 ;
        RECT 2905.430 2.760 2905.750 2.820 ;
        RECT 2910.950 2.760 2911.270 2.820 ;
      LAYER via ;
        RECT 724.140 141.140 724.400 141.400 ;
        RECT 2905.460 141.140 2905.720 141.400 ;
        RECT 2905.460 2.760 2905.720 3.020 ;
        RECT 2910.980 2.760 2911.240 3.020 ;
      LAYER met2 ;
        RECT 721.050 510.410 721.330 514.000 ;
        RECT 721.050 510.270 724.340 510.410 ;
        RECT 721.050 510.000 721.330 510.270 ;
        RECT 724.200 141.430 724.340 510.270 ;
        RECT 724.140 141.110 724.400 141.430 ;
        RECT 2905.460 141.110 2905.720 141.430 ;
        RECT 2905.520 3.050 2905.660 141.110 ;
        RECT 2905.460 2.730 2905.720 3.050 ;
        RECT 2910.980 2.730 2911.240 3.050 ;
        RECT 2911.040 2.400 2911.180 2.730 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 382.790 1497.600 383.110 1497.660 ;
        RECT 396.130 1497.600 396.450 1497.660 ;
        RECT 382.790 1497.460 396.450 1497.600 ;
        RECT 382.790 1497.400 383.110 1497.460 ;
        RECT 396.130 1497.400 396.450 1497.460 ;
        RECT 382.790 369.480 383.110 369.540 ;
        RECT 855.670 369.480 855.990 369.540 ;
        RECT 382.790 369.340 855.990 369.480 ;
        RECT 382.790 369.280 383.110 369.340 ;
        RECT 855.670 369.280 855.990 369.340 ;
        RECT 855.670 2.960 855.990 3.020 ;
        RECT 858.890 2.960 859.210 3.020 ;
        RECT 855.670 2.820 859.210 2.960 ;
        RECT 855.670 2.760 855.990 2.820 ;
        RECT 858.890 2.760 859.210 2.820 ;
      LAYER via ;
        RECT 382.820 1497.400 383.080 1497.660 ;
        RECT 396.160 1497.400 396.420 1497.660 ;
        RECT 382.820 369.280 383.080 369.540 ;
        RECT 855.700 369.280 855.960 369.540 ;
        RECT 855.700 2.760 855.960 3.020 ;
        RECT 858.920 2.760 859.180 3.020 ;
      LAYER met2 ;
        RECT 396.150 1500.235 396.430 1500.605 ;
        RECT 396.220 1497.690 396.360 1500.235 ;
        RECT 382.820 1497.370 383.080 1497.690 ;
        RECT 396.160 1497.370 396.420 1497.690 ;
        RECT 382.880 369.570 383.020 1497.370 ;
        RECT 382.820 369.250 383.080 369.570 ;
        RECT 855.700 369.250 855.960 369.570 ;
        RECT 855.760 3.050 855.900 369.250 ;
        RECT 855.700 2.730 855.960 3.050 ;
        RECT 858.920 2.730 859.180 3.050 ;
        RECT 858.980 2.400 859.120 2.730 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 396.150 1500.280 396.430 1500.560 ;
      LAYER met3 ;
        RECT 396.125 1500.570 396.455 1500.585 ;
        RECT 410.000 1500.570 414.000 1500.720 ;
        RECT 396.125 1500.270 414.000 1500.570 ;
        RECT 396.125 1500.255 396.455 1500.270 ;
        RECT 410.000 1500.120 414.000 1500.270 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2125.805 3001.265 2125.975 3006.535 ;
      LAYER mcon ;
        RECT 2125.805 3006.365 2125.975 3006.535 ;
      LAYER met1 ;
        RECT 2125.730 3006.520 2126.050 3006.580 ;
        RECT 2125.535 3006.380 2126.050 3006.520 ;
        RECT 2125.730 3006.320 2126.050 3006.380 ;
        RECT 2125.745 3001.420 2126.035 3001.465 ;
        RECT 2507.530 3001.420 2507.850 3001.480 ;
        RECT 2125.745 3001.280 2507.850 3001.420 ;
        RECT 2125.745 3001.235 2126.035 3001.280 ;
        RECT 2507.530 3001.220 2507.850 3001.280 ;
        RECT 876.830 16.560 877.150 16.620 ;
        RECT 882.810 16.560 883.130 16.620 ;
        RECT 876.830 16.420 883.130 16.560 ;
        RECT 876.830 16.360 877.150 16.420 ;
        RECT 882.810 16.360 883.130 16.420 ;
      LAYER via ;
        RECT 2125.760 3006.320 2126.020 3006.580 ;
        RECT 2507.560 3001.220 2507.820 3001.480 ;
        RECT 876.860 16.360 877.120 16.620 ;
        RECT 882.840 16.360 883.100 16.620 ;
      LAYER met2 ;
        RECT 2124.050 3006.690 2124.330 3010.000 ;
        RECT 2124.050 3006.610 2125.960 3006.690 ;
        RECT 2124.050 3006.550 2126.020 3006.610 ;
        RECT 2124.050 3006.000 2124.330 3006.550 ;
        RECT 2125.760 3006.290 2126.020 3006.550 ;
        RECT 2507.560 3001.365 2507.820 3001.510 ;
        RECT 2507.550 3000.995 2507.830 3001.365 ;
        RECT 882.830 506.755 883.110 507.125 ;
        RECT 882.900 16.650 883.040 506.755 ;
        RECT 876.860 16.330 877.120 16.650 ;
        RECT 882.840 16.330 883.100 16.650 ;
        RECT 876.920 2.400 877.060 16.330 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 2507.550 3001.040 2507.830 3001.320 ;
        RECT 882.830 506.800 883.110 507.080 ;
      LAYER met3 ;
        RECT 2498.990 3001.330 2499.370 3001.340 ;
        RECT 2507.525 3001.330 2507.855 3001.345 ;
        RECT 2498.990 3001.030 2507.855 3001.330 ;
        RECT 2498.990 3001.020 2499.370 3001.030 ;
        RECT 2507.525 3001.015 2507.855 3001.030 ;
        RECT 882.805 507.090 883.135 507.105 ;
        RECT 2468.630 507.090 2469.010 507.100 ;
        RECT 882.805 506.790 2469.010 507.090 ;
        RECT 882.805 506.775 883.135 506.790 ;
        RECT 2468.630 506.780 2469.010 506.790 ;
      LAYER via3 ;
        RECT 2499.020 3001.020 2499.340 3001.340 ;
        RECT 2468.660 506.780 2468.980 507.100 ;
      LAYER met4 ;
        RECT 2499.015 3001.015 2499.345 3001.345 ;
        RECT 2499.030 2538.690 2499.330 3001.015 ;
        RECT 2471.910 2537.510 2473.090 2538.690 ;
        RECT 2498.590 2537.510 2499.770 2538.690 ;
        RECT 2472.350 2382.290 2472.650 2537.510 ;
        RECT 2467.310 2381.110 2468.490 2382.290 ;
        RECT 2471.910 2381.110 2473.090 2382.290 ;
        RECT 2467.750 2347.850 2468.050 2381.110 ;
        RECT 2467.750 2347.550 2472.650 2347.850 ;
        RECT 2472.350 2279.850 2472.650 2347.550 ;
        RECT 2470.510 2279.550 2472.650 2279.850 ;
        RECT 2470.510 2256.490 2470.810 2279.550 ;
        RECT 2470.070 2255.310 2471.250 2256.490 ;
        RECT 2470.070 2242.450 2471.250 2242.890 ;
        RECT 2467.750 2242.150 2471.250 2242.450 ;
        RECT 2467.750 2201.650 2468.050 2242.150 ;
        RECT 2470.070 2241.710 2471.250 2242.150 ;
        RECT 2467.750 2201.350 2470.810 2201.650 ;
        RECT 2470.510 2147.250 2470.810 2201.350 ;
        RECT 2468.670 2146.950 2470.810 2147.250 ;
        RECT 2468.670 2086.050 2468.970 2146.950 ;
        RECT 2468.670 2085.750 2471.730 2086.050 ;
        RECT 2471.430 2035.050 2471.730 2085.750 ;
        RECT 2467.750 2034.750 2471.730 2035.050 ;
        RECT 2467.750 1984.490 2468.050 2034.750 ;
        RECT 2467.310 1983.310 2468.490 1984.490 ;
        RECT 2471.910 1983.310 2473.090 1984.490 ;
        RECT 2472.350 1878.650 2472.650 1983.310 ;
        RECT 2471.430 1878.350 2472.650 1878.650 ;
        RECT 2471.430 1871.850 2471.730 1878.350 ;
        RECT 2471.430 1871.550 2472.650 1871.850 ;
        RECT 2472.350 1810.650 2472.650 1871.550 ;
        RECT 2470.510 1810.350 2472.650 1810.650 ;
        RECT 2470.510 1766.450 2470.810 1810.350 ;
        RECT 2470.510 1766.150 2471.730 1766.450 ;
        RECT 2471.430 1701.850 2471.730 1766.150 ;
        RECT 2471.430 1701.550 2474.490 1701.850 ;
        RECT 2474.190 1678.050 2474.490 1701.550 ;
        RECT 2474.190 1677.750 2476.330 1678.050 ;
        RECT 2476.030 1667.850 2476.330 1677.750 ;
        RECT 2471.430 1667.550 2476.330 1667.850 ;
        RECT 2471.430 1610.490 2471.730 1667.550 ;
        RECT 2466.390 1609.310 2467.570 1610.490 ;
        RECT 2470.990 1609.310 2472.170 1610.490 ;
        RECT 2466.830 1593.050 2467.130 1609.310 ;
        RECT 2466.830 1592.750 2472.650 1593.050 ;
        RECT 2472.350 1545.450 2472.650 1592.750 ;
        RECT 2470.510 1545.150 2472.650 1545.450 ;
        RECT 2470.510 1498.290 2470.810 1545.150 ;
        RECT 2470.070 1497.110 2471.250 1498.290 ;
        RECT 2475.590 1497.110 2476.770 1498.290 ;
        RECT 2476.030 1409.450 2476.330 1497.110 ;
        RECT 2475.110 1409.150 2476.330 1409.450 ;
        RECT 2475.110 1406.050 2475.410 1409.150 ;
        RECT 2471.430 1405.750 2475.410 1406.050 ;
        RECT 2471.430 1375.450 2471.730 1405.750 ;
        RECT 2471.430 1375.150 2472.650 1375.450 ;
        RECT 2472.350 1351.650 2472.650 1375.150 ;
        RECT 2471.430 1351.350 2472.650 1351.650 ;
        RECT 2471.430 1327.850 2471.730 1351.350 ;
        RECT 2469.590 1327.550 2471.730 1327.850 ;
        RECT 2469.590 1317.650 2469.890 1327.550 ;
        RECT 2469.590 1317.350 2471.730 1317.650 ;
        RECT 2471.430 1297.690 2471.730 1317.350 ;
        RECT 2470.990 1296.510 2472.170 1297.690 ;
        RECT 2484.790 1296.510 2485.970 1297.690 ;
        RECT 2485.230 1267.090 2485.530 1296.510 ;
        RECT 2466.390 1265.910 2467.570 1267.090 ;
        RECT 2484.790 1265.910 2485.970 1267.090 ;
        RECT 2466.830 1239.450 2467.130 1265.910 ;
        RECT 2466.830 1239.150 2472.650 1239.450 ;
        RECT 2472.350 1212.250 2472.650 1239.150 ;
        RECT 2467.750 1211.950 2472.650 1212.250 ;
        RECT 2467.750 1188.890 2468.050 1211.950 ;
        RECT 2467.310 1187.710 2468.490 1188.890 ;
        RECT 2471.910 1187.710 2473.090 1188.890 ;
        RECT 2472.350 1086.890 2472.650 1187.710 ;
        RECT 2468.230 1085.710 2469.410 1086.890 ;
        RECT 2471.910 1085.710 2473.090 1086.890 ;
        RECT 2468.670 1066.050 2468.970 1085.710 ;
        RECT 2468.670 1065.750 2472.650 1066.050 ;
        RECT 2472.350 1042.250 2472.650 1065.750 ;
        RECT 2471.430 1041.950 2472.650 1042.250 ;
        RECT 2471.430 981.050 2471.730 1041.950 ;
        RECT 2471.430 980.750 2472.650 981.050 ;
        RECT 2472.350 902.850 2472.650 980.750 ;
        RECT 2470.510 902.550 2472.650 902.850 ;
        RECT 2470.510 899.890 2470.810 902.550 ;
        RECT 2470.070 898.710 2471.250 899.890 ;
        RECT 2471.910 885.110 2473.090 886.290 ;
        RECT 2472.350 511.850 2472.650 885.110 ;
        RECT 2468.670 511.550 2472.650 511.850 ;
        RECT 2468.670 507.105 2468.970 511.550 ;
        RECT 2468.655 506.775 2468.985 507.105 ;
      LAYER met5 ;
        RECT 2471.700 2537.300 2499.980 2538.900 ;
        RECT 2467.100 2380.900 2473.300 2382.500 ;
        RECT 2469.860 2255.100 2473.300 2256.700 ;
        RECT 2471.700 2243.100 2473.300 2255.100 ;
        RECT 2469.860 2241.500 2473.300 2243.100 ;
        RECT 2467.100 1983.100 2473.300 1984.700 ;
        RECT 2466.180 1609.100 2472.380 1610.700 ;
        RECT 2469.860 1496.900 2476.980 1498.500 ;
        RECT 2470.780 1296.300 2486.180 1297.900 ;
        RECT 2466.180 1265.700 2486.180 1267.300 ;
        RECT 2467.100 1187.500 2473.300 1189.100 ;
        RECT 2468.020 1085.500 2473.300 1087.100 ;
        RECT 2469.860 898.500 2473.300 900.100 ;
        RECT 2471.700 884.900 2473.300 898.500 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 37.980 895.090 38.040 ;
        RECT 2214.970 37.980 2215.290 38.040 ;
        RECT 894.770 37.840 2215.290 37.980 ;
        RECT 894.770 37.780 895.090 37.840 ;
        RECT 2214.970 37.780 2215.290 37.840 ;
      LAYER via ;
        RECT 894.800 37.780 895.060 38.040 ;
        RECT 2215.000 37.780 2215.260 38.040 ;
      LAYER met2 ;
        RECT 2216.050 510.410 2216.330 514.000 ;
        RECT 2215.060 510.270 2216.330 510.410 ;
        RECT 2215.060 38.070 2215.200 510.270 ;
        RECT 2216.050 510.000 2216.330 510.270 ;
        RECT 894.800 37.750 895.060 38.070 ;
        RECT 2215.000 37.750 2215.260 38.070 ;
        RECT 894.860 2.400 895.000 37.750 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1249.060 2520.730 1249.120 ;
        RECT 2590.330 1249.060 2590.650 1249.120 ;
        RECT 2520.410 1248.920 2590.650 1249.060 ;
        RECT 2520.410 1248.860 2520.730 1248.920 ;
        RECT 2590.330 1248.860 2590.650 1248.920 ;
        RECT 917.310 466.040 917.630 466.100 ;
        RECT 2590.330 466.040 2590.650 466.100 ;
        RECT 917.310 465.900 2590.650 466.040 ;
        RECT 917.310 465.840 917.630 465.900 ;
        RECT 2590.330 465.840 2590.650 465.900 ;
        RECT 912.710 16.560 913.030 16.620 ;
        RECT 917.310 16.560 917.630 16.620 ;
        RECT 912.710 16.420 917.630 16.560 ;
        RECT 912.710 16.360 913.030 16.420 ;
        RECT 917.310 16.360 917.630 16.420 ;
      LAYER via ;
        RECT 2520.440 1248.860 2520.700 1249.120 ;
        RECT 2590.360 1248.860 2590.620 1249.120 ;
        RECT 917.340 465.840 917.600 466.100 ;
        RECT 2590.360 465.840 2590.620 466.100 ;
        RECT 912.740 16.360 913.000 16.620 ;
        RECT 917.340 16.360 917.600 16.620 ;
      LAYER met2 ;
        RECT 2520.430 1251.355 2520.710 1251.725 ;
        RECT 2520.500 1249.150 2520.640 1251.355 ;
        RECT 2520.440 1248.830 2520.700 1249.150 ;
        RECT 2590.360 1248.830 2590.620 1249.150 ;
        RECT 2590.420 466.130 2590.560 1248.830 ;
        RECT 917.340 465.810 917.600 466.130 ;
        RECT 2590.360 465.810 2590.620 466.130 ;
        RECT 917.400 16.650 917.540 465.810 ;
        RECT 912.740 16.330 913.000 16.650 ;
        RECT 917.340 16.330 917.600 16.650 ;
        RECT 912.800 2.400 912.940 16.330 ;
        RECT 912.590 -4.800 913.150 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1251.400 2520.710 1251.680 ;
      LAYER met3 ;
        RECT 2506.000 1251.690 2510.000 1251.840 ;
        RECT 2520.405 1251.690 2520.735 1251.705 ;
        RECT 2506.000 1251.390 2520.735 1251.690 ;
        RECT 2506.000 1251.240 2510.000 1251.390 ;
        RECT 2520.405 1251.375 2520.735 1251.390 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1338.820 2520.730 1338.880 ;
        RECT 2576.530 1338.820 2576.850 1338.880 ;
        RECT 2520.410 1338.680 2576.850 1338.820 ;
        RECT 2520.410 1338.620 2520.730 1338.680 ;
        RECT 2576.530 1338.620 2576.850 1338.680 ;
        RECT 931.110 466.380 931.430 466.440 ;
        RECT 2576.530 466.380 2576.850 466.440 ;
        RECT 931.110 466.240 2576.850 466.380 ;
        RECT 931.110 466.180 931.430 466.240 ;
        RECT 2576.530 466.180 2576.850 466.240 ;
      LAYER via ;
        RECT 2520.440 1338.620 2520.700 1338.880 ;
        RECT 2576.560 1338.620 2576.820 1338.880 ;
        RECT 931.140 466.180 931.400 466.440 ;
        RECT 2576.560 466.180 2576.820 466.440 ;
      LAYER met2 ;
        RECT 2520.430 1343.835 2520.710 1344.205 ;
        RECT 2520.500 1338.910 2520.640 1343.835 ;
        RECT 2520.440 1338.590 2520.700 1338.910 ;
        RECT 2576.560 1338.590 2576.820 1338.910 ;
        RECT 2576.620 466.470 2576.760 1338.590 ;
        RECT 931.140 466.150 931.400 466.470 ;
        RECT 2576.560 466.150 2576.820 466.470 ;
        RECT 931.200 3.130 931.340 466.150 ;
        RECT 930.280 2.990 931.340 3.130 ;
        RECT 930.280 2.400 930.420 2.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1343.880 2520.710 1344.160 ;
      LAYER met3 ;
        RECT 2506.000 1344.170 2510.000 1344.320 ;
        RECT 2520.405 1344.170 2520.735 1344.185 ;
        RECT 2506.000 1343.870 2520.735 1344.170 ;
        RECT 2506.000 1343.720 2510.000 1343.870 ;
        RECT 2520.405 1343.855 2520.735 1343.870 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 16.900 948.450 16.960 ;
        RECT 951.810 16.900 952.130 16.960 ;
        RECT 948.130 16.760 952.130 16.900 ;
        RECT 948.130 16.700 948.450 16.760 ;
        RECT 951.810 16.700 952.130 16.760 ;
      LAYER via ;
        RECT 948.160 16.700 948.420 16.960 ;
        RECT 951.840 16.700 952.100 16.960 ;
      LAYER met2 ;
        RECT 951.830 230.675 952.110 231.045 ;
        RECT 951.900 16.990 952.040 230.675 ;
        RECT 948.160 16.670 948.420 16.990 ;
        RECT 951.840 16.670 952.100 16.990 ;
        RECT 948.220 2.400 948.360 16.670 ;
        RECT 948.010 -4.800 948.570 2.400 ;
      LAYER via2 ;
        RECT 951.830 230.720 952.110 231.000 ;
      LAYER met3 ;
        RECT 2506.000 2330.170 2510.000 2330.320 ;
        RECT 2533.030 2330.170 2533.410 2330.180 ;
        RECT 2506.000 2329.870 2533.410 2330.170 ;
        RECT 2506.000 2329.720 2510.000 2329.870 ;
        RECT 2533.030 2329.860 2533.410 2329.870 ;
        RECT 951.805 231.010 952.135 231.025 ;
        RECT 2533.030 231.010 2533.410 231.020 ;
        RECT 951.805 230.710 2533.410 231.010 ;
        RECT 951.805 230.695 952.135 230.710 ;
        RECT 2533.030 230.700 2533.410 230.710 ;
      LAYER via3 ;
        RECT 2533.060 2329.860 2533.380 2330.180 ;
        RECT 2533.060 230.700 2533.380 231.020 ;
      LAYER met4 ;
        RECT 2533.055 2329.855 2533.385 2330.185 ;
        RECT 2533.070 231.025 2533.370 2329.855 ;
        RECT 2533.055 230.695 2533.385 231.025 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 399.810 3023.860 400.130 3023.920 ;
        RECT 1629.850 3023.860 1630.170 3023.920 ;
        RECT 399.810 3023.720 1630.170 3023.860 ;
        RECT 399.810 3023.660 400.130 3023.720 ;
        RECT 1629.850 3023.660 1630.170 3023.720 ;
        RECT 399.810 883.560 400.130 883.620 ;
        RECT 403.490 883.560 403.810 883.620 ;
        RECT 399.810 883.420 403.810 883.560 ;
        RECT 399.810 883.360 400.130 883.420 ;
        RECT 403.490 883.360 403.810 883.420 ;
        RECT 403.490 494.600 403.810 494.660 ;
        RECT 966.070 494.600 966.390 494.660 ;
        RECT 403.490 494.460 966.390 494.600 ;
        RECT 403.490 494.400 403.810 494.460 ;
        RECT 966.070 494.400 966.390 494.460 ;
      LAYER via ;
        RECT 399.840 3023.660 400.100 3023.920 ;
        RECT 1629.880 3023.660 1630.140 3023.920 ;
        RECT 399.840 883.360 400.100 883.620 ;
        RECT 403.520 883.360 403.780 883.620 ;
        RECT 403.520 494.400 403.780 494.660 ;
        RECT 966.100 494.400 966.360 494.660 ;
      LAYER met2 ;
        RECT 399.840 3023.630 400.100 3023.950 ;
        RECT 1629.880 3023.630 1630.140 3023.950 ;
        RECT 399.900 883.650 400.040 3023.630 ;
        RECT 1629.940 3010.000 1630.080 3023.630 ;
        RECT 1629.940 3009.340 1630.290 3010.000 ;
        RECT 1630.010 3006.000 1630.290 3009.340 ;
        RECT 399.840 883.330 400.100 883.650 ;
        RECT 403.520 883.330 403.780 883.650 ;
        RECT 403.580 494.690 403.720 883.330 ;
        RECT 403.520 494.370 403.780 494.690 ;
        RECT 966.100 494.370 966.360 494.690 ;
        RECT 966.160 2.400 966.300 494.370 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.690 493.920 390.010 493.980 ;
        RECT 979.870 493.920 980.190 493.980 ;
        RECT 389.690 493.780 980.190 493.920 ;
        RECT 389.690 493.720 390.010 493.780 ;
        RECT 979.870 493.720 980.190 493.780 ;
        RECT 979.870 2.960 980.190 3.020 ;
        RECT 984.010 2.960 984.330 3.020 ;
        RECT 979.870 2.820 984.330 2.960 ;
        RECT 979.870 2.760 980.190 2.820 ;
        RECT 984.010 2.760 984.330 2.820 ;
      LAYER via ;
        RECT 389.720 493.720 389.980 493.980 ;
        RECT 979.900 493.720 980.160 493.980 ;
        RECT 979.900 2.760 980.160 3.020 ;
        RECT 984.040 2.760 984.300 3.020 ;
      LAYER met2 ;
        RECT 389.710 988.875 389.990 989.245 ;
        RECT 389.780 494.010 389.920 988.875 ;
        RECT 389.720 493.690 389.980 494.010 ;
        RECT 979.900 493.690 980.160 494.010 ;
        RECT 979.960 3.050 980.100 493.690 ;
        RECT 979.900 2.730 980.160 3.050 ;
        RECT 984.040 2.730 984.300 3.050 ;
        RECT 984.100 2.400 984.240 2.730 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 389.710 988.920 389.990 989.200 ;
      LAYER met3 ;
        RECT 389.685 989.210 390.015 989.225 ;
        RECT 410.000 989.210 414.000 989.360 ;
        RECT 389.685 988.910 414.000 989.210 ;
        RECT 389.685 988.895 390.015 988.910 ;
        RECT 410.000 988.760 414.000 988.910 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 391.990 496.300 392.310 496.360 ;
        RECT 662.930 496.300 663.250 496.360 ;
        RECT 391.990 496.160 663.250 496.300 ;
        RECT 391.990 496.100 392.310 496.160 ;
        RECT 662.930 496.100 663.250 496.160 ;
      LAYER via ;
        RECT 392.020 496.100 392.280 496.360 ;
        RECT 662.960 496.100 663.220 496.360 ;
      LAYER met2 ;
        RECT 392.010 1974.875 392.290 1975.245 ;
        RECT 392.080 496.390 392.220 1974.875 ;
        RECT 392.020 496.070 392.280 496.390 ;
        RECT 662.960 496.070 663.220 496.390 ;
        RECT 663.020 2.400 663.160 496.070 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 392.010 1974.920 392.290 1975.200 ;
      LAYER met3 ;
        RECT 391.985 1975.210 392.315 1975.225 ;
        RECT 410.000 1975.210 414.000 1975.360 ;
        RECT 391.985 1974.910 414.000 1975.210 ;
        RECT 391.985 1974.895 392.315 1974.910 ;
        RECT 410.000 1974.760 414.000 1974.910 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 432.040 1007.330 432.100 ;
        RECT 1373.170 432.040 1373.490 432.100 ;
        RECT 1007.010 431.900 1373.490 432.040 ;
        RECT 1007.010 431.840 1007.330 431.900 ;
        RECT 1373.170 431.840 1373.490 431.900 ;
        RECT 1001.950 15.880 1002.270 15.940 ;
        RECT 1007.010 15.880 1007.330 15.940 ;
        RECT 1001.950 15.740 1007.330 15.880 ;
        RECT 1001.950 15.680 1002.270 15.740 ;
        RECT 1007.010 15.680 1007.330 15.740 ;
      LAYER via ;
        RECT 1007.040 431.840 1007.300 432.100 ;
        RECT 1373.200 431.840 1373.460 432.100 ;
        RECT 1001.980 15.680 1002.240 15.940 ;
        RECT 1007.040 15.680 1007.300 15.940 ;
      LAYER met2 ;
        RECT 1376.090 510.410 1376.370 514.000 ;
        RECT 1373.260 510.270 1376.370 510.410 ;
        RECT 1373.260 432.130 1373.400 510.270 ;
        RECT 1376.090 510.000 1376.370 510.270 ;
        RECT 1007.040 431.810 1007.300 432.130 ;
        RECT 1373.200 431.810 1373.460 432.130 ;
        RECT 1007.100 15.970 1007.240 431.810 ;
        RECT 1001.980 15.650 1002.240 15.970 ;
        RECT 1007.040 15.650 1007.300 15.970 ;
        RECT 1002.040 2.400 1002.180 15.650 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1019.505 2.805 1019.675 14.195 ;
      LAYER mcon ;
        RECT 1019.505 14.025 1019.675 14.195 ;
      LAYER met1 ;
        RECT 2519.950 1835.560 2520.270 1835.620 ;
        RECT 2534.210 1835.560 2534.530 1835.620 ;
        RECT 2519.950 1835.420 2534.530 1835.560 ;
        RECT 2519.950 1835.360 2520.270 1835.420 ;
        RECT 2534.210 1835.360 2534.530 1835.420 ;
        RECT 1020.350 148.140 1020.670 148.200 ;
        RECT 2534.210 148.140 2534.530 148.200 ;
        RECT 1020.350 148.000 2534.530 148.140 ;
        RECT 1020.350 147.940 1020.670 148.000 ;
        RECT 2534.210 147.940 2534.530 148.000 ;
        RECT 1019.445 14.180 1019.735 14.225 ;
        RECT 1020.350 14.180 1020.670 14.240 ;
        RECT 1019.445 14.040 1020.670 14.180 ;
        RECT 1019.445 13.995 1019.735 14.040 ;
        RECT 1020.350 13.980 1020.670 14.040 ;
        RECT 1019.430 2.960 1019.750 3.020 ;
        RECT 1019.235 2.820 1019.750 2.960 ;
        RECT 1019.430 2.760 1019.750 2.820 ;
      LAYER via ;
        RECT 2519.980 1835.360 2520.240 1835.620 ;
        RECT 2534.240 1835.360 2534.500 1835.620 ;
        RECT 1020.380 147.940 1020.640 148.200 ;
        RECT 2534.240 147.940 2534.500 148.200 ;
        RECT 1020.380 13.980 1020.640 14.240 ;
        RECT 1019.460 2.760 1019.720 3.020 ;
      LAYER met2 ;
        RECT 2519.970 1836.155 2520.250 1836.525 ;
        RECT 2520.040 1835.650 2520.180 1836.155 ;
        RECT 2519.980 1835.330 2520.240 1835.650 ;
        RECT 2534.240 1835.330 2534.500 1835.650 ;
        RECT 2534.300 148.230 2534.440 1835.330 ;
        RECT 1020.380 147.910 1020.640 148.230 ;
        RECT 2534.240 147.910 2534.500 148.230 ;
        RECT 1020.440 14.270 1020.580 147.910 ;
        RECT 1020.380 13.950 1020.640 14.270 ;
        RECT 1019.460 2.730 1019.720 3.050 ;
        RECT 1019.520 2.400 1019.660 2.730 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 2519.970 1836.200 2520.250 1836.480 ;
      LAYER met3 ;
        RECT 2506.000 1836.490 2510.000 1836.640 ;
        RECT 2519.945 1836.490 2520.275 1836.505 ;
        RECT 2506.000 1836.190 2520.275 1836.490 ;
        RECT 2506.000 1836.040 2510.000 1836.190 ;
        RECT 2519.945 1836.175 2520.275 1836.190 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 405.790 3031.680 406.110 3031.740 ;
        RECT 1593.050 3031.680 1593.370 3031.740 ;
        RECT 405.790 3031.540 1593.370 3031.680 ;
        RECT 405.790 3031.480 406.110 3031.540 ;
        RECT 1593.050 3031.480 1593.370 3031.540 ;
        RECT 405.790 493.240 406.110 493.300 ;
        RECT 1035.070 493.240 1035.390 493.300 ;
        RECT 405.790 493.100 1035.390 493.240 ;
        RECT 405.790 493.040 406.110 493.100 ;
        RECT 1035.070 493.040 1035.390 493.100 ;
        RECT 1035.070 20.300 1035.390 20.360 ;
        RECT 1037.370 20.300 1037.690 20.360 ;
        RECT 1035.070 20.160 1037.690 20.300 ;
        RECT 1035.070 20.100 1035.390 20.160 ;
        RECT 1037.370 20.100 1037.690 20.160 ;
      LAYER via ;
        RECT 405.820 3031.480 406.080 3031.740 ;
        RECT 1593.080 3031.480 1593.340 3031.740 ;
        RECT 405.820 493.040 406.080 493.300 ;
        RECT 1035.100 493.040 1035.360 493.300 ;
        RECT 1035.100 20.100 1035.360 20.360 ;
        RECT 1037.400 20.100 1037.660 20.360 ;
      LAYER met2 ;
        RECT 405.820 3031.450 406.080 3031.770 ;
        RECT 1593.080 3031.450 1593.340 3031.770 ;
        RECT 405.880 493.330 406.020 3031.450 ;
        RECT 1593.140 3010.000 1593.280 3031.450 ;
        RECT 1593.140 3009.340 1593.490 3010.000 ;
        RECT 1593.210 3006.000 1593.490 3009.340 ;
        RECT 405.820 493.010 406.080 493.330 ;
        RECT 1035.100 493.010 1035.360 493.330 ;
        RECT 1035.160 20.390 1035.300 493.010 ;
        RECT 1035.100 20.070 1035.360 20.390 ;
        RECT 1037.400 20.070 1037.660 20.390 ;
        RECT 1037.460 2.400 1037.600 20.070 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1054.925 234.685 1055.095 241.655 ;
        RECT 1054.925 96.305 1055.095 137.955 ;
      LAYER mcon ;
        RECT 1054.925 241.485 1055.095 241.655 ;
        RECT 1054.925 137.785 1055.095 137.955 ;
      LAYER met1 ;
        RECT 1054.850 327.660 1055.170 327.720 ;
        RECT 2520.410 327.660 2520.730 327.720 ;
        RECT 1054.850 327.520 2520.730 327.660 ;
        RECT 1054.850 327.460 1055.170 327.520 ;
        RECT 2520.410 327.460 2520.730 327.520 ;
        RECT 1054.850 241.640 1055.170 241.700 ;
        RECT 1054.655 241.500 1055.170 241.640 ;
        RECT 1054.850 241.440 1055.170 241.500 ;
        RECT 1054.850 234.840 1055.170 234.900 ;
        RECT 1054.655 234.700 1055.170 234.840 ;
        RECT 1054.850 234.640 1055.170 234.700 ;
        RECT 1054.850 186.560 1055.170 186.620 ;
        RECT 1055.310 186.560 1055.630 186.620 ;
        RECT 1054.850 186.420 1055.630 186.560 ;
        RECT 1054.850 186.360 1055.170 186.420 ;
        RECT 1055.310 186.360 1055.630 186.420 ;
        RECT 1054.850 137.940 1055.170 138.000 ;
        RECT 1054.655 137.800 1055.170 137.940 ;
        RECT 1054.850 137.740 1055.170 137.800 ;
        RECT 1054.865 96.460 1055.155 96.505 ;
        RECT 1055.770 96.460 1056.090 96.520 ;
        RECT 1054.865 96.320 1056.090 96.460 ;
        RECT 1054.865 96.275 1055.155 96.320 ;
        RECT 1055.770 96.260 1056.090 96.320 ;
      LAYER via ;
        RECT 1054.880 327.460 1055.140 327.720 ;
        RECT 2520.440 327.460 2520.700 327.720 ;
        RECT 1054.880 241.440 1055.140 241.700 ;
        RECT 1054.880 234.640 1055.140 234.900 ;
        RECT 1054.880 186.360 1055.140 186.620 ;
        RECT 1055.340 186.360 1055.600 186.620 ;
        RECT 1054.880 137.740 1055.140 138.000 ;
        RECT 1055.800 96.260 1056.060 96.520 ;
      LAYER met2 ;
        RECT 2520.430 1014.715 2520.710 1015.085 ;
        RECT 2520.500 327.750 2520.640 1014.715 ;
        RECT 1054.880 327.430 1055.140 327.750 ;
        RECT 2520.440 327.430 2520.700 327.750 ;
        RECT 1054.940 241.730 1055.080 327.430 ;
        RECT 1054.880 241.410 1055.140 241.730 ;
        RECT 1054.880 234.610 1055.140 234.930 ;
        RECT 1054.940 234.330 1055.080 234.610 ;
        RECT 1054.940 234.190 1055.540 234.330 ;
        RECT 1055.400 186.650 1055.540 234.190 ;
        RECT 1054.880 186.330 1055.140 186.650 ;
        RECT 1055.340 186.330 1055.600 186.650 ;
        RECT 1054.940 138.030 1055.080 186.330 ;
        RECT 1054.880 137.710 1055.140 138.030 ;
        RECT 1055.800 96.230 1056.060 96.550 ;
        RECT 1055.860 24.380 1056.000 96.230 ;
        RECT 1055.400 24.240 1056.000 24.380 ;
        RECT 1055.400 2.400 1055.540 24.240 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1014.760 2520.710 1015.040 ;
      LAYER met3 ;
        RECT 2506.000 1015.050 2510.000 1015.200 ;
        RECT 2520.405 1015.050 2520.735 1015.065 ;
        RECT 2506.000 1014.750 2520.735 1015.050 ;
        RECT 2506.000 1014.600 2510.000 1014.750 ;
        RECT 2520.405 1014.735 2520.735 1014.750 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1069.570 62.120 1069.890 62.180 ;
        RECT 1073.250 62.120 1073.570 62.180 ;
        RECT 1069.570 61.980 1073.570 62.120 ;
        RECT 1069.570 61.920 1069.890 61.980 ;
        RECT 1073.250 61.920 1073.570 61.980 ;
      LAYER via ;
        RECT 1069.600 61.920 1069.860 62.180 ;
        RECT 1073.280 61.920 1073.540 62.180 ;
      LAYER met2 ;
        RECT 1069.590 431.275 1069.870 431.645 ;
        RECT 1069.660 62.210 1069.800 431.275 ;
        RECT 1069.600 61.890 1069.860 62.210 ;
        RECT 1073.280 61.890 1073.540 62.210 ;
        RECT 1073.340 2.400 1073.480 61.890 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 1069.590 431.320 1069.870 431.600 ;
      LAYER met3 ;
        RECT 410.000 2375.960 414.000 2376.560 ;
        RECT 412.470 2375.060 412.770 2375.960 ;
        RECT 412.430 2374.740 412.810 2375.060 ;
        RECT 417.030 431.610 417.410 431.620 ;
        RECT 1069.565 431.610 1069.895 431.625 ;
        RECT 417.030 431.310 1069.895 431.610 ;
        RECT 417.030 431.300 417.410 431.310 ;
        RECT 1069.565 431.295 1069.895 431.310 ;
      LAYER via3 ;
        RECT 412.460 2374.740 412.780 2375.060 ;
        RECT 417.060 431.300 417.380 431.620 ;
      LAYER met4 ;
        RECT 412.455 2375.050 412.785 2375.065 ;
        RECT 412.455 2374.750 414.610 2375.050 ;
        RECT 412.455 2374.735 412.785 2374.750 ;
        RECT 414.310 2368.250 414.610 2374.750 ;
        RECT 414.310 2367.950 417.370 2368.250 ;
        RECT 417.070 431.625 417.370 2367.950 ;
        RECT 417.055 431.295 417.385 431.625 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2235.740 2519.810 2235.800 ;
        RECT 2532.830 2235.740 2533.150 2235.800 ;
        RECT 2519.490 2235.600 2533.150 2235.740 ;
        RECT 2519.490 2235.540 2519.810 2235.600 ;
        RECT 2532.830 2235.540 2533.150 2235.600 ;
        RECT 1096.250 293.320 1096.570 293.380 ;
        RECT 2532.830 293.320 2533.150 293.380 ;
        RECT 1096.250 293.180 2533.150 293.320 ;
        RECT 1096.250 293.120 1096.570 293.180 ;
        RECT 2532.830 293.120 2533.150 293.180 ;
        RECT 1090.730 16.220 1091.050 16.280 ;
        RECT 1096.250 16.220 1096.570 16.280 ;
        RECT 1090.730 16.080 1096.570 16.220 ;
        RECT 1090.730 16.020 1091.050 16.080 ;
        RECT 1096.250 16.020 1096.570 16.080 ;
      LAYER via ;
        RECT 2519.520 2235.540 2519.780 2235.800 ;
        RECT 2532.860 2235.540 2533.120 2235.800 ;
        RECT 1096.280 293.120 1096.540 293.380 ;
        RECT 2532.860 293.120 2533.120 293.380 ;
        RECT 1090.760 16.020 1091.020 16.280 ;
        RECT 1096.280 16.020 1096.540 16.280 ;
      LAYER met2 ;
        RECT 2519.510 2238.715 2519.790 2239.085 ;
        RECT 2519.580 2235.830 2519.720 2238.715 ;
        RECT 2519.520 2235.510 2519.780 2235.830 ;
        RECT 2532.860 2235.510 2533.120 2235.830 ;
        RECT 2532.920 293.410 2533.060 2235.510 ;
        RECT 1096.280 293.090 1096.540 293.410 ;
        RECT 2532.860 293.090 2533.120 293.410 ;
        RECT 1096.340 16.310 1096.480 293.090 ;
        RECT 1090.760 15.990 1091.020 16.310 ;
        RECT 1096.280 15.990 1096.540 16.310 ;
        RECT 1090.820 2.400 1090.960 15.990 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2238.760 2519.790 2239.040 ;
      LAYER met3 ;
        RECT 2506.000 2239.050 2510.000 2239.200 ;
        RECT 2519.485 2239.050 2519.815 2239.065 ;
        RECT 2506.000 2238.750 2519.815 2239.050 ;
        RECT 2506.000 2238.600 2510.000 2238.750 ;
        RECT 2519.485 2238.735 2519.815 2238.750 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 308.280 1110.830 308.340 ;
        RECT 1345.570 308.280 1345.890 308.340 ;
        RECT 1110.510 308.140 1345.890 308.280 ;
        RECT 1110.510 308.080 1110.830 308.140 ;
        RECT 1345.570 308.080 1345.890 308.140 ;
      LAYER via ;
        RECT 1110.540 308.080 1110.800 308.340 ;
        RECT 1345.600 308.080 1345.860 308.340 ;
      LAYER met2 ;
        RECT 1351.250 510.410 1351.530 514.000 ;
        RECT 1345.660 510.270 1351.530 510.410 ;
        RECT 1345.660 308.370 1345.800 510.270 ;
        RECT 1351.250 510.000 1351.530 510.270 ;
        RECT 1110.540 308.050 1110.800 308.370 ;
        RECT 1345.600 308.050 1345.860 308.370 ;
        RECT 1110.600 3.130 1110.740 308.050 ;
        RECT 1108.760 2.990 1110.740 3.130 ;
        RECT 1108.760 2.400 1108.900 2.990 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1030.010 501.400 1030.330 501.460 ;
        RECT 1034.610 501.400 1034.930 501.460 ;
        RECT 1030.010 501.260 1034.930 501.400 ;
        RECT 1030.010 501.200 1030.330 501.260 ;
        RECT 1034.610 501.200 1034.930 501.260 ;
        RECT 1034.610 24.380 1034.930 24.440 ;
        RECT 1126.610 24.380 1126.930 24.440 ;
        RECT 1034.610 24.240 1126.930 24.380 ;
        RECT 1034.610 24.180 1034.930 24.240 ;
        RECT 1126.610 24.180 1126.930 24.240 ;
      LAYER via ;
        RECT 1030.040 501.200 1030.300 501.460 ;
        RECT 1034.640 501.200 1034.900 501.460 ;
        RECT 1034.640 24.180 1034.900 24.440 ;
        RECT 1126.640 24.180 1126.900 24.440 ;
      LAYER met2 ;
        RECT 1030.170 510.340 1030.450 514.000 ;
        RECT 1030.100 510.000 1030.450 510.340 ;
        RECT 1030.100 501.490 1030.240 510.000 ;
        RECT 1030.040 501.170 1030.300 501.490 ;
        RECT 1034.640 501.170 1034.900 501.490 ;
        RECT 1034.700 24.470 1034.840 501.170 ;
        RECT 1034.640 24.150 1034.900 24.470 ;
        RECT 1126.640 24.150 1126.900 24.470 ;
        RECT 1126.700 2.400 1126.840 24.150 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.090 189.960 1144.410 190.020 ;
        RECT 2507.530 189.960 2507.850 190.020 ;
        RECT 1144.090 189.820 2507.850 189.960 ;
        RECT 1144.090 189.760 1144.410 189.820 ;
        RECT 2507.530 189.760 2507.850 189.820 ;
      LAYER via ;
        RECT 1144.120 189.760 1144.380 190.020 ;
        RECT 2507.560 189.760 2507.820 190.020 ;
      LAYER met2 ;
        RECT 2507.550 682.875 2507.830 683.245 ;
        RECT 2507.620 190.050 2507.760 682.875 ;
        RECT 1144.120 189.730 1144.380 190.050 ;
        RECT 2507.560 189.730 2507.820 190.050 ;
        RECT 1144.180 17.410 1144.320 189.730 ;
        RECT 1144.180 17.270 1144.780 17.410 ;
        RECT 1144.640 2.400 1144.780 17.270 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 2507.550 682.920 2507.830 683.200 ;
      LAYER met3 ;
        RECT 2506.000 685.480 2510.000 686.080 ;
        RECT 2507.310 683.225 2507.610 685.480 ;
        RECT 2507.310 682.910 2507.855 683.225 ;
        RECT 2507.525 682.895 2507.855 682.910 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 375.940 1166.030 376.000 ;
        RECT 1546.130 375.940 1546.450 376.000 ;
        RECT 1165.710 375.800 1546.450 375.940 ;
        RECT 1165.710 375.740 1166.030 375.800 ;
        RECT 1546.130 375.740 1546.450 375.800 ;
        RECT 1162.490 16.900 1162.810 16.960 ;
        RECT 1165.710 16.900 1166.030 16.960 ;
        RECT 1162.490 16.760 1166.030 16.900 ;
        RECT 1162.490 16.700 1162.810 16.760 ;
        RECT 1165.710 16.700 1166.030 16.760 ;
      LAYER via ;
        RECT 1165.740 375.740 1166.000 376.000 ;
        RECT 1546.160 375.740 1546.420 376.000 ;
        RECT 1162.520 16.700 1162.780 16.960 ;
        RECT 1165.740 16.700 1166.000 16.960 ;
      LAYER met2 ;
        RECT 1549.050 510.410 1549.330 514.000 ;
        RECT 1546.220 510.270 1549.330 510.410 ;
        RECT 1546.220 376.030 1546.360 510.270 ;
        RECT 1549.050 510.000 1549.330 510.270 ;
        RECT 1165.740 375.710 1166.000 376.030 ;
        RECT 1546.160 375.710 1546.420 376.030 ;
        RECT 1165.800 16.990 1165.940 375.710 ;
        RECT 1162.520 16.670 1162.780 16.990 ;
        RECT 1165.740 16.670 1166.000 16.990 ;
        RECT 1162.580 2.400 1162.720 16.670 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 279.380 683.030 279.440 ;
        RECT 2519.030 279.380 2519.350 279.440 ;
        RECT 682.710 279.240 2519.350 279.380 ;
        RECT 682.710 279.180 683.030 279.240 ;
        RECT 2519.030 279.180 2519.350 279.240 ;
        RECT 680.410 16.900 680.730 16.960 ;
        RECT 682.710 16.900 683.030 16.960 ;
        RECT 680.410 16.760 683.030 16.900 ;
        RECT 680.410 16.700 680.730 16.760 ;
        RECT 682.710 16.700 683.030 16.760 ;
      LAYER via ;
        RECT 682.740 279.180 683.000 279.440 ;
        RECT 2519.060 279.180 2519.320 279.440 ;
        RECT 680.440 16.700 680.700 16.960 ;
        RECT 682.740 16.700 683.000 16.960 ;
      LAYER met2 ;
        RECT 2519.050 886.875 2519.330 887.245 ;
        RECT 2519.120 279.470 2519.260 886.875 ;
        RECT 682.740 279.150 683.000 279.470 ;
        RECT 2519.060 279.150 2519.320 279.470 ;
        RECT 682.800 16.990 682.940 279.150 ;
        RECT 680.440 16.670 680.700 16.990 ;
        RECT 682.740 16.670 683.000 16.990 ;
        RECT 680.500 2.400 680.640 16.670 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 2519.050 886.920 2519.330 887.200 ;
      LAYER met3 ;
        RECT 2506.000 887.210 2510.000 887.360 ;
        RECT 2519.025 887.210 2519.355 887.225 ;
        RECT 2506.000 886.910 2519.355 887.210 ;
        RECT 2506.000 886.760 2510.000 886.910 ;
        RECT 2519.025 886.895 2519.355 886.910 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 155.280 1186.270 155.340 ;
        RECT 1559.470 155.280 1559.790 155.340 ;
        RECT 1185.950 155.140 1559.790 155.280 ;
        RECT 1185.950 155.080 1186.270 155.140 ;
        RECT 1559.470 155.080 1559.790 155.140 ;
        RECT 1179.970 18.260 1180.290 18.320 ;
        RECT 1185.950 18.260 1186.270 18.320 ;
        RECT 1179.970 18.120 1186.270 18.260 ;
        RECT 1179.970 18.060 1180.290 18.120 ;
        RECT 1185.950 18.060 1186.270 18.120 ;
      LAYER via ;
        RECT 1185.980 155.080 1186.240 155.340 ;
        RECT 1559.500 155.080 1559.760 155.340 ;
        RECT 1180.000 18.060 1180.260 18.320 ;
        RECT 1185.980 18.060 1186.240 18.320 ;
      LAYER met2 ;
        RECT 1561.010 510.410 1561.290 514.000 ;
        RECT 1559.560 510.270 1561.290 510.410 ;
        RECT 1559.560 155.370 1559.700 510.270 ;
        RECT 1561.010 510.000 1561.290 510.270 ;
        RECT 1185.980 155.050 1186.240 155.370 ;
        RECT 1559.500 155.050 1559.760 155.370 ;
        RECT 1186.040 18.350 1186.180 155.050 ;
        RECT 1180.000 18.030 1180.260 18.350 ;
        RECT 1185.980 18.030 1186.240 18.350 ;
        RECT 1180.060 2.400 1180.200 18.030 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 369.820 1200.530 369.880 ;
        RECT 1925.170 369.820 1925.490 369.880 ;
        RECT 1200.210 369.680 1925.490 369.820 ;
        RECT 1200.210 369.620 1200.530 369.680 ;
        RECT 1925.170 369.620 1925.490 369.680 ;
        RECT 1197.910 16.900 1198.230 16.960 ;
        RECT 1200.210 16.900 1200.530 16.960 ;
        RECT 1197.910 16.760 1200.530 16.900 ;
        RECT 1197.910 16.700 1198.230 16.760 ;
        RECT 1200.210 16.700 1200.530 16.760 ;
      LAYER via ;
        RECT 1200.240 369.620 1200.500 369.880 ;
        RECT 1925.200 369.620 1925.460 369.880 ;
        RECT 1197.940 16.700 1198.200 16.960 ;
        RECT 1200.240 16.700 1200.500 16.960 ;
      LAYER met2 ;
        RECT 1931.770 510.410 1932.050 514.000 ;
        RECT 1925.260 510.270 1932.050 510.410 ;
        RECT 1925.260 369.910 1925.400 510.270 ;
        RECT 1931.770 510.000 1932.050 510.270 ;
        RECT 1200.240 369.590 1200.500 369.910 ;
        RECT 1925.200 369.590 1925.460 369.910 ;
        RECT 1200.300 16.990 1200.440 369.590 ;
        RECT 1197.940 16.670 1198.200 16.990 ;
        RECT 1200.240 16.670 1200.500 16.990 ;
        RECT 1198.000 2.400 1198.140 16.670 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 383.080 427.730 383.140 ;
        RECT 1214.470 383.080 1214.790 383.140 ;
        RECT 427.410 382.940 1214.790 383.080 ;
        RECT 427.410 382.880 427.730 382.940 ;
        RECT 1214.470 382.880 1214.790 382.940 ;
      LAYER via ;
        RECT 427.440 382.880 427.700 383.140 ;
        RECT 1214.500 382.880 1214.760 383.140 ;
      LAYER met2 ;
        RECT 424.810 510.410 425.090 514.000 ;
        RECT 424.810 510.270 427.640 510.410 ;
        RECT 424.810 510.000 425.090 510.270 ;
        RECT 427.500 383.170 427.640 510.270 ;
        RECT 427.440 382.850 427.700 383.170 ;
        RECT 1214.500 382.850 1214.760 383.170 ;
        RECT 1214.560 3.130 1214.700 382.850 ;
        RECT 1214.560 2.990 1216.080 3.130 ;
        RECT 1215.940 2.400 1216.080 2.990 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 128.420 1235.030 128.480 ;
        RECT 2311.570 128.420 2311.890 128.480 ;
        RECT 1234.710 128.280 2311.890 128.420 ;
        RECT 1234.710 128.220 1235.030 128.280 ;
        RECT 2311.570 128.220 2311.890 128.280 ;
      LAYER via ;
        RECT 1234.740 128.220 1235.000 128.480 ;
        RECT 2311.600 128.220 2311.860 128.480 ;
      LAYER met2 ;
        RECT 2314.490 510.410 2314.770 514.000 ;
        RECT 2311.660 510.270 2314.770 510.410 ;
        RECT 2311.660 128.510 2311.800 510.270 ;
        RECT 2314.490 510.000 2314.770 510.270 ;
        RECT 1234.740 128.190 1235.000 128.510 ;
        RECT 2311.600 128.190 2311.860 128.510 ;
        RECT 1234.800 3.130 1234.940 128.190 ;
        RECT 1233.880 2.990 1234.940 3.130 ;
        RECT 1233.880 2.400 1234.020 2.990 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 494.260 1255.730 494.320 ;
        RECT 2519.950 494.260 2520.270 494.320 ;
        RECT 1255.410 494.120 2520.270 494.260 ;
        RECT 1255.410 494.060 1255.730 494.120 ;
        RECT 2519.950 494.060 2520.270 494.120 ;
        RECT 1251.730 16.900 1252.050 16.960 ;
        RECT 1255.410 16.900 1255.730 16.960 ;
        RECT 1251.730 16.760 1255.730 16.900 ;
        RECT 1251.730 16.700 1252.050 16.760 ;
        RECT 1255.410 16.700 1255.730 16.760 ;
      LAYER via ;
        RECT 1255.440 494.060 1255.700 494.320 ;
        RECT 2519.980 494.060 2520.240 494.320 ;
        RECT 1251.760 16.700 1252.020 16.960 ;
        RECT 1255.440 16.700 1255.700 16.960 ;
      LAYER met2 ;
        RECT 2519.970 594.475 2520.250 594.845 ;
        RECT 2520.040 494.350 2520.180 594.475 ;
        RECT 1255.440 494.030 1255.700 494.350 ;
        RECT 2519.980 494.030 2520.240 494.350 ;
        RECT 1255.500 16.990 1255.640 494.030 ;
        RECT 1251.760 16.670 1252.020 16.990 ;
        RECT 1255.440 16.670 1255.700 16.990 ;
        RECT 1251.820 2.400 1251.960 16.670 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
      LAYER via2 ;
        RECT 2519.970 594.520 2520.250 594.800 ;
      LAYER met3 ;
        RECT 2506.000 594.810 2510.000 594.960 ;
        RECT 2519.945 594.810 2520.275 594.825 ;
        RECT 2506.000 594.510 2520.275 594.810 ;
        RECT 2506.000 594.360 2510.000 594.510 ;
        RECT 2519.945 594.495 2520.275 594.510 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.550 3017.315 851.830 3017.685 ;
        RECT 851.620 3010.000 851.760 3017.315 ;
        RECT 851.620 3009.340 851.970 3010.000 ;
        RECT 851.690 3006.000 851.970 3009.340 ;
        RECT 334.970 2890.835 335.250 2891.205 ;
        RECT 335.040 2863.325 335.180 2890.835 ;
        RECT 334.970 2862.955 335.250 2863.325 ;
        RECT 334.970 2671.195 335.250 2671.565 ;
        RECT 335.040 2657.965 335.180 2671.195 ;
        RECT 334.970 2657.595 335.250 2657.965 ;
        RECT 332.670 2607.955 332.950 2608.325 ;
        RECT 332.740 2561.405 332.880 2607.955 ;
        RECT 332.670 2561.035 332.950 2561.405 ;
        RECT 333.130 2551.515 333.410 2551.885 ;
        RECT 333.200 2504.965 333.340 2551.515 ;
        RECT 333.130 2504.595 333.410 2504.965 ;
        RECT 334.970 2455.635 335.250 2456.005 ;
        RECT 335.040 2418.605 335.180 2455.635 ;
        RECT 334.970 2418.235 335.250 2418.605 ;
        RECT 334.970 2393.755 335.250 2394.125 ;
        RECT 335.040 2347.205 335.180 2393.755 ;
        RECT 334.970 2346.835 335.250 2347.205 ;
        RECT 334.510 2345.475 334.790 2345.845 ;
        RECT 334.580 2298.925 334.720 2345.475 ;
        RECT 334.510 2298.555 334.790 2298.925 ;
        RECT 333.590 2231.915 333.870 2232.285 ;
        RECT 333.660 2173.805 333.800 2231.915 ;
        RECT 333.590 2173.435 333.870 2173.805 ;
        RECT 334.510 1994.595 334.790 1994.965 ;
        RECT 334.580 1980.685 334.720 1994.595 ;
        RECT 334.510 1980.315 334.790 1980.685 ;
        RECT 334.970 1917.075 335.250 1917.445 ;
        RECT 335.040 1870.525 335.180 1917.075 ;
        RECT 334.970 1870.155 335.250 1870.525 ;
        RECT 333.590 1682.475 333.870 1682.845 ;
        RECT 333.660 1636.605 333.800 1682.475 ;
        RECT 333.590 1636.235 333.870 1636.605 ;
        RECT 334.970 1496.155 335.250 1496.525 ;
        RECT 335.040 1450.285 335.180 1496.155 ;
        RECT 334.970 1449.915 335.250 1450.285 ;
        RECT 334.510 1400.275 334.790 1400.645 ;
        RECT 334.580 1353.725 334.720 1400.275 ;
        RECT 334.510 1353.355 334.790 1353.725 ;
        RECT 335.430 1200.355 335.710 1200.725 ;
        RECT 335.500 1112.325 335.640 1200.355 ;
        RECT 335.430 1111.955 335.710 1112.325 ;
        RECT 333.590 1006.555 333.870 1006.925 ;
        RECT 333.660 977.685 333.800 1006.555 ;
        RECT 333.590 977.315 333.870 977.685 ;
        RECT 335.430 957.595 335.710 957.965 ;
        RECT 335.500 870.925 335.640 957.595 ;
        RECT 335.430 870.555 335.710 870.925 ;
        RECT 335.430 572.035 335.710 572.405 ;
        RECT 335.500 566.965 335.640 572.035 ;
        RECT 335.430 566.595 335.710 566.965 ;
        RECT 335.430 516.275 335.710 516.645 ;
        RECT 335.500 448.645 335.640 516.275 ;
        RECT 335.430 448.275 335.710 448.645 ;
        RECT 336.350 361.915 336.630 362.285 ;
        RECT 336.420 338.485 336.560 361.915 ;
        RECT 336.350 338.115 336.630 338.485 ;
        RECT 335.430 289.155 335.710 289.525 ;
        RECT 335.500 254.845 335.640 289.155 ;
        RECT 335.430 254.475 335.710 254.845 ;
        RECT 1268.770 46.395 1269.050 46.765 ;
        RECT 1268.840 17.410 1268.980 46.395 ;
        RECT 1268.840 17.270 1269.440 17.410 ;
        RECT 1269.300 2.400 1269.440 17.270 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 851.550 3017.360 851.830 3017.640 ;
        RECT 334.970 2890.880 335.250 2891.160 ;
        RECT 334.970 2863.000 335.250 2863.280 ;
        RECT 334.970 2671.240 335.250 2671.520 ;
        RECT 334.970 2657.640 335.250 2657.920 ;
        RECT 332.670 2608.000 332.950 2608.280 ;
        RECT 332.670 2561.080 332.950 2561.360 ;
        RECT 333.130 2551.560 333.410 2551.840 ;
        RECT 333.130 2504.640 333.410 2504.920 ;
        RECT 334.970 2455.680 335.250 2455.960 ;
        RECT 334.970 2418.280 335.250 2418.560 ;
        RECT 334.970 2393.800 335.250 2394.080 ;
        RECT 334.970 2346.880 335.250 2347.160 ;
        RECT 334.510 2345.520 334.790 2345.800 ;
        RECT 334.510 2298.600 334.790 2298.880 ;
        RECT 333.590 2231.960 333.870 2232.240 ;
        RECT 333.590 2173.480 333.870 2173.760 ;
        RECT 334.510 1994.640 334.790 1994.920 ;
        RECT 334.510 1980.360 334.790 1980.640 ;
        RECT 334.970 1917.120 335.250 1917.400 ;
        RECT 334.970 1870.200 335.250 1870.480 ;
        RECT 333.590 1682.520 333.870 1682.800 ;
        RECT 333.590 1636.280 333.870 1636.560 ;
        RECT 334.970 1496.200 335.250 1496.480 ;
        RECT 334.970 1449.960 335.250 1450.240 ;
        RECT 334.510 1400.320 334.790 1400.600 ;
        RECT 334.510 1353.400 334.790 1353.680 ;
        RECT 335.430 1200.400 335.710 1200.680 ;
        RECT 335.430 1112.000 335.710 1112.280 ;
        RECT 333.590 1006.600 333.870 1006.880 ;
        RECT 333.590 977.360 333.870 977.640 ;
        RECT 335.430 957.640 335.710 957.920 ;
        RECT 335.430 870.600 335.710 870.880 ;
        RECT 335.430 572.080 335.710 572.360 ;
        RECT 335.430 566.640 335.710 566.920 ;
        RECT 335.430 516.320 335.710 516.600 ;
        RECT 335.430 448.320 335.710 448.600 ;
        RECT 336.350 361.960 336.630 362.240 ;
        RECT 336.350 338.160 336.630 338.440 ;
        RECT 335.430 289.200 335.710 289.480 ;
        RECT 335.430 254.520 335.710 254.800 ;
        RECT 1268.770 46.440 1269.050 46.720 ;
      LAYER met3 ;
        RECT 448.310 3017.650 448.690 3017.660 ;
        RECT 851.525 3017.650 851.855 3017.665 ;
        RECT 448.310 3017.350 851.855 3017.650 ;
        RECT 448.310 3017.340 448.690 3017.350 ;
        RECT 851.525 3017.335 851.855 3017.350 ;
        RECT 404.150 3000.650 404.530 3000.660 ;
        RECT 448.310 3000.650 448.690 3000.660 ;
        RECT 404.150 3000.350 448.690 3000.650 ;
        RECT 404.150 3000.340 404.530 3000.350 ;
        RECT 448.310 3000.340 448.690 3000.350 ;
        RECT 334.230 2911.940 334.610 2912.260 ;
        RECT 334.270 2910.890 334.570 2911.940 ;
        RECT 335.150 2910.890 335.530 2910.900 ;
        RECT 334.270 2910.590 335.530 2910.890 ;
        RECT 335.150 2910.580 335.530 2910.590 ;
        RECT 334.945 2891.180 335.275 2891.185 ;
        RECT 334.945 2891.170 335.530 2891.180 ;
        RECT 334.720 2890.870 335.530 2891.170 ;
        RECT 334.945 2890.860 335.530 2890.870 ;
        RECT 334.945 2890.855 335.275 2890.860 ;
        RECT 334.945 2863.300 335.275 2863.305 ;
        RECT 334.945 2863.290 335.530 2863.300 ;
        RECT 334.945 2862.990 335.730 2863.290 ;
        RECT 334.945 2862.980 335.530 2862.990 ;
        RECT 334.945 2862.975 335.275 2862.980 ;
        RECT 334.230 2767.100 334.610 2767.420 ;
        RECT 334.270 2766.050 334.570 2767.100 ;
        RECT 335.150 2766.050 335.530 2766.060 ;
        RECT 334.270 2765.750 335.530 2766.050 ;
        RECT 335.150 2765.740 335.530 2765.750 ;
        RECT 335.150 2719.500 335.530 2719.820 ;
        RECT 335.190 2717.780 335.490 2719.500 ;
        RECT 335.150 2717.460 335.530 2717.780 ;
        RECT 334.945 2671.540 335.275 2671.545 ;
        RECT 334.945 2671.530 335.530 2671.540 ;
        RECT 334.720 2671.230 335.530 2671.530 ;
        RECT 334.945 2671.220 335.530 2671.230 ;
        RECT 334.945 2671.215 335.275 2671.220 ;
        RECT 334.945 2657.930 335.275 2657.945 ;
        RECT 334.945 2657.615 335.490 2657.930 ;
        RECT 335.190 2657.260 335.490 2657.615 ;
        RECT 335.150 2656.940 335.530 2657.260 ;
        RECT 335.150 2623.930 335.530 2623.940 ;
        RECT 333.350 2623.630 335.530 2623.930 ;
        RECT 333.350 2621.220 333.650 2623.630 ;
        RECT 335.150 2623.620 335.530 2623.630 ;
        RECT 333.310 2620.900 333.690 2621.220 ;
        RECT 332.645 2608.290 332.975 2608.305 ;
        RECT 333.310 2608.290 333.690 2608.300 ;
        RECT 332.645 2607.990 333.690 2608.290 ;
        RECT 332.645 2607.975 332.975 2607.990 ;
        RECT 333.310 2607.980 333.690 2607.990 ;
        RECT 332.645 2561.370 332.975 2561.385 ;
        RECT 332.430 2561.055 332.975 2561.370 ;
        RECT 332.430 2560.700 332.730 2561.055 ;
        RECT 332.390 2560.380 332.770 2560.700 ;
        RECT 332.390 2552.220 332.770 2552.540 ;
        RECT 332.430 2551.850 332.730 2552.220 ;
        RECT 333.105 2551.850 333.435 2551.865 ;
        RECT 332.430 2551.550 333.435 2551.850 ;
        RECT 333.105 2551.535 333.435 2551.550 ;
        RECT 333.105 2504.930 333.435 2504.945 ;
        RECT 335.150 2504.930 335.530 2504.940 ;
        RECT 333.105 2504.630 335.530 2504.930 ;
        RECT 333.105 2504.615 333.435 2504.630 ;
        RECT 335.150 2504.620 335.530 2504.630 ;
        RECT 334.945 2455.980 335.275 2455.985 ;
        RECT 334.945 2455.970 335.530 2455.980 ;
        RECT 334.720 2455.670 335.530 2455.970 ;
        RECT 334.945 2455.660 335.530 2455.670 ;
        RECT 334.945 2455.655 335.275 2455.660 ;
        RECT 334.945 2418.580 335.275 2418.585 ;
        RECT 334.945 2418.570 335.530 2418.580 ;
        RECT 334.720 2418.270 335.530 2418.570 ;
        RECT 334.945 2418.260 335.530 2418.270 ;
        RECT 334.945 2418.255 335.275 2418.260 ;
        RECT 334.945 2394.100 335.275 2394.105 ;
        RECT 334.945 2394.090 335.530 2394.100 ;
        RECT 334.720 2393.790 335.530 2394.090 ;
        RECT 334.945 2393.780 335.530 2393.790 ;
        RECT 334.945 2393.775 335.275 2393.780 ;
        RECT 334.945 2347.180 335.275 2347.185 ;
        RECT 334.945 2347.170 335.530 2347.180 ;
        RECT 334.945 2346.870 335.730 2347.170 ;
        RECT 334.945 2346.860 335.530 2346.870 ;
        RECT 334.945 2346.855 335.275 2346.860 ;
        RECT 334.485 2345.810 334.815 2345.825 ;
        RECT 335.150 2345.810 335.530 2345.820 ;
        RECT 334.485 2345.510 335.530 2345.810 ;
        RECT 334.485 2345.495 334.815 2345.510 ;
        RECT 335.150 2345.500 335.530 2345.510 ;
        RECT 334.485 2298.890 334.815 2298.905 ;
        RECT 334.270 2298.575 334.815 2298.890 ;
        RECT 334.270 2298.220 334.570 2298.575 ;
        RECT 334.230 2297.900 334.610 2298.220 ;
        RECT 333.565 2232.250 333.895 2232.265 ;
        RECT 335.150 2232.250 335.530 2232.260 ;
        RECT 333.565 2231.950 335.530 2232.250 ;
        RECT 333.565 2231.935 333.895 2231.950 ;
        RECT 335.150 2231.940 335.530 2231.950 ;
        RECT 333.565 2173.780 333.895 2173.785 ;
        RECT 333.310 2173.770 333.895 2173.780 ;
        RECT 333.110 2173.470 333.895 2173.770 ;
        RECT 333.310 2173.460 333.895 2173.470 ;
        RECT 333.565 2173.455 333.895 2173.460 ;
        RECT 334.485 1994.930 334.815 1994.945 ;
        RECT 336.070 1994.930 336.450 1994.940 ;
        RECT 334.485 1994.630 336.450 1994.930 ;
        RECT 334.485 1994.615 334.815 1994.630 ;
        RECT 336.070 1994.620 336.450 1994.630 ;
        RECT 334.485 1980.660 334.815 1980.665 ;
        RECT 334.230 1980.650 334.815 1980.660 ;
        RECT 334.030 1980.350 334.815 1980.650 ;
        RECT 334.230 1980.340 334.815 1980.350 ;
        RECT 334.485 1980.335 334.815 1980.340 ;
        RECT 334.230 1972.860 334.610 1973.180 ;
        RECT 334.270 1972.490 334.570 1972.860 ;
        RECT 335.150 1972.490 335.530 1972.500 ;
        RECT 334.270 1972.190 335.530 1972.490 ;
        RECT 335.150 1972.180 335.530 1972.190 ;
        RECT 335.150 1917.780 335.530 1918.100 ;
        RECT 335.190 1917.425 335.490 1917.780 ;
        RECT 334.945 1917.110 335.490 1917.425 ;
        RECT 334.945 1917.095 335.275 1917.110 ;
        RECT 334.945 1870.490 335.275 1870.505 ;
        RECT 336.070 1870.490 336.450 1870.500 ;
        RECT 334.945 1870.190 336.450 1870.490 ;
        RECT 334.945 1870.175 335.275 1870.190 ;
        RECT 336.070 1870.180 336.450 1870.190 ;
        RECT 334.230 1869.130 334.610 1869.140 ;
        RECT 336.070 1869.130 336.450 1869.140 ;
        RECT 334.230 1868.830 336.450 1869.130 ;
        RECT 334.230 1868.820 334.610 1868.830 ;
        RECT 336.070 1868.820 336.450 1868.830 ;
        RECT 336.070 1753.530 336.450 1753.540 ;
        RECT 334.270 1753.230 336.450 1753.530 ;
        RECT 334.270 1752.860 334.570 1753.230 ;
        RECT 336.070 1753.220 336.450 1753.230 ;
        RECT 334.230 1752.540 334.610 1752.860 ;
        RECT 334.230 1704.940 334.610 1705.260 ;
        RECT 334.270 1703.890 334.570 1704.940 ;
        RECT 335.150 1703.890 335.530 1703.900 ;
        RECT 334.270 1703.590 335.530 1703.890 ;
        RECT 335.150 1703.580 335.530 1703.590 ;
        RECT 335.150 1683.180 335.530 1683.500 ;
        RECT 333.565 1682.810 333.895 1682.825 ;
        RECT 335.190 1682.810 335.490 1683.180 ;
        RECT 333.565 1682.510 335.490 1682.810 ;
        RECT 333.565 1682.495 333.895 1682.510 ;
        RECT 333.565 1636.570 333.895 1636.585 ;
        RECT 333.350 1636.255 333.895 1636.570 ;
        RECT 333.350 1635.900 333.650 1636.255 ;
        RECT 333.310 1635.580 333.690 1635.900 ;
        RECT 335.150 1560.410 335.530 1560.420 ;
        RECT 334.270 1560.110 335.530 1560.410 ;
        RECT 334.270 1559.060 334.570 1560.110 ;
        RECT 335.150 1560.100 335.530 1560.110 ;
        RECT 334.230 1558.740 334.610 1559.060 ;
        RECT 333.310 1511.140 333.690 1511.460 ;
        RECT 333.350 1510.770 333.650 1511.140 ;
        RECT 334.230 1510.770 334.610 1510.780 ;
        RECT 333.350 1510.470 334.610 1510.770 ;
        RECT 334.230 1510.460 334.610 1510.470 ;
        RECT 335.150 1496.860 335.530 1497.180 ;
        RECT 335.190 1496.505 335.490 1496.860 ;
        RECT 334.945 1496.190 335.490 1496.505 ;
        RECT 334.945 1496.175 335.275 1496.190 ;
        RECT 334.945 1450.250 335.275 1450.265 ;
        RECT 334.945 1449.935 335.490 1450.250 ;
        RECT 335.190 1449.580 335.490 1449.935 ;
        RECT 335.150 1449.260 335.530 1449.580 ;
        RECT 334.485 1400.610 334.815 1400.625 ;
        RECT 335.150 1400.610 335.530 1400.620 ;
        RECT 334.485 1400.310 335.530 1400.610 ;
        RECT 334.485 1400.295 334.815 1400.310 ;
        RECT 335.150 1400.300 335.530 1400.310 ;
        RECT 334.485 1353.690 334.815 1353.705 ;
        RECT 334.270 1353.375 334.815 1353.690 ;
        RECT 334.270 1353.020 334.570 1353.375 ;
        RECT 334.230 1352.700 334.610 1353.020 ;
        RECT 333.310 1304.050 333.690 1304.060 ;
        RECT 335.150 1304.050 335.530 1304.060 ;
        RECT 333.310 1303.750 335.530 1304.050 ;
        RECT 333.310 1303.740 333.690 1303.750 ;
        RECT 335.150 1303.740 335.530 1303.750 ;
        RECT 336.070 1255.460 336.450 1255.780 ;
        RECT 335.150 1255.090 335.530 1255.100 ;
        RECT 336.110 1255.090 336.410 1255.460 ;
        RECT 335.150 1254.790 336.410 1255.090 ;
        RECT 335.150 1254.780 335.530 1254.790 ;
        RECT 335.405 1200.690 335.735 1200.705 ;
        RECT 336.070 1200.690 336.450 1200.700 ;
        RECT 335.405 1200.390 336.450 1200.690 ;
        RECT 335.405 1200.375 335.735 1200.390 ;
        RECT 336.070 1200.380 336.450 1200.390 ;
        RECT 335.405 1112.290 335.735 1112.305 ;
        RECT 335.190 1111.975 335.735 1112.290 ;
        RECT 335.190 1111.620 335.490 1111.975 ;
        RECT 335.150 1111.300 335.530 1111.620 ;
        RECT 335.150 1077.610 335.530 1077.620 ;
        RECT 334.270 1077.310 335.530 1077.610 ;
        RECT 334.270 1076.260 334.570 1077.310 ;
        RECT 335.150 1077.300 335.530 1077.310 ;
        RECT 334.230 1075.940 334.610 1076.260 ;
        RECT 333.565 1006.900 333.895 1006.905 ;
        RECT 333.310 1006.890 333.895 1006.900 ;
        RECT 333.310 1006.590 334.120 1006.890 ;
        RECT 333.310 1006.580 333.895 1006.590 ;
        RECT 333.565 1006.575 333.895 1006.580 ;
        RECT 332.390 977.650 332.770 977.660 ;
        RECT 333.565 977.650 333.895 977.665 ;
        RECT 332.390 977.350 333.895 977.650 ;
        RECT 332.390 977.340 332.770 977.350 ;
        RECT 333.565 977.335 333.895 977.350 ;
        RECT 332.390 958.300 332.770 958.620 ;
        RECT 332.430 957.930 332.730 958.300 ;
        RECT 335.405 957.930 335.735 957.945 ;
        RECT 332.430 957.630 335.735 957.930 ;
        RECT 335.405 957.615 335.735 957.630 ;
        RECT 335.405 870.890 335.735 870.905 ;
        RECT 335.405 870.590 336.410 870.890 ;
        RECT 335.405 870.575 335.735 870.590 ;
        RECT 336.110 870.220 336.410 870.590 ;
        RECT 336.070 869.900 336.450 870.220 ;
        RECT 333.310 724.690 333.690 724.700 ;
        RECT 334.230 724.690 334.610 724.700 ;
        RECT 333.310 724.390 334.610 724.690 ;
        RECT 333.310 724.380 333.690 724.390 ;
        RECT 334.230 724.380 334.610 724.390 ;
        RECT 333.310 689.330 333.690 689.340 ;
        RECT 336.070 689.330 336.450 689.340 ;
        RECT 333.310 689.030 336.450 689.330 ;
        RECT 333.310 689.020 333.690 689.030 ;
        RECT 336.070 689.020 336.450 689.030 ;
        RECT 335.405 572.380 335.735 572.385 ;
        RECT 335.150 572.370 335.735 572.380 ;
        RECT 335.150 572.070 335.960 572.370 ;
        RECT 335.150 572.060 335.735 572.070 ;
        RECT 335.405 572.055 335.735 572.060 ;
        RECT 335.405 566.930 335.735 566.945 ;
        RECT 335.190 566.615 335.735 566.930 ;
        RECT 335.190 566.260 335.490 566.615 ;
        RECT 335.150 565.940 335.530 566.260 ;
        RECT 335.150 516.980 335.530 517.300 ;
        RECT 335.190 516.625 335.490 516.980 ;
        RECT 335.190 516.310 335.735 516.625 ;
        RECT 335.405 516.295 335.735 516.310 ;
        RECT 335.405 448.620 335.735 448.625 ;
        RECT 335.150 448.610 335.735 448.620 ;
        RECT 334.950 448.310 335.735 448.610 ;
        RECT 335.150 448.300 335.735 448.310 ;
        RECT 335.405 448.295 335.735 448.300 ;
        RECT 336.325 362.260 336.655 362.265 ;
        RECT 336.070 362.250 336.655 362.260 ;
        RECT 336.070 361.950 336.880 362.250 ;
        RECT 336.070 361.940 336.655 361.950 ;
        RECT 336.325 361.935 336.655 361.940 ;
        RECT 336.325 338.460 336.655 338.465 ;
        RECT 336.070 338.450 336.655 338.460 ;
        RECT 335.870 338.150 336.655 338.450 ;
        RECT 336.070 338.140 336.655 338.150 ;
        RECT 336.325 338.135 336.655 338.140 ;
        RECT 336.070 304.450 336.450 304.460 ;
        RECT 335.190 304.150 336.450 304.450 ;
        RECT 335.190 303.100 335.490 304.150 ;
        RECT 336.070 304.140 336.450 304.150 ;
        RECT 335.150 302.780 335.530 303.100 ;
        RECT 335.405 289.500 335.735 289.505 ;
        RECT 335.150 289.490 335.735 289.500 ;
        RECT 335.150 289.190 335.960 289.490 ;
        RECT 335.150 289.180 335.735 289.190 ;
        RECT 335.405 289.175 335.735 289.180 ;
        RECT 335.405 254.820 335.735 254.825 ;
        RECT 335.150 254.810 335.735 254.820 ;
        RECT 334.950 254.510 335.735 254.810 ;
        RECT 335.150 254.500 335.735 254.510 ;
        RECT 335.405 254.495 335.735 254.500 ;
        RECT 333.310 46.730 333.690 46.740 ;
        RECT 1268.745 46.730 1269.075 46.745 ;
        RECT 333.310 46.430 1269.075 46.730 ;
        RECT 333.310 46.420 333.690 46.430 ;
        RECT 1268.745 46.415 1269.075 46.430 ;
      LAYER via3 ;
        RECT 448.340 3017.340 448.660 3017.660 ;
        RECT 404.180 3000.340 404.500 3000.660 ;
        RECT 448.340 3000.340 448.660 3000.660 ;
        RECT 334.260 2911.940 334.580 2912.260 ;
        RECT 335.180 2910.580 335.500 2910.900 ;
        RECT 335.180 2890.860 335.500 2891.180 ;
        RECT 335.180 2862.980 335.500 2863.300 ;
        RECT 334.260 2767.100 334.580 2767.420 ;
        RECT 335.180 2765.740 335.500 2766.060 ;
        RECT 335.180 2719.500 335.500 2719.820 ;
        RECT 335.180 2717.460 335.500 2717.780 ;
        RECT 335.180 2671.220 335.500 2671.540 ;
        RECT 335.180 2656.940 335.500 2657.260 ;
        RECT 335.180 2623.620 335.500 2623.940 ;
        RECT 333.340 2620.900 333.660 2621.220 ;
        RECT 333.340 2607.980 333.660 2608.300 ;
        RECT 332.420 2560.380 332.740 2560.700 ;
        RECT 332.420 2552.220 332.740 2552.540 ;
        RECT 335.180 2504.620 335.500 2504.940 ;
        RECT 335.180 2455.660 335.500 2455.980 ;
        RECT 335.180 2418.260 335.500 2418.580 ;
        RECT 335.180 2393.780 335.500 2394.100 ;
        RECT 335.180 2346.860 335.500 2347.180 ;
        RECT 335.180 2345.500 335.500 2345.820 ;
        RECT 334.260 2297.900 334.580 2298.220 ;
        RECT 335.180 2231.940 335.500 2232.260 ;
        RECT 333.340 2173.460 333.660 2173.780 ;
        RECT 336.100 1994.620 336.420 1994.940 ;
        RECT 334.260 1980.340 334.580 1980.660 ;
        RECT 334.260 1972.860 334.580 1973.180 ;
        RECT 335.180 1972.180 335.500 1972.500 ;
        RECT 335.180 1917.780 335.500 1918.100 ;
        RECT 336.100 1870.180 336.420 1870.500 ;
        RECT 334.260 1868.820 334.580 1869.140 ;
        RECT 336.100 1868.820 336.420 1869.140 ;
        RECT 336.100 1753.220 336.420 1753.540 ;
        RECT 334.260 1752.540 334.580 1752.860 ;
        RECT 334.260 1704.940 334.580 1705.260 ;
        RECT 335.180 1703.580 335.500 1703.900 ;
        RECT 335.180 1683.180 335.500 1683.500 ;
        RECT 333.340 1635.580 333.660 1635.900 ;
        RECT 335.180 1560.100 335.500 1560.420 ;
        RECT 334.260 1558.740 334.580 1559.060 ;
        RECT 333.340 1511.140 333.660 1511.460 ;
        RECT 334.260 1510.460 334.580 1510.780 ;
        RECT 335.180 1496.860 335.500 1497.180 ;
        RECT 335.180 1449.260 335.500 1449.580 ;
        RECT 335.180 1400.300 335.500 1400.620 ;
        RECT 334.260 1352.700 334.580 1353.020 ;
        RECT 333.340 1303.740 333.660 1304.060 ;
        RECT 335.180 1303.740 335.500 1304.060 ;
        RECT 336.100 1255.460 336.420 1255.780 ;
        RECT 335.180 1254.780 335.500 1255.100 ;
        RECT 336.100 1200.380 336.420 1200.700 ;
        RECT 335.180 1111.300 335.500 1111.620 ;
        RECT 335.180 1077.300 335.500 1077.620 ;
        RECT 334.260 1075.940 334.580 1076.260 ;
        RECT 333.340 1006.580 333.660 1006.900 ;
        RECT 332.420 977.340 332.740 977.660 ;
        RECT 332.420 958.300 332.740 958.620 ;
        RECT 336.100 869.900 336.420 870.220 ;
        RECT 333.340 724.380 333.660 724.700 ;
        RECT 334.260 724.380 334.580 724.700 ;
        RECT 333.340 689.020 333.660 689.340 ;
        RECT 336.100 689.020 336.420 689.340 ;
        RECT 335.180 572.060 335.500 572.380 ;
        RECT 335.180 565.940 335.500 566.260 ;
        RECT 335.180 516.980 335.500 517.300 ;
        RECT 335.180 448.300 335.500 448.620 ;
        RECT 336.100 361.940 336.420 362.260 ;
        RECT 336.100 338.140 336.420 338.460 ;
        RECT 336.100 304.140 336.420 304.460 ;
        RECT 335.180 302.780 335.500 303.100 ;
        RECT 335.180 289.180 335.500 289.500 ;
        RECT 335.180 254.500 335.500 254.820 ;
        RECT 333.340 46.420 333.660 46.740 ;
      LAYER met4 ;
        RECT 448.335 3017.335 448.665 3017.665 ;
        RECT 448.350 3000.665 448.650 3017.335 ;
        RECT 404.175 3000.335 404.505 3000.665 ;
        RECT 448.335 3000.335 448.665 3000.665 ;
        RECT 404.190 2994.290 404.490 3000.335 ;
        RECT 333.830 2993.850 335.010 2994.290 ;
        RECT 333.830 2993.550 336.410 2993.850 ;
        RECT 333.830 2993.110 335.010 2993.550 ;
        RECT 336.110 2959.850 336.410 2993.550 ;
        RECT 403.750 2993.110 404.930 2994.290 ;
        RECT 334.270 2959.550 336.410 2959.850 ;
        RECT 334.270 2912.265 334.570 2959.550 ;
        RECT 334.255 2911.935 334.585 2912.265 ;
        RECT 335.175 2910.575 335.505 2910.905 ;
        RECT 335.190 2891.185 335.490 2910.575 ;
        RECT 335.175 2890.855 335.505 2891.185 ;
        RECT 335.175 2862.975 335.505 2863.305 ;
        RECT 335.190 2813.650 335.490 2862.975 ;
        RECT 334.270 2813.350 335.490 2813.650 ;
        RECT 334.270 2767.425 334.570 2813.350 ;
        RECT 334.255 2767.095 334.585 2767.425 ;
        RECT 335.175 2765.735 335.505 2766.065 ;
        RECT 335.190 2719.825 335.490 2765.735 ;
        RECT 335.175 2719.495 335.505 2719.825 ;
        RECT 335.175 2717.455 335.505 2717.785 ;
        RECT 335.190 2671.545 335.490 2717.455 ;
        RECT 335.175 2671.215 335.505 2671.545 ;
        RECT 335.175 2656.935 335.505 2657.265 ;
        RECT 335.190 2623.945 335.490 2656.935 ;
        RECT 335.175 2623.615 335.505 2623.945 ;
        RECT 333.335 2620.895 333.665 2621.225 ;
        RECT 333.350 2608.305 333.650 2620.895 ;
        RECT 333.335 2607.975 333.665 2608.305 ;
        RECT 332.415 2560.375 332.745 2560.705 ;
        RECT 332.430 2552.545 332.730 2560.375 ;
        RECT 332.415 2552.215 332.745 2552.545 ;
        RECT 335.175 2504.615 335.505 2504.945 ;
        RECT 335.190 2455.985 335.490 2504.615 ;
        RECT 335.175 2455.655 335.505 2455.985 ;
        RECT 335.175 2418.255 335.505 2418.585 ;
        RECT 335.190 2394.105 335.490 2418.255 ;
        RECT 335.175 2393.775 335.505 2394.105 ;
        RECT 335.175 2346.855 335.505 2347.185 ;
        RECT 335.190 2345.825 335.490 2346.855 ;
        RECT 335.175 2345.495 335.505 2345.825 ;
        RECT 334.255 2297.895 334.585 2298.225 ;
        RECT 334.270 2279.850 334.570 2297.895 ;
        RECT 334.270 2279.550 335.490 2279.850 ;
        RECT 335.190 2232.265 335.490 2279.550 ;
        RECT 335.175 2231.935 335.505 2232.265 ;
        RECT 333.335 2173.455 333.665 2173.785 ;
        RECT 333.350 2133.650 333.650 2173.455 ;
        RECT 333.350 2133.350 336.410 2133.650 ;
        RECT 336.110 1994.945 336.410 2133.350 ;
        RECT 336.095 1994.615 336.425 1994.945 ;
        RECT 334.255 1980.335 334.585 1980.665 ;
        RECT 334.270 1973.185 334.570 1980.335 ;
        RECT 334.255 1972.855 334.585 1973.185 ;
        RECT 335.175 1972.175 335.505 1972.505 ;
        RECT 335.190 1918.105 335.490 1972.175 ;
        RECT 335.175 1917.775 335.505 1918.105 ;
        RECT 336.095 1870.175 336.425 1870.505 ;
        RECT 336.110 1869.145 336.410 1870.175 ;
        RECT 334.255 1868.815 334.585 1869.145 ;
        RECT 336.095 1868.815 336.425 1869.145 ;
        RECT 334.270 1844.650 334.570 1868.815 ;
        RECT 334.270 1844.350 336.410 1844.650 ;
        RECT 336.110 1753.545 336.410 1844.350 ;
        RECT 336.095 1753.215 336.425 1753.545 ;
        RECT 334.255 1752.535 334.585 1752.865 ;
        RECT 334.270 1705.265 334.570 1752.535 ;
        RECT 334.255 1704.935 334.585 1705.265 ;
        RECT 335.175 1703.575 335.505 1703.905 ;
        RECT 335.190 1683.505 335.490 1703.575 ;
        RECT 335.175 1683.175 335.505 1683.505 ;
        RECT 333.335 1635.575 333.665 1635.905 ;
        RECT 333.350 1606.650 333.650 1635.575 ;
        RECT 333.350 1606.350 335.490 1606.650 ;
        RECT 335.190 1560.425 335.490 1606.350 ;
        RECT 335.175 1560.095 335.505 1560.425 ;
        RECT 334.255 1558.735 334.585 1559.065 ;
        RECT 334.270 1545.450 334.570 1558.735 ;
        RECT 333.350 1545.150 334.570 1545.450 ;
        RECT 333.350 1511.465 333.650 1545.150 ;
        RECT 333.335 1511.135 333.665 1511.465 ;
        RECT 334.255 1510.455 334.585 1510.785 ;
        RECT 334.270 1501.250 334.570 1510.455 ;
        RECT 334.270 1500.950 335.260 1501.250 ;
        RECT 334.960 1497.850 335.260 1500.950 ;
        RECT 334.960 1497.550 335.490 1497.850 ;
        RECT 335.190 1497.185 335.490 1497.550 ;
        RECT 335.175 1496.855 335.505 1497.185 ;
        RECT 335.175 1449.255 335.505 1449.585 ;
        RECT 335.190 1400.625 335.490 1449.255 ;
        RECT 335.175 1400.295 335.505 1400.625 ;
        RECT 334.255 1352.695 334.585 1353.025 ;
        RECT 334.270 1321.050 334.570 1352.695 ;
        RECT 332.430 1320.750 334.570 1321.050 ;
        RECT 332.430 1317.650 332.730 1320.750 ;
        RECT 332.430 1317.350 333.650 1317.650 ;
        RECT 333.350 1304.065 333.650 1317.350 ;
        RECT 333.335 1303.735 333.665 1304.065 ;
        RECT 335.175 1303.735 335.505 1304.065 ;
        RECT 335.190 1263.250 335.490 1303.735 ;
        RECT 335.190 1262.950 336.410 1263.250 ;
        RECT 336.110 1255.785 336.410 1262.950 ;
        RECT 336.095 1255.455 336.425 1255.785 ;
        RECT 335.175 1254.775 335.505 1255.105 ;
        RECT 335.190 1208.850 335.490 1254.775 ;
        RECT 335.190 1208.550 336.410 1208.850 ;
        RECT 336.110 1200.705 336.410 1208.550 ;
        RECT 336.095 1200.375 336.425 1200.705 ;
        RECT 335.175 1111.295 335.505 1111.625 ;
        RECT 335.190 1077.625 335.490 1111.295 ;
        RECT 335.175 1077.295 335.505 1077.625 ;
        RECT 334.255 1075.935 334.585 1076.265 ;
        RECT 334.270 1028.650 334.570 1075.935 ;
        RECT 333.350 1028.350 334.570 1028.650 ;
        RECT 333.350 1006.905 333.650 1028.350 ;
        RECT 333.335 1006.575 333.665 1006.905 ;
        RECT 332.415 977.335 332.745 977.665 ;
        RECT 332.430 958.625 332.730 977.335 ;
        RECT 332.415 958.295 332.745 958.625 ;
        RECT 336.095 869.895 336.425 870.225 ;
        RECT 336.110 834.850 336.410 869.895 ;
        RECT 335.190 834.550 336.410 834.850 ;
        RECT 335.190 787.250 335.490 834.550 ;
        RECT 334.270 786.950 335.490 787.250 ;
        RECT 334.270 724.705 334.570 786.950 ;
        RECT 333.335 724.375 333.665 724.705 ;
        RECT 334.255 724.375 334.585 724.705 ;
        RECT 333.350 689.345 333.650 724.375 ;
        RECT 333.335 689.015 333.665 689.345 ;
        RECT 336.095 689.015 336.425 689.345 ;
        RECT 336.110 641.050 336.410 689.015 ;
        RECT 335.190 640.750 336.410 641.050 ;
        RECT 335.190 572.385 335.490 640.750 ;
        RECT 335.175 572.055 335.505 572.385 ;
        RECT 335.175 565.935 335.505 566.265 ;
        RECT 335.190 517.305 335.490 565.935 ;
        RECT 335.175 516.975 335.505 517.305 ;
        RECT 335.175 448.295 335.505 448.625 ;
        RECT 335.190 389.450 335.490 448.295 ;
        RECT 335.190 389.150 336.410 389.450 ;
        RECT 336.110 362.265 336.410 389.150 ;
        RECT 336.095 361.935 336.425 362.265 ;
        RECT 336.095 338.135 336.425 338.465 ;
        RECT 336.110 304.465 336.410 338.135 ;
        RECT 336.095 304.135 336.425 304.465 ;
        RECT 335.175 302.775 335.505 303.105 ;
        RECT 335.190 289.505 335.490 302.775 ;
        RECT 335.175 289.175 335.505 289.505 ;
        RECT 335.175 254.495 335.505 254.825 ;
        RECT 335.190 205.850 335.490 254.495 ;
        RECT 334.270 205.550 335.490 205.850 ;
        RECT 334.270 161.650 334.570 205.550 ;
        RECT 332.430 161.350 334.570 161.650 ;
        RECT 332.430 158.250 332.730 161.350 ;
        RECT 332.430 157.950 333.650 158.250 ;
        RECT 333.350 110.650 333.650 157.950 ;
        RECT 333.350 110.350 334.570 110.650 ;
        RECT 334.270 63.050 334.570 110.350 ;
        RECT 333.350 62.750 334.570 63.050 ;
        RECT 333.350 46.745 333.650 62.750 ;
        RECT 333.335 46.415 333.665 46.745 ;
      LAYER met5 ;
        RECT 333.620 2992.900 405.140 2994.500 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 3010.940 372.530 3011.000 ;
        RECT 678.570 3010.940 678.890 3011.000 ;
        RECT 372.210 3010.800 678.890 3010.940 ;
        RECT 372.210 3010.740 372.530 3010.800 ;
        RECT 678.570 3010.740 678.890 3010.800 ;
        RECT 1287.150 19.280 1287.470 19.340 ;
        RECT 1256.880 19.140 1287.470 19.280 ;
        RECT 372.210 18.600 372.530 18.660 ;
        RECT 1256.880 18.600 1257.020 19.140 ;
        RECT 1287.150 19.080 1287.470 19.140 ;
        RECT 372.210 18.460 1257.020 18.600 ;
        RECT 372.210 18.400 372.530 18.460 ;
      LAYER via ;
        RECT 372.240 3010.740 372.500 3011.000 ;
        RECT 678.600 3010.740 678.860 3011.000 ;
        RECT 372.240 18.400 372.500 18.660 ;
        RECT 1287.180 19.080 1287.440 19.340 ;
      LAYER met2 ;
        RECT 372.240 3010.710 372.500 3011.030 ;
        RECT 678.600 3010.710 678.860 3011.030 ;
        RECT 372.300 18.690 372.440 3010.710 ;
        RECT 678.660 3010.000 678.800 3010.710 ;
        RECT 678.660 3009.340 679.010 3010.000 ;
        RECT 678.730 3006.000 679.010 3009.340 ;
        RECT 1287.180 19.050 1287.440 19.370 ;
        RECT 372.240 18.370 372.500 18.690 ;
        RECT 1287.240 2.400 1287.380 19.050 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 455.545 3001.945 455.715 3006.535 ;
      LAYER mcon ;
        RECT 455.545 3006.365 455.715 3006.535 ;
      LAYER met1 ;
        RECT 455.470 3006.520 455.790 3006.580 ;
        RECT 455.275 3006.380 455.790 3006.520 ;
        RECT 455.470 3006.320 455.790 3006.380 ;
        RECT 309.650 3002.100 309.970 3002.160 ;
        RECT 455.485 3002.100 455.775 3002.145 ;
        RECT 309.650 3001.960 455.775 3002.100 ;
        RECT 309.650 3001.900 309.970 3001.960 ;
        RECT 455.485 3001.915 455.775 3001.960 ;
        RECT 309.650 61.440 309.970 61.500 ;
        RECT 1304.170 61.440 1304.490 61.500 ;
        RECT 309.650 61.300 1304.490 61.440 ;
        RECT 309.650 61.240 309.970 61.300 ;
        RECT 1304.170 61.240 1304.490 61.300 ;
      LAYER via ;
        RECT 455.500 3006.320 455.760 3006.580 ;
        RECT 309.680 3001.900 309.940 3002.160 ;
        RECT 309.680 61.240 309.940 61.500 ;
        RECT 1304.200 61.240 1304.460 61.500 ;
      LAYER met2 ;
        RECT 456.090 3006.690 456.370 3010.000 ;
        RECT 455.560 3006.610 456.370 3006.690 ;
        RECT 455.500 3006.550 456.370 3006.610 ;
        RECT 455.500 3006.290 455.760 3006.550 ;
        RECT 456.090 3006.000 456.370 3006.550 ;
        RECT 309.680 3001.870 309.940 3002.190 ;
        RECT 309.740 61.530 309.880 3001.870 ;
        RECT 309.680 61.210 309.940 61.530 ;
        RECT 1304.200 61.210 1304.460 61.530 ;
        RECT 1304.260 17.410 1304.400 61.210 ;
        RECT 1304.260 17.270 1305.320 17.410 ;
        RECT 1305.180 2.400 1305.320 17.270 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 376.810 2284.020 377.130 2284.080 ;
        RECT 393.370 2284.020 393.690 2284.080 ;
        RECT 376.810 2283.880 393.690 2284.020 ;
        RECT 376.810 2283.820 377.130 2283.880 ;
        RECT 393.370 2283.820 393.690 2283.880 ;
        RECT 376.810 390.560 377.130 390.620 ;
        RECT 1317.970 390.560 1318.290 390.620 ;
        RECT 376.810 390.420 1318.290 390.560 ;
        RECT 376.810 390.360 377.130 390.420 ;
        RECT 1317.970 390.360 1318.290 390.420 ;
      LAYER via ;
        RECT 376.840 2283.820 377.100 2284.080 ;
        RECT 393.400 2283.820 393.660 2284.080 ;
        RECT 376.840 390.360 377.100 390.620 ;
        RECT 1318.000 390.360 1318.260 390.620 ;
      LAYER met2 ;
        RECT 393.390 2284.955 393.670 2285.325 ;
        RECT 393.460 2284.110 393.600 2284.955 ;
        RECT 376.840 2283.790 377.100 2284.110 ;
        RECT 393.400 2283.790 393.660 2284.110 ;
        RECT 376.900 390.650 377.040 2283.790 ;
        RECT 376.840 390.330 377.100 390.650 ;
        RECT 1318.000 390.330 1318.260 390.650 ;
        RECT 1318.060 17.410 1318.200 390.330 ;
        RECT 1318.060 17.270 1323.260 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
      LAYER via2 ;
        RECT 393.390 2285.000 393.670 2285.280 ;
      LAYER met3 ;
        RECT 393.365 2285.290 393.695 2285.305 ;
        RECT 410.000 2285.290 414.000 2285.440 ;
        RECT 393.365 2284.990 414.000 2285.290 ;
        RECT 393.365 2284.975 393.695 2284.990 ;
        RECT 410.000 2284.840 414.000 2284.990 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 376.350 1787.280 376.670 1787.340 ;
        RECT 393.370 1787.280 393.690 1787.340 ;
        RECT 376.350 1787.140 393.690 1787.280 ;
        RECT 376.350 1787.080 376.670 1787.140 ;
        RECT 393.370 1787.080 393.690 1787.140 ;
        RECT 376.350 307.940 376.670 308.000 ;
        RECT 1338.670 307.940 1338.990 308.000 ;
        RECT 376.350 307.800 1338.990 307.940 ;
        RECT 376.350 307.740 376.670 307.800 ;
        RECT 1338.670 307.740 1338.990 307.800 ;
      LAYER via ;
        RECT 376.380 1787.080 376.640 1787.340 ;
        RECT 393.400 1787.080 393.660 1787.340 ;
        RECT 376.380 307.740 376.640 308.000 ;
        RECT 1338.700 307.740 1338.960 308.000 ;
      LAYER met2 ;
        RECT 393.390 1791.275 393.670 1791.645 ;
        RECT 393.460 1787.370 393.600 1791.275 ;
        RECT 376.380 1787.050 376.640 1787.370 ;
        RECT 393.400 1787.050 393.660 1787.370 ;
        RECT 376.440 308.030 376.580 1787.050 ;
        RECT 376.380 307.710 376.640 308.030 ;
        RECT 1338.700 307.710 1338.960 308.030 ;
        RECT 1338.760 17.410 1338.900 307.710 ;
        RECT 1338.760 17.270 1340.740 17.410 ;
        RECT 1340.600 2.400 1340.740 17.270 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
      LAYER via2 ;
        RECT 393.390 1791.320 393.670 1791.600 ;
      LAYER met3 ;
        RECT 393.365 1791.610 393.695 1791.625 ;
        RECT 410.000 1791.610 414.000 1791.760 ;
        RECT 393.365 1791.310 414.000 1791.610 ;
        RECT 393.365 1791.295 393.695 1791.310 ;
        RECT 410.000 1791.160 414.000 1791.310 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 14.520 698.670 14.580 ;
        RECT 703.410 14.520 703.730 14.580 ;
        RECT 698.350 14.380 703.730 14.520 ;
        RECT 698.350 14.320 698.670 14.380 ;
        RECT 703.410 14.320 703.730 14.380 ;
      LAYER via ;
        RECT 698.380 14.320 698.640 14.580 ;
        RECT 703.440 14.320 703.700 14.580 ;
      LAYER met2 ;
        RECT 703.430 223.875 703.710 224.245 ;
        RECT 703.500 14.610 703.640 223.875 ;
        RECT 698.380 14.290 698.640 14.610 ;
        RECT 703.440 14.290 703.700 14.610 ;
        RECT 698.440 2.400 698.580 14.290 ;
        RECT 698.230 -4.800 698.790 2.400 ;
      LAYER via2 ;
        RECT 703.430 223.920 703.710 224.200 ;
      LAYER met3 ;
        RECT 2506.000 2274.410 2510.000 2274.560 ;
        RECT 2533.950 2274.410 2534.330 2274.420 ;
        RECT 2506.000 2274.110 2534.330 2274.410 ;
        RECT 2506.000 2273.960 2510.000 2274.110 ;
        RECT 2533.950 2274.100 2534.330 2274.110 ;
        RECT 703.405 224.210 703.735 224.225 ;
        RECT 2533.950 224.210 2534.330 224.220 ;
        RECT 703.405 223.910 2534.330 224.210 ;
        RECT 703.405 223.895 703.735 223.910 ;
        RECT 2533.950 223.900 2534.330 223.910 ;
      LAYER via3 ;
        RECT 2533.980 2274.100 2534.300 2274.420 ;
        RECT 2533.980 223.900 2534.300 224.220 ;
      LAYER met4 ;
        RECT 2533.975 2274.095 2534.305 2274.425 ;
        RECT 2533.990 224.225 2534.290 2274.095 ;
        RECT 2533.975 223.895 2534.305 224.225 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2622.320 2519.810 2622.380 ;
        RECT 2532.370 2622.320 2532.690 2622.380 ;
        RECT 2519.490 2622.180 2532.690 2622.320 ;
        RECT 2519.490 2622.120 2519.810 2622.180 ;
        RECT 2532.370 2622.120 2532.690 2622.180 ;
        RECT 1358.910 397.020 1359.230 397.080 ;
        RECT 2532.370 397.020 2532.690 397.080 ;
        RECT 1358.910 396.880 2532.690 397.020 ;
        RECT 1358.910 396.820 1359.230 396.880 ;
        RECT 2532.370 396.820 2532.690 396.880 ;
      LAYER via ;
        RECT 2519.520 2622.120 2519.780 2622.380 ;
        RECT 2532.400 2622.120 2532.660 2622.380 ;
        RECT 1358.940 396.820 1359.200 397.080 ;
        RECT 2532.400 396.820 2532.660 397.080 ;
      LAYER met2 ;
        RECT 2519.510 2622.235 2519.790 2622.605 ;
        RECT 2519.520 2622.090 2519.780 2622.235 ;
        RECT 2532.400 2622.090 2532.660 2622.410 ;
        RECT 2532.460 397.110 2532.600 2622.090 ;
        RECT 1358.940 396.790 1359.200 397.110 ;
        RECT 2532.400 396.790 2532.660 397.110 ;
        RECT 1359.000 17.410 1359.140 396.790 ;
        RECT 1358.540 17.270 1359.140 17.410 ;
        RECT 1358.540 2.400 1358.680 17.270 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2622.280 2519.790 2622.560 ;
      LAYER met3 ;
        RECT 2506.000 2622.570 2510.000 2622.720 ;
        RECT 2519.485 2622.570 2519.815 2622.585 ;
        RECT 2506.000 2622.270 2519.815 2622.570 ;
        RECT 2506.000 2622.120 2510.000 2622.270 ;
        RECT 2519.485 2622.255 2519.815 2622.270 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.610 480.320 1379.930 480.380 ;
        RECT 2553.530 480.320 2553.850 480.380 ;
        RECT 1379.610 480.180 2553.850 480.320 ;
        RECT 1379.610 480.120 1379.930 480.180 ;
        RECT 2553.530 480.120 2553.850 480.180 ;
        RECT 1376.390 20.300 1376.710 20.360 ;
        RECT 1379.610 20.300 1379.930 20.360 ;
        RECT 1376.390 20.160 1379.930 20.300 ;
        RECT 1376.390 20.100 1376.710 20.160 ;
        RECT 1379.610 20.100 1379.930 20.160 ;
      LAYER via ;
        RECT 1379.640 480.120 1379.900 480.380 ;
        RECT 2553.560 480.120 2553.820 480.380 ;
        RECT 1376.420 20.100 1376.680 20.360 ;
        RECT 1379.640 20.100 1379.900 20.360 ;
      LAYER met2 ;
        RECT 2248.110 3015.955 2248.390 3016.325 ;
        RECT 2553.550 3015.955 2553.830 3016.325 ;
        RECT 2248.180 3010.000 2248.320 3015.955 ;
        RECT 2248.180 3009.340 2248.530 3010.000 ;
        RECT 2248.250 3006.000 2248.530 3009.340 ;
        RECT 2553.620 480.410 2553.760 3015.955 ;
        RECT 1379.640 480.090 1379.900 480.410 ;
        RECT 2553.560 480.090 2553.820 480.410 ;
        RECT 1379.700 20.390 1379.840 480.090 ;
        RECT 1376.420 20.070 1376.680 20.390 ;
        RECT 1379.640 20.070 1379.900 20.390 ;
        RECT 1376.480 2.400 1376.620 20.070 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
      LAYER via2 ;
        RECT 2248.110 3016.000 2248.390 3016.280 ;
        RECT 2553.550 3016.000 2553.830 3016.280 ;
      LAYER met3 ;
        RECT 2248.085 3016.290 2248.415 3016.305 ;
        RECT 2553.525 3016.290 2553.855 3016.305 ;
        RECT 2248.085 3015.990 2553.855 3016.290 ;
        RECT 2248.085 3015.975 2248.415 3015.990 ;
        RECT 2553.525 3015.975 2553.855 3015.990 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2307.820 2519.810 2307.880 ;
        RECT 2540.190 2307.820 2540.510 2307.880 ;
        RECT 2519.490 2307.680 2540.510 2307.820 ;
        RECT 2519.490 2307.620 2519.810 2307.680 ;
        RECT 2540.190 2307.620 2540.510 2307.680 ;
        RECT 1400.310 444.960 1400.630 445.020 ;
        RECT 2540.190 444.960 2540.510 445.020 ;
        RECT 1400.310 444.820 2540.510 444.960 ;
        RECT 1400.310 444.760 1400.630 444.820 ;
        RECT 2540.190 444.760 2540.510 444.820 ;
        RECT 1394.330 20.300 1394.650 20.360 ;
        RECT 1400.310 20.300 1400.630 20.360 ;
        RECT 1394.330 20.160 1400.630 20.300 ;
        RECT 1394.330 20.100 1394.650 20.160 ;
        RECT 1400.310 20.100 1400.630 20.160 ;
      LAYER via ;
        RECT 2519.520 2307.620 2519.780 2307.880 ;
        RECT 2540.220 2307.620 2540.480 2307.880 ;
        RECT 1400.340 444.760 1400.600 445.020 ;
        RECT 2540.220 444.760 2540.480 445.020 ;
        RECT 1394.360 20.100 1394.620 20.360 ;
        RECT 1400.340 20.100 1400.600 20.360 ;
      LAYER met2 ;
        RECT 2519.510 2310.795 2519.790 2311.165 ;
        RECT 2519.580 2307.910 2519.720 2310.795 ;
        RECT 2519.520 2307.590 2519.780 2307.910 ;
        RECT 2540.220 2307.590 2540.480 2307.910 ;
        RECT 2540.280 445.050 2540.420 2307.590 ;
        RECT 1400.340 444.730 1400.600 445.050 ;
        RECT 2540.220 444.730 2540.480 445.050 ;
        RECT 1400.400 20.390 1400.540 444.730 ;
        RECT 1394.360 20.070 1394.620 20.390 ;
        RECT 1400.340 20.070 1400.600 20.390 ;
        RECT 1394.420 2.400 1394.560 20.070 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2310.840 2519.790 2311.120 ;
      LAYER met3 ;
        RECT 2506.000 2311.130 2510.000 2311.280 ;
        RECT 2519.485 2311.130 2519.815 2311.145 ;
        RECT 2506.000 2310.830 2519.815 2311.130 ;
        RECT 2506.000 2310.680 2510.000 2310.830 ;
        RECT 2519.485 2310.815 2519.815 2310.830 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 378.650 2885.820 378.970 2885.880 ;
        RECT 394.750 2885.820 395.070 2885.880 ;
        RECT 378.650 2885.680 395.070 2885.820 ;
        RECT 378.650 2885.620 378.970 2885.680 ;
        RECT 394.750 2885.620 395.070 2885.680 ;
        RECT 378.650 120.600 378.970 120.660 ;
        RECT 1407.670 120.600 1407.990 120.660 ;
        RECT 378.650 120.460 1407.990 120.600 ;
        RECT 378.650 120.400 378.970 120.460 ;
        RECT 1407.670 120.400 1407.990 120.460 ;
        RECT 1407.670 62.120 1407.990 62.180 ;
        RECT 1412.270 62.120 1412.590 62.180 ;
        RECT 1407.670 61.980 1412.590 62.120 ;
        RECT 1407.670 61.920 1407.990 61.980 ;
        RECT 1412.270 61.920 1412.590 61.980 ;
      LAYER via ;
        RECT 378.680 2885.620 378.940 2885.880 ;
        RECT 394.780 2885.620 395.040 2885.880 ;
        RECT 378.680 120.400 378.940 120.660 ;
        RECT 1407.700 120.400 1407.960 120.660 ;
        RECT 1407.700 61.920 1407.960 62.180 ;
        RECT 1412.300 61.920 1412.560 62.180 ;
      LAYER met2 ;
        RECT 394.770 2887.435 395.050 2887.805 ;
        RECT 394.840 2885.910 394.980 2887.435 ;
        RECT 378.680 2885.590 378.940 2885.910 ;
        RECT 394.780 2885.590 395.040 2885.910 ;
        RECT 378.740 120.690 378.880 2885.590 ;
        RECT 378.680 120.370 378.940 120.690 ;
        RECT 1407.700 120.370 1407.960 120.690 ;
        RECT 1407.760 62.210 1407.900 120.370 ;
        RECT 1407.700 61.890 1407.960 62.210 ;
        RECT 1412.300 61.890 1412.560 62.210 ;
        RECT 1412.360 2.400 1412.500 61.890 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
      LAYER via2 ;
        RECT 394.770 2887.480 395.050 2887.760 ;
      LAYER met3 ;
        RECT 394.745 2887.770 395.075 2887.785 ;
        RECT 410.000 2887.770 414.000 2887.920 ;
        RECT 394.745 2887.470 414.000 2887.770 ;
        RECT 394.745 2887.455 395.075 2887.470 ;
        RECT 410.000 2887.320 414.000 2887.470 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 79.800 1435.130 79.860 ;
        RECT 2513.970 79.800 2514.290 79.860 ;
        RECT 1434.810 79.660 2514.290 79.800 ;
        RECT 1434.810 79.600 1435.130 79.660 ;
        RECT 2513.970 79.600 2514.290 79.660 ;
        RECT 1429.750 16.900 1430.070 16.960 ;
        RECT 1434.810 16.900 1435.130 16.960 ;
        RECT 1429.750 16.760 1435.130 16.900 ;
        RECT 1429.750 16.700 1430.070 16.760 ;
        RECT 1434.810 16.700 1435.130 16.760 ;
      LAYER via ;
        RECT 1434.840 79.600 1435.100 79.860 ;
        RECT 2514.000 79.600 2514.260 79.860 ;
        RECT 1429.780 16.700 1430.040 16.960 ;
        RECT 1434.840 16.700 1435.100 16.960 ;
      LAYER met2 ;
        RECT 2513.990 795.755 2514.270 796.125 ;
        RECT 2514.060 79.890 2514.200 795.755 ;
        RECT 1434.840 79.570 1435.100 79.890 ;
        RECT 2514.000 79.570 2514.260 79.890 ;
        RECT 1434.900 16.990 1435.040 79.570 ;
        RECT 1429.780 16.670 1430.040 16.990 ;
        RECT 1434.840 16.670 1435.100 16.990 ;
        RECT 1429.840 2.400 1429.980 16.670 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 2513.990 795.800 2514.270 796.080 ;
      LAYER met3 ;
        RECT 2506.000 796.090 2510.000 796.240 ;
        RECT 2513.965 796.090 2514.295 796.105 ;
        RECT 2506.000 795.790 2514.295 796.090 ;
        RECT 2506.000 795.640 2510.000 795.790 ;
        RECT 2513.965 795.775 2514.295 795.790 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2186.525 3003.985 2186.695 3006.535 ;
      LAYER mcon ;
        RECT 2186.525 3006.365 2186.695 3006.535 ;
      LAYER met1 ;
        RECT 2186.450 3006.520 2186.770 3006.580 ;
        RECT 2186.255 3006.380 2186.770 3006.520 ;
        RECT 2186.450 3006.320 2186.770 3006.380 ;
        RECT 2186.465 3004.140 2186.755 3004.185 ;
        RECT 2546.630 3004.140 2546.950 3004.200 ;
        RECT 2186.465 3004.000 2546.950 3004.140 ;
        RECT 2186.465 3003.955 2186.755 3004.000 ;
        RECT 2546.630 3003.940 2546.950 3004.000 ;
      LAYER via ;
        RECT 2186.480 3006.320 2186.740 3006.580 ;
        RECT 2546.660 3003.940 2546.920 3004.200 ;
      LAYER met2 ;
        RECT 2185.690 3006.690 2185.970 3010.000 ;
        RECT 2185.690 3006.610 2186.680 3006.690 ;
        RECT 2185.690 3006.550 2186.740 3006.610 ;
        RECT 2185.690 3006.000 2185.970 3006.550 ;
        RECT 2186.480 3006.290 2186.740 3006.550 ;
        RECT 2546.660 3003.910 2546.920 3004.230 ;
        RECT 2546.720 494.885 2546.860 3003.910 ;
        RECT 1448.630 494.515 1448.910 494.885 ;
        RECT 2546.650 494.515 2546.930 494.885 ;
        RECT 1448.700 17.410 1448.840 494.515 ;
        RECT 1447.780 17.270 1448.840 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
      LAYER via2 ;
        RECT 1448.630 494.560 1448.910 494.840 ;
        RECT 2546.650 494.560 2546.930 494.840 ;
      LAYER met3 ;
        RECT 1448.605 494.850 1448.935 494.865 ;
        RECT 2546.625 494.850 2546.955 494.865 ;
        RECT 1448.605 494.550 2546.955 494.850 ;
        RECT 1448.605 494.535 1448.935 494.550 ;
        RECT 2546.625 494.535 2546.955 494.550 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2162.640 2519.810 2162.700 ;
        RECT 2533.750 2162.640 2534.070 2162.700 ;
        RECT 2519.490 2162.500 2534.070 2162.640 ;
        RECT 2519.490 2162.440 2519.810 2162.500 ;
        RECT 2533.750 2162.440 2534.070 2162.500 ;
        RECT 1469.310 438.160 1469.630 438.220 ;
        RECT 2533.750 438.160 2534.070 438.220 ;
        RECT 1469.310 438.020 2534.070 438.160 ;
        RECT 1469.310 437.960 1469.630 438.020 ;
        RECT 2533.750 437.960 2534.070 438.020 ;
        RECT 1465.630 16.900 1465.950 16.960 ;
        RECT 1469.310 16.900 1469.630 16.960 ;
        RECT 1465.630 16.760 1469.630 16.900 ;
        RECT 1465.630 16.700 1465.950 16.760 ;
        RECT 1469.310 16.700 1469.630 16.760 ;
      LAYER via ;
        RECT 2519.520 2162.440 2519.780 2162.700 ;
        RECT 2533.780 2162.440 2534.040 2162.700 ;
        RECT 1469.340 437.960 1469.600 438.220 ;
        RECT 2533.780 437.960 2534.040 438.220 ;
        RECT 1465.660 16.700 1465.920 16.960 ;
        RECT 1469.340 16.700 1469.600 16.960 ;
      LAYER met2 ;
        RECT 2519.510 2165.275 2519.790 2165.645 ;
        RECT 2519.580 2162.730 2519.720 2165.275 ;
        RECT 2519.520 2162.410 2519.780 2162.730 ;
        RECT 2533.780 2162.410 2534.040 2162.730 ;
        RECT 2533.840 438.250 2533.980 2162.410 ;
        RECT 1469.340 437.930 1469.600 438.250 ;
        RECT 2533.780 437.930 2534.040 438.250 ;
        RECT 1469.400 16.990 1469.540 437.930 ;
        RECT 1465.660 16.670 1465.920 16.990 ;
        RECT 1469.340 16.670 1469.600 16.990 ;
        RECT 1465.720 2.400 1465.860 16.670 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2165.320 2519.790 2165.600 ;
      LAYER met3 ;
        RECT 2506.000 2165.610 2510.000 2165.760 ;
        RECT 2519.485 2165.610 2519.815 2165.625 ;
        RECT 2506.000 2165.310 2519.815 2165.610 ;
        RECT 2506.000 2165.160 2510.000 2165.310 ;
        RECT 2519.485 2165.295 2519.815 2165.310 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1373.500 2520.730 1373.560 ;
        RECT 2596.770 1373.500 2597.090 1373.560 ;
        RECT 2520.410 1373.360 2597.090 1373.500 ;
        RECT 2520.410 1373.300 2520.730 1373.360 ;
        RECT 2596.770 1373.300 2597.090 1373.360 ;
        RECT 1490.010 452.100 1490.330 452.160 ;
        RECT 2596.770 452.100 2597.090 452.160 ;
        RECT 1490.010 451.960 2597.090 452.100 ;
        RECT 1490.010 451.900 1490.330 451.960 ;
        RECT 2596.770 451.900 2597.090 451.960 ;
        RECT 1483.570 16.900 1483.890 16.960 ;
        RECT 1490.010 16.900 1490.330 16.960 ;
        RECT 1483.570 16.760 1490.330 16.900 ;
        RECT 1483.570 16.700 1483.890 16.760 ;
        RECT 1490.010 16.700 1490.330 16.760 ;
      LAYER via ;
        RECT 2520.440 1373.300 2520.700 1373.560 ;
        RECT 2596.800 1373.300 2597.060 1373.560 ;
        RECT 1490.040 451.900 1490.300 452.160 ;
        RECT 2596.800 451.900 2597.060 452.160 ;
        RECT 1483.600 16.700 1483.860 16.960 ;
        RECT 1490.040 16.700 1490.300 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1379.195 2520.710 1379.565 ;
        RECT 2520.500 1373.590 2520.640 1379.195 ;
        RECT 2520.440 1373.270 2520.700 1373.590 ;
        RECT 2596.800 1373.270 2597.060 1373.590 ;
        RECT 2596.860 452.190 2597.000 1373.270 ;
        RECT 1490.040 451.870 1490.300 452.190 ;
        RECT 2596.800 451.870 2597.060 452.190 ;
        RECT 1490.100 16.990 1490.240 451.870 ;
        RECT 1483.600 16.670 1483.860 16.990 ;
        RECT 1490.040 16.670 1490.300 16.990 ;
        RECT 1483.660 2.400 1483.800 16.670 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1379.240 2520.710 1379.520 ;
      LAYER met3 ;
        RECT 2506.000 1379.530 2510.000 1379.680 ;
        RECT 2520.405 1379.530 2520.735 1379.545 ;
        RECT 2506.000 1379.230 2520.735 1379.530 ;
        RECT 2506.000 1379.080 2510.000 1379.230 ;
        RECT 2520.405 1379.215 2520.735 1379.230 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1506.570 3015.700 1506.890 3015.760 ;
        RECT 1731.970 3015.700 1732.290 3015.760 ;
        RECT 1506.570 3015.560 1732.290 3015.700 ;
        RECT 1506.570 3015.500 1506.890 3015.560 ;
        RECT 1731.970 3015.500 1732.290 3015.560 ;
        RECT 2415.070 455.500 2415.390 455.560 ;
        RECT 2443.130 455.500 2443.450 455.560 ;
        RECT 2415.070 455.360 2443.450 455.500 ;
        RECT 2415.070 455.300 2415.390 455.360 ;
        RECT 2443.130 455.300 2443.450 455.360 ;
        RECT 2414.610 421.160 2414.930 421.220 ;
        RECT 2394.460 421.020 2414.930 421.160 ;
        RECT 2380.570 420.820 2380.890 420.880 ;
        RECT 2394.460 420.820 2394.600 421.020 ;
        RECT 2414.610 420.960 2414.930 421.020 ;
        RECT 2380.570 420.680 2394.600 420.820 ;
        RECT 2380.570 420.620 2380.890 420.680 ;
        RECT 2373.210 400.420 2373.530 400.480 ;
        RECT 2380.570 400.420 2380.890 400.480 ;
        RECT 2373.210 400.280 2380.890 400.420 ;
        RECT 2373.210 400.220 2373.530 400.280 ;
        RECT 2380.570 400.220 2380.890 400.280 ;
        RECT 2356.190 390.560 2356.510 390.620 ;
        RECT 2373.210 390.560 2373.530 390.620 ;
        RECT 2356.190 390.420 2373.530 390.560 ;
        RECT 2356.190 390.360 2356.510 390.420 ;
        RECT 2373.210 390.360 2373.530 390.420 ;
        RECT 2346.530 359.960 2346.850 360.020 ;
        RECT 2356.190 359.960 2356.510 360.020 ;
        RECT 2346.530 359.820 2356.510 359.960 ;
        RECT 2346.530 359.760 2346.850 359.820 ;
        RECT 2356.190 359.760 2356.510 359.820 ;
        RECT 2335.490 337.520 2335.810 337.580 ;
        RECT 2346.530 337.520 2346.850 337.580 ;
        RECT 2335.490 337.380 2346.850 337.520 ;
        RECT 2335.490 337.320 2335.810 337.380 ;
        RECT 2346.530 337.320 2346.850 337.380 ;
        RECT 2328.590 117.540 2328.910 117.600 ;
        RECT 2335.490 117.540 2335.810 117.600 ;
        RECT 2328.590 117.400 2335.810 117.540 ;
        RECT 2328.590 117.340 2328.910 117.400 ;
        RECT 2335.490 117.340 2335.810 117.400 ;
        RECT 2311.570 44.440 2311.890 44.500 ;
        RECT 2328.590 44.440 2328.910 44.500 ;
        RECT 2311.570 44.300 2328.910 44.440 ;
        RECT 2311.570 44.240 2311.890 44.300 ;
        RECT 2328.590 44.240 2328.910 44.300 ;
        RECT 1893.430 25.400 1893.750 25.460 ;
        RECT 2311.110 25.400 2311.430 25.460 ;
        RECT 1893.430 25.260 2311.430 25.400 ;
        RECT 1893.430 25.200 1893.750 25.260 ;
        RECT 2311.110 25.200 2311.430 25.260 ;
        RECT 1501.510 18.940 1501.830 19.000 ;
        RECT 1893.430 18.940 1893.750 19.000 ;
        RECT 1501.510 18.800 1893.750 18.940 ;
        RECT 1501.510 18.740 1501.830 18.800 ;
        RECT 1893.430 18.740 1893.750 18.800 ;
      LAYER via ;
        RECT 1506.600 3015.500 1506.860 3015.760 ;
        RECT 1732.000 3015.500 1732.260 3015.760 ;
        RECT 2415.100 455.300 2415.360 455.560 ;
        RECT 2443.160 455.300 2443.420 455.560 ;
        RECT 2380.600 420.620 2380.860 420.880 ;
        RECT 2414.640 420.960 2414.900 421.220 ;
        RECT 2373.240 400.220 2373.500 400.480 ;
        RECT 2380.600 400.220 2380.860 400.480 ;
        RECT 2356.220 390.360 2356.480 390.620 ;
        RECT 2373.240 390.360 2373.500 390.620 ;
        RECT 2346.560 359.760 2346.820 360.020 ;
        RECT 2356.220 359.760 2356.480 360.020 ;
        RECT 2335.520 337.320 2335.780 337.580 ;
        RECT 2346.560 337.320 2346.820 337.580 ;
        RECT 2328.620 117.340 2328.880 117.600 ;
        RECT 2335.520 117.340 2335.780 117.600 ;
        RECT 2311.600 44.240 2311.860 44.500 ;
        RECT 2328.620 44.240 2328.880 44.500 ;
        RECT 1893.460 25.200 1893.720 25.460 ;
        RECT 2311.140 25.200 2311.400 25.460 ;
        RECT 1501.540 18.740 1501.800 19.000 ;
        RECT 1893.460 18.740 1893.720 19.000 ;
      LAYER met2 ;
        RECT 1506.600 3015.470 1506.860 3015.790 ;
        RECT 1732.000 3015.470 1732.260 3015.790 ;
        RECT 1506.660 3010.000 1506.800 3015.470 ;
        RECT 1732.060 3012.245 1732.200 3015.470 ;
        RECT 1731.990 3011.875 1732.270 3012.245 ;
        RECT 1506.660 3009.340 1507.010 3010.000 ;
        RECT 1506.730 3006.000 1507.010 3009.340 ;
        RECT 2443.150 482.955 2443.430 483.325 ;
        RECT 2443.220 455.590 2443.360 482.955 ;
        RECT 2415.100 455.270 2415.360 455.590 ;
        RECT 2443.160 455.270 2443.420 455.590 ;
        RECT 2415.160 428.130 2415.300 455.270 ;
        RECT 2414.700 427.990 2415.300 428.130 ;
        RECT 2414.700 421.250 2414.840 427.990 ;
        RECT 2414.640 420.930 2414.900 421.250 ;
        RECT 2380.600 420.590 2380.860 420.910 ;
        RECT 2380.660 400.510 2380.800 420.590 ;
        RECT 2373.240 400.190 2373.500 400.510 ;
        RECT 2380.600 400.190 2380.860 400.510 ;
        RECT 2373.300 390.650 2373.440 400.190 ;
        RECT 2356.220 390.330 2356.480 390.650 ;
        RECT 2373.240 390.330 2373.500 390.650 ;
        RECT 2356.280 360.050 2356.420 390.330 ;
        RECT 2346.560 359.730 2346.820 360.050 ;
        RECT 2356.220 359.730 2356.480 360.050 ;
        RECT 2346.620 337.610 2346.760 359.730 ;
        RECT 2335.520 337.290 2335.780 337.610 ;
        RECT 2346.560 337.290 2346.820 337.610 ;
        RECT 2335.580 117.630 2335.720 337.290 ;
        RECT 2328.620 117.310 2328.880 117.630 ;
        RECT 2335.520 117.310 2335.780 117.630 ;
        RECT 2328.680 44.530 2328.820 117.310 ;
        RECT 2311.600 44.210 2311.860 44.530 ;
        RECT 2328.620 44.210 2328.880 44.530 ;
        RECT 2311.660 41.210 2311.800 44.210 ;
        RECT 2311.200 41.070 2311.800 41.210 ;
        RECT 2311.200 25.490 2311.340 41.070 ;
        RECT 1893.460 25.170 1893.720 25.490 ;
        RECT 2311.140 25.170 2311.400 25.490 ;
        RECT 1893.520 19.030 1893.660 25.170 ;
        RECT 1501.540 18.710 1501.800 19.030 ;
        RECT 1893.460 18.710 1893.720 19.030 ;
        RECT 1501.600 2.400 1501.740 18.710 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
      LAYER via2 ;
        RECT 1731.990 3011.920 1732.270 3012.200 ;
        RECT 2443.150 483.000 2443.430 483.280 ;
      LAYER met3 ;
        RECT 1731.965 3012.210 1732.295 3012.225 ;
        RECT 2414.350 3012.210 2414.730 3012.220 ;
        RECT 1731.965 3011.910 2414.730 3012.210 ;
        RECT 1731.965 3011.895 1732.295 3011.910 ;
        RECT 2414.350 3011.900 2414.730 3011.910 ;
        RECT 2414.350 2999.970 2414.730 2999.980 ;
        RECT 2449.310 2999.970 2449.690 2999.980 ;
        RECT 2414.350 2999.670 2449.690 2999.970 ;
        RECT 2414.350 2999.660 2414.730 2999.670 ;
        RECT 2449.310 2999.660 2449.690 2999.670 ;
        RECT 2443.125 483.290 2443.455 483.305 ;
        RECT 2449.310 483.290 2449.690 483.300 ;
        RECT 2443.125 482.990 2449.690 483.290 ;
        RECT 2443.125 482.975 2443.455 482.990 ;
        RECT 2449.310 482.980 2449.690 482.990 ;
      LAYER via3 ;
        RECT 2414.380 3011.900 2414.700 3012.220 ;
        RECT 2414.380 2999.660 2414.700 2999.980 ;
        RECT 2449.340 2999.660 2449.660 2999.980 ;
        RECT 2449.340 482.980 2449.660 483.300 ;
      LAYER met4 ;
        RECT 2414.375 3011.895 2414.705 3012.225 ;
        RECT 2414.390 2999.985 2414.690 3011.895 ;
        RECT 2414.375 2999.655 2414.705 2999.985 ;
        RECT 2449.335 2999.655 2449.665 2999.985 ;
        RECT 2449.350 2021.450 2449.650 2999.655 ;
        RECT 2449.350 2021.150 2450.570 2021.450 ;
        RECT 2450.270 2001.050 2450.570 2021.150 ;
        RECT 2449.350 2000.750 2450.570 2001.050 ;
        RECT 2449.350 483.305 2449.650 2000.750 ;
        RECT 2449.335 482.975 2449.665 483.305 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1518.990 16.900 1519.310 16.960 ;
        RECT 1524.510 16.900 1524.830 16.960 ;
        RECT 1518.990 16.760 1524.830 16.900 ;
        RECT 1518.990 16.700 1519.310 16.760 ;
        RECT 1524.510 16.700 1524.830 16.760 ;
      LAYER via ;
        RECT 1519.020 16.700 1519.280 16.960 ;
        RECT 1524.540 16.700 1524.800 16.960 ;
      LAYER met2 ;
        RECT 1654.710 3037.715 1654.990 3038.085 ;
        RECT 1654.780 3010.000 1654.920 3037.715 ;
        RECT 1654.780 3009.340 1655.130 3010.000 ;
        RECT 1654.850 3006.000 1655.130 3009.340 ;
        RECT 2415.090 510.835 2415.370 511.205 ;
        RECT 2415.160 486.725 2415.300 510.835 ;
        RECT 1524.530 486.355 1524.810 486.725 ;
        RECT 2415.090 486.355 2415.370 486.725 ;
        RECT 1524.600 16.990 1524.740 486.355 ;
        RECT 1519.020 16.670 1519.280 16.990 ;
        RECT 1524.540 16.670 1524.800 16.990 ;
        RECT 1519.080 2.400 1519.220 16.670 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
      LAYER via2 ;
        RECT 1654.710 3037.760 1654.990 3038.040 ;
        RECT 2415.090 510.880 2415.370 511.160 ;
        RECT 1524.530 486.400 1524.810 486.680 ;
        RECT 2415.090 486.400 2415.370 486.680 ;
      LAYER met3 ;
        RECT 1654.685 3038.050 1655.015 3038.065 ;
        RECT 2449.310 3038.050 2449.690 3038.060 ;
        RECT 1654.685 3037.750 2449.690 3038.050 ;
        RECT 1654.685 3037.735 1655.015 3037.750 ;
        RECT 2449.310 3037.740 2449.690 3037.750 ;
        RECT 2415.065 511.170 2415.395 511.185 ;
        RECT 2435.510 511.170 2435.890 511.180 ;
        RECT 2415.065 510.870 2435.890 511.170 ;
        RECT 2415.065 510.855 2415.395 510.870 ;
        RECT 2435.510 510.860 2435.890 510.870 ;
        RECT 1524.505 486.690 1524.835 486.705 ;
        RECT 2415.065 486.690 2415.395 486.705 ;
        RECT 1524.505 486.390 2415.395 486.690 ;
        RECT 1524.505 486.375 1524.835 486.390 ;
        RECT 2415.065 486.375 2415.395 486.390 ;
      LAYER via3 ;
        RECT 2449.340 3037.740 2449.660 3038.060 ;
        RECT 2435.540 510.860 2435.860 511.180 ;
      LAYER met4 ;
        RECT 2449.335 3037.735 2449.665 3038.065 ;
        RECT 2449.350 3007.450 2449.650 3037.735 ;
        RECT 2448.430 3007.150 2449.650 3007.450 ;
        RECT 2448.430 2959.850 2448.730 3007.150 ;
        RECT 2446.590 2959.550 2448.730 2959.850 ;
        RECT 2446.590 2908.850 2446.890 2959.550 ;
        RECT 2446.590 2908.550 2447.810 2908.850 ;
        RECT 2447.510 2011.250 2447.810 2908.550 ;
        RECT 2445.670 2010.950 2447.810 2011.250 ;
        RECT 2445.670 1950.050 2445.970 2010.950 ;
        RECT 2445.670 1949.750 2448.730 1950.050 ;
        RECT 2448.430 1922.850 2448.730 1949.750 ;
        RECT 2443.830 1922.550 2448.730 1922.850 ;
        RECT 2443.830 1875.690 2444.130 1922.550 ;
        RECT 2436.030 1874.510 2437.210 1875.690 ;
        RECT 2443.390 1874.510 2444.570 1875.690 ;
        RECT 2436.470 1827.650 2436.770 1874.510 ;
        RECT 2436.470 1827.350 2437.690 1827.650 ;
        RECT 2437.390 1800.450 2437.690 1827.350 ;
        RECT 2437.390 1800.150 2438.610 1800.450 ;
        RECT 2438.310 1780.050 2438.610 1800.150 ;
        RECT 2437.390 1779.750 2438.610 1780.050 ;
        RECT 2437.390 1742.650 2437.690 1779.750 ;
        RECT 2436.470 1742.350 2437.690 1742.650 ;
        RECT 2436.470 1708.650 2436.770 1742.350 ;
        RECT 2436.470 1708.350 2438.610 1708.650 ;
        RECT 2438.310 1684.850 2438.610 1708.350 ;
        RECT 2437.390 1684.550 2438.610 1684.850 ;
        RECT 2437.390 1657.650 2437.690 1684.550 ;
        RECT 2437.390 1657.350 2438.610 1657.650 ;
        RECT 2438.310 1620.250 2438.610 1657.350 ;
        RECT 2438.310 1619.950 2440.450 1620.250 ;
        RECT 2440.150 1593.050 2440.450 1619.950 ;
        RECT 2438.310 1592.750 2440.450 1593.050 ;
        RECT 2438.310 1528.450 2438.610 1592.750 ;
        RECT 2437.390 1528.150 2438.610 1528.450 ;
        RECT 2437.390 1491.050 2437.690 1528.150 ;
        RECT 2436.470 1490.750 2437.690 1491.050 ;
        RECT 2436.470 1028.650 2436.770 1490.750 ;
        RECT 2436.470 1028.350 2438.610 1028.650 ;
        RECT 2438.310 981.050 2438.610 1028.350 ;
        RECT 2435.550 980.750 2438.610 981.050 ;
        RECT 2435.550 926.650 2435.850 980.750 ;
        RECT 2435.550 926.350 2436.770 926.650 ;
        RECT 2436.470 909.650 2436.770 926.350 ;
        RECT 2436.470 909.350 2438.610 909.650 ;
        RECT 2438.310 855.250 2438.610 909.350 ;
        RECT 2437.390 854.950 2438.610 855.250 ;
        RECT 2437.390 787.250 2437.690 854.950 ;
        RECT 2436.470 786.950 2437.690 787.250 ;
        RECT 2436.470 770.250 2436.770 786.950 ;
        RECT 2434.630 769.950 2436.770 770.250 ;
        RECT 2434.630 726.490 2434.930 769.950 ;
        RECT 2434.190 725.310 2435.370 726.490 ;
        RECT 2434.190 721.910 2435.370 723.090 ;
        RECT 2434.630 678.450 2434.930 721.910 ;
        RECT 2434.630 678.150 2438.610 678.450 ;
        RECT 2438.310 620.650 2438.610 678.150 ;
        RECT 2437.390 620.350 2438.610 620.650 ;
        RECT 2437.390 573.050 2437.690 620.350 ;
        RECT 2435.550 572.750 2437.690 573.050 ;
        RECT 2435.550 511.185 2435.850 572.750 ;
        RECT 2435.535 510.855 2435.865 511.185 ;
      LAYER met5 ;
        RECT 2435.820 1874.300 2444.780 1875.900 ;
        RECT 2433.980 725.100 2438.340 726.700 ;
        RECT 2436.740 723.300 2438.340 725.100 ;
        RECT 2433.980 721.700 2438.340 723.300 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.050 3012.980 351.370 3013.040 ;
        RECT 1160.650 3012.980 1160.970 3013.040 ;
        RECT 351.050 3012.840 1160.970 3012.980 ;
        RECT 351.050 3012.780 351.370 3012.840 ;
        RECT 1160.650 3012.780 1160.970 3012.840 ;
        RECT 351.050 495.960 351.370 496.020 ;
        RECT 710.770 495.960 711.090 496.020 ;
        RECT 351.050 495.820 711.090 495.960 ;
        RECT 351.050 495.760 351.370 495.820 ;
        RECT 710.770 495.760 711.090 495.820 ;
        RECT 710.770 20.300 711.090 20.360 ;
        RECT 716.290 20.300 716.610 20.360 ;
        RECT 710.770 20.160 716.610 20.300 ;
        RECT 710.770 20.100 711.090 20.160 ;
        RECT 716.290 20.100 716.610 20.160 ;
      LAYER via ;
        RECT 351.080 3012.780 351.340 3013.040 ;
        RECT 1160.680 3012.780 1160.940 3013.040 ;
        RECT 351.080 495.760 351.340 496.020 ;
        RECT 710.800 495.760 711.060 496.020 ;
        RECT 710.800 20.100 711.060 20.360 ;
        RECT 716.320 20.100 716.580 20.360 ;
      LAYER met2 ;
        RECT 351.080 3012.750 351.340 3013.070 ;
        RECT 1160.680 3012.750 1160.940 3013.070 ;
        RECT 351.140 496.050 351.280 3012.750 ;
        RECT 1160.740 3010.000 1160.880 3012.750 ;
        RECT 1160.740 3009.340 1161.090 3010.000 ;
        RECT 1160.810 3006.000 1161.090 3009.340 ;
        RECT 351.080 495.730 351.340 496.050 ;
        RECT 710.800 495.730 711.060 496.050 ;
        RECT 710.860 20.390 711.000 495.730 ;
        RECT 710.800 20.070 711.060 20.390 ;
        RECT 716.320 20.070 716.580 20.390 ;
        RECT 716.380 2.400 716.520 20.070 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2509.830 2118.440 2510.150 2118.500 ;
        RECT 2510.290 2118.440 2510.610 2118.500 ;
        RECT 2509.830 2118.300 2510.610 2118.440 ;
        RECT 2509.830 2118.240 2510.150 2118.300 ;
        RECT 2510.290 2118.240 2510.610 2118.300 ;
      LAYER via ;
        RECT 2509.860 2118.240 2510.120 2118.500 ;
        RECT 2510.320 2118.240 2510.580 2118.500 ;
      LAYER met2 ;
        RECT 2136.930 3008.730 2137.210 3010.000 ;
        RECT 2138.630 3008.730 2138.910 3008.845 ;
        RECT 2136.930 3008.590 2138.910 3008.730 ;
        RECT 2136.930 3006.000 2137.210 3008.590 ;
        RECT 2138.630 3008.475 2138.910 3008.590 ;
        RECT 2509.390 2623.595 2509.670 2623.965 ;
        RECT 2509.460 2611.725 2509.600 2623.595 ;
        RECT 2509.390 2611.355 2509.670 2611.725 ;
        RECT 2510.310 2538.595 2510.590 2538.965 ;
        RECT 2510.380 2492.045 2510.520 2538.595 ;
        RECT 2510.310 2491.675 2510.590 2492.045 ;
        RECT 2509.850 2407.355 2510.130 2407.725 ;
        RECT 2509.920 2360.125 2510.060 2407.355 ;
        RECT 2509.850 2359.755 2510.130 2360.125 ;
        RECT 2510.310 2359.075 2510.590 2359.445 ;
        RECT 2510.380 2313.205 2510.520 2359.075 ;
        RECT 2510.310 2312.835 2510.590 2313.205 ;
        RECT 2509.850 2294.475 2510.130 2294.845 ;
        RECT 2509.920 2263.565 2510.060 2294.475 ;
        RECT 2509.850 2263.195 2510.130 2263.565 ;
        RECT 2510.310 2214.235 2510.590 2214.605 ;
        RECT 2510.380 2167.005 2510.520 2214.235 ;
        RECT 2510.310 2166.635 2510.590 2167.005 ;
        RECT 2510.310 2142.155 2510.590 2142.525 ;
        RECT 2510.380 2118.530 2510.520 2142.155 ;
        RECT 2509.860 2118.210 2510.120 2118.530 ;
        RECT 2510.320 2118.210 2510.580 2118.530 ;
        RECT 2509.920 2077.245 2510.060 2118.210 ;
        RECT 2509.850 2076.875 2510.130 2077.245 ;
        RECT 2510.310 2069.395 2510.590 2069.765 ;
        RECT 2510.380 2022.845 2510.520 2069.395 ;
        RECT 2510.310 2022.475 2510.590 2022.845 ;
        RECT 2510.310 1972.835 2510.590 1973.205 ;
        RECT 2510.380 1926.285 2510.520 1972.835 ;
        RECT 2510.310 1925.915 2510.590 1926.285 ;
        RECT 2510.310 1804.195 2510.590 1804.565 ;
        RECT 2510.380 1780.765 2510.520 1804.195 ;
        RECT 2510.310 1780.395 2510.590 1780.765 ;
        RECT 2511.230 1772.915 2511.510 1773.285 ;
        RECT 2511.300 1726.365 2511.440 1772.915 ;
        RECT 2511.230 1725.995 2511.510 1726.365 ;
        RECT 2510.310 1676.355 2510.590 1676.725 ;
        RECT 2510.380 1629.125 2510.520 1676.355 ;
        RECT 2510.310 1628.755 2510.590 1629.125 ;
        RECT 2509.850 1143.915 2510.130 1144.285 ;
        RECT 2509.920 1104.845 2510.060 1143.915 ;
        RECT 2509.850 1104.475 2510.130 1104.845 ;
        RECT 1538.330 512.875 1538.610 513.245 ;
        RECT 1538.400 17.410 1538.540 512.875 ;
        RECT 1537.020 17.270 1538.540 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
      LAYER via2 ;
        RECT 2138.630 3008.520 2138.910 3008.800 ;
        RECT 2509.390 2623.640 2509.670 2623.920 ;
        RECT 2509.390 2611.400 2509.670 2611.680 ;
        RECT 2510.310 2538.640 2510.590 2538.920 ;
        RECT 2510.310 2491.720 2510.590 2492.000 ;
        RECT 2509.850 2407.400 2510.130 2407.680 ;
        RECT 2509.850 2359.800 2510.130 2360.080 ;
        RECT 2510.310 2359.120 2510.590 2359.400 ;
        RECT 2510.310 2312.880 2510.590 2313.160 ;
        RECT 2509.850 2294.520 2510.130 2294.800 ;
        RECT 2509.850 2263.240 2510.130 2263.520 ;
        RECT 2510.310 2214.280 2510.590 2214.560 ;
        RECT 2510.310 2166.680 2510.590 2166.960 ;
        RECT 2510.310 2142.200 2510.590 2142.480 ;
        RECT 2509.850 2076.920 2510.130 2077.200 ;
        RECT 2510.310 2069.440 2510.590 2069.720 ;
        RECT 2510.310 2022.520 2510.590 2022.800 ;
        RECT 2510.310 1972.880 2510.590 1973.160 ;
        RECT 2510.310 1925.960 2510.590 1926.240 ;
        RECT 2510.310 1804.240 2510.590 1804.520 ;
        RECT 2510.310 1780.440 2510.590 1780.720 ;
        RECT 2511.230 1772.960 2511.510 1773.240 ;
        RECT 2511.230 1726.040 2511.510 1726.320 ;
        RECT 2510.310 1676.400 2510.590 1676.680 ;
        RECT 2510.310 1628.800 2510.590 1629.080 ;
        RECT 2509.850 1143.960 2510.130 1144.240 ;
        RECT 2509.850 1104.520 2510.130 1104.800 ;
        RECT 1538.330 512.920 1538.610 513.200 ;
      LAYER met3 ;
        RECT 2138.605 3008.810 2138.935 3008.825 ;
        RECT 2508.190 3008.810 2508.570 3008.820 ;
        RECT 2138.605 3008.510 2508.570 3008.810 ;
        RECT 2138.605 3008.495 2138.935 3008.510 ;
        RECT 2508.190 3008.500 2508.570 3008.510 ;
        RECT 2508.190 2946.620 2508.570 2946.940 ;
        RECT 2508.230 2945.570 2508.530 2946.620 ;
        RECT 2509.110 2945.570 2509.490 2945.580 ;
        RECT 2508.230 2945.270 2509.490 2945.570 ;
        RECT 2509.110 2945.260 2509.490 2945.270 ;
        RECT 2508.190 2898.340 2508.570 2898.660 ;
        RECT 2508.230 2897.980 2508.530 2898.340 ;
        RECT 2508.190 2897.660 2508.570 2897.980 ;
        RECT 2508.190 2774.580 2508.570 2774.900 ;
        RECT 2508.230 2774.210 2508.530 2774.580 ;
        RECT 2509.110 2774.210 2509.490 2774.220 ;
        RECT 2508.230 2773.910 2509.490 2774.210 ;
        RECT 2509.110 2773.900 2509.490 2773.910 ;
        RECT 2509.365 2623.930 2509.695 2623.945 ;
        RECT 2510.030 2623.930 2510.410 2623.940 ;
        RECT 2509.365 2623.630 2510.410 2623.930 ;
        RECT 2509.365 2623.615 2509.695 2623.630 ;
        RECT 2510.030 2623.620 2510.410 2623.630 ;
        RECT 2509.365 2611.700 2509.695 2611.705 ;
        RECT 2509.110 2611.690 2509.695 2611.700 ;
        RECT 2508.910 2611.390 2509.695 2611.690 ;
        RECT 2509.110 2611.380 2509.695 2611.390 ;
        RECT 2509.365 2611.375 2509.695 2611.380 ;
        RECT 2510.285 2538.940 2510.615 2538.945 ;
        RECT 2510.030 2538.930 2510.615 2538.940 ;
        RECT 2510.030 2538.630 2510.840 2538.930 ;
        RECT 2510.030 2538.620 2510.615 2538.630 ;
        RECT 2510.285 2538.615 2510.615 2538.620 ;
        RECT 2510.285 2492.010 2510.615 2492.025 ;
        RECT 2510.070 2491.695 2510.615 2492.010 ;
        RECT 2510.070 2491.340 2510.370 2491.695 ;
        RECT 2510.030 2491.020 2510.410 2491.340 ;
        RECT 2508.190 2437.610 2508.570 2437.620 ;
        RECT 2510.030 2437.610 2510.410 2437.620 ;
        RECT 2508.190 2437.310 2510.410 2437.610 ;
        RECT 2508.190 2437.300 2508.570 2437.310 ;
        RECT 2510.030 2437.300 2510.410 2437.310 ;
        RECT 2509.825 2407.700 2510.155 2407.705 ;
        RECT 2509.825 2407.690 2510.410 2407.700 ;
        RECT 2509.600 2407.390 2510.410 2407.690 ;
        RECT 2509.825 2407.380 2510.410 2407.390 ;
        RECT 2509.825 2407.375 2510.155 2407.380 ;
        RECT 2509.825 2360.100 2510.155 2360.105 ;
        RECT 2509.825 2360.090 2510.410 2360.100 ;
        RECT 2509.825 2359.790 2510.610 2360.090 ;
        RECT 2509.825 2359.780 2510.410 2359.790 ;
        RECT 2509.825 2359.775 2510.155 2359.780 ;
        RECT 2510.285 2359.420 2510.615 2359.425 ;
        RECT 2510.030 2359.410 2510.615 2359.420 ;
        RECT 2510.030 2359.110 2510.840 2359.410 ;
        RECT 2510.030 2359.100 2510.615 2359.110 ;
        RECT 2510.285 2359.095 2510.615 2359.100 ;
        RECT 2510.285 2313.180 2510.615 2313.185 ;
        RECT 2510.030 2313.170 2510.615 2313.180 ;
        RECT 2509.830 2312.870 2510.615 2313.170 ;
        RECT 2510.030 2312.860 2510.615 2312.870 ;
        RECT 2510.285 2312.855 2510.615 2312.860 ;
        RECT 2508.190 2294.810 2508.570 2294.820 ;
        RECT 2509.825 2294.810 2510.155 2294.825 ;
        RECT 2508.190 2294.510 2510.155 2294.810 ;
        RECT 2508.190 2294.500 2508.570 2294.510 ;
        RECT 2509.825 2294.495 2510.155 2294.510 ;
        RECT 2509.825 2263.540 2510.155 2263.545 ;
        RECT 2509.825 2263.530 2510.410 2263.540 ;
        RECT 2509.825 2263.230 2510.610 2263.530 ;
        RECT 2509.825 2263.220 2510.410 2263.230 ;
        RECT 2509.825 2263.215 2510.155 2263.220 ;
        RECT 2510.285 2214.580 2510.615 2214.585 ;
        RECT 2510.030 2214.570 2510.615 2214.580 ;
        RECT 2510.030 2214.270 2510.840 2214.570 ;
        RECT 2510.030 2214.260 2510.615 2214.270 ;
        RECT 2510.285 2214.255 2510.615 2214.260 ;
        RECT 2510.285 2166.980 2510.615 2166.985 ;
        RECT 2510.030 2166.970 2510.615 2166.980 ;
        RECT 2509.830 2166.670 2510.615 2166.970 ;
        RECT 2510.030 2166.660 2510.615 2166.670 ;
        RECT 2510.285 2166.655 2510.615 2166.660 ;
        RECT 2510.285 2142.500 2510.615 2142.505 ;
        RECT 2510.030 2142.490 2510.615 2142.500 ;
        RECT 2510.030 2142.190 2510.840 2142.490 ;
        RECT 2510.030 2142.180 2510.615 2142.190 ;
        RECT 2510.285 2142.175 2510.615 2142.180 ;
        RECT 2509.825 2077.220 2510.155 2077.225 ;
        RECT 2509.825 2077.210 2510.410 2077.220 ;
        RECT 2509.825 2076.910 2510.610 2077.210 ;
        RECT 2509.825 2076.900 2510.410 2076.910 ;
        RECT 2509.825 2076.895 2510.155 2076.900 ;
        RECT 2510.285 2069.740 2510.615 2069.745 ;
        RECT 2510.030 2069.730 2510.615 2069.740 ;
        RECT 2510.030 2069.430 2510.840 2069.730 ;
        RECT 2510.030 2069.420 2510.615 2069.430 ;
        RECT 2510.285 2069.415 2510.615 2069.420 ;
        RECT 2510.285 2022.810 2510.615 2022.825 ;
        RECT 2510.070 2022.495 2510.615 2022.810 ;
        RECT 2510.070 2022.140 2510.370 2022.495 ;
        RECT 2510.030 2021.820 2510.410 2022.140 ;
        RECT 2510.285 1973.180 2510.615 1973.185 ;
        RECT 2510.030 1973.170 2510.615 1973.180 ;
        RECT 2510.030 1972.870 2510.840 1973.170 ;
        RECT 2510.030 1972.860 2510.615 1972.870 ;
        RECT 2510.285 1972.855 2510.615 1972.860 ;
        RECT 2510.285 1926.250 2510.615 1926.265 ;
        RECT 2510.070 1925.935 2510.615 1926.250 ;
        RECT 2510.070 1925.580 2510.370 1925.935 ;
        RECT 2510.030 1925.260 2510.410 1925.580 ;
        RECT 2509.110 1804.530 2509.490 1804.540 ;
        RECT 2510.285 1804.530 2510.615 1804.545 ;
        RECT 2509.110 1804.230 2510.615 1804.530 ;
        RECT 2509.110 1804.220 2509.490 1804.230 ;
        RECT 2510.285 1804.215 2510.615 1804.230 ;
        RECT 2510.285 1780.730 2510.615 1780.745 ;
        RECT 2510.950 1780.730 2511.330 1780.740 ;
        RECT 2510.285 1780.430 2511.330 1780.730 ;
        RECT 2510.285 1780.415 2510.615 1780.430 ;
        RECT 2510.950 1780.420 2511.330 1780.430 ;
        RECT 2511.205 1773.260 2511.535 1773.265 ;
        RECT 2510.950 1773.250 2511.535 1773.260 ;
        RECT 2510.950 1772.950 2511.760 1773.250 ;
        RECT 2510.950 1772.940 2511.535 1772.950 ;
        RECT 2511.205 1772.935 2511.535 1772.940 ;
        RECT 2511.205 1726.330 2511.535 1726.345 ;
        RECT 2510.990 1726.015 2511.535 1726.330 ;
        RECT 2510.990 1725.660 2511.290 1726.015 ;
        RECT 2510.950 1725.340 2511.330 1725.660 ;
        RECT 2510.950 1698.450 2511.330 1698.460 ;
        RECT 2510.070 1698.150 2511.330 1698.450 ;
        RECT 2510.070 1697.100 2510.370 1698.150 ;
        RECT 2510.950 1698.140 2511.330 1698.150 ;
        RECT 2510.030 1696.780 2510.410 1697.100 ;
        RECT 2510.285 1676.700 2510.615 1676.705 ;
        RECT 2510.030 1676.690 2510.615 1676.700 ;
        RECT 2509.830 1676.390 2510.615 1676.690 ;
        RECT 2510.030 1676.380 2510.615 1676.390 ;
        RECT 2510.285 1676.375 2510.615 1676.380 ;
        RECT 2510.285 1629.090 2510.615 1629.105 ;
        RECT 2510.950 1629.090 2511.330 1629.100 ;
        RECT 2510.285 1628.790 2511.330 1629.090 ;
        RECT 2510.285 1628.775 2510.615 1628.790 ;
        RECT 2510.950 1628.780 2511.330 1628.790 ;
        RECT 2509.110 1346.210 2509.490 1346.220 ;
        RECT 2510.030 1346.210 2510.410 1346.220 ;
        RECT 2509.110 1345.910 2510.410 1346.210 ;
        RECT 2509.110 1345.900 2509.490 1345.910 ;
        RECT 2510.030 1345.900 2510.410 1345.910 ;
        RECT 2508.190 1144.250 2508.570 1144.260 ;
        RECT 2509.825 1144.250 2510.155 1144.265 ;
        RECT 2508.190 1143.950 2510.155 1144.250 ;
        RECT 2508.190 1143.940 2508.570 1143.950 ;
        RECT 2509.825 1143.935 2510.155 1143.950 ;
        RECT 2509.825 1104.810 2510.155 1104.825 ;
        RECT 2509.110 1104.640 2509.490 1104.650 ;
        RECT 2509.825 1104.640 2510.370 1104.810 ;
        RECT 2509.110 1104.340 2510.370 1104.640 ;
        RECT 2509.110 1104.330 2509.490 1104.340 ;
        RECT 2509.110 1034.460 2509.490 1034.780 ;
        RECT 2509.150 1034.090 2509.450 1034.460 ;
        RECT 2510.030 1034.090 2510.410 1034.100 ;
        RECT 2509.150 1033.790 2510.410 1034.090 ;
        RECT 2510.030 1033.780 2510.410 1033.790 ;
        RECT 2510.030 938.580 2510.410 938.900 ;
        RECT 2510.070 937.530 2510.370 938.580 ;
        RECT 2510.950 937.530 2511.330 937.540 ;
        RECT 2510.070 937.230 2511.330 937.530 ;
        RECT 2510.950 937.220 2511.330 937.230 ;
        RECT 2509.110 914.410 2509.490 914.420 ;
        RECT 2510.950 914.410 2511.330 914.420 ;
        RECT 2509.110 914.110 2511.330 914.410 ;
        RECT 2509.110 914.100 2509.490 914.110 ;
        RECT 2510.950 914.100 2511.330 914.110 ;
        RECT 1538.305 513.210 1538.635 513.225 ;
        RECT 2488.870 513.210 2489.250 513.220 ;
        RECT 1538.305 512.910 2489.250 513.210 ;
        RECT 1538.305 512.895 1538.635 512.910 ;
        RECT 2488.870 512.900 2489.250 512.910 ;
      LAYER via3 ;
        RECT 2508.220 3008.500 2508.540 3008.820 ;
        RECT 2508.220 2946.620 2508.540 2946.940 ;
        RECT 2509.140 2945.260 2509.460 2945.580 ;
        RECT 2508.220 2898.340 2508.540 2898.660 ;
        RECT 2508.220 2897.660 2508.540 2897.980 ;
        RECT 2508.220 2774.580 2508.540 2774.900 ;
        RECT 2509.140 2773.900 2509.460 2774.220 ;
        RECT 2510.060 2623.620 2510.380 2623.940 ;
        RECT 2509.140 2611.380 2509.460 2611.700 ;
        RECT 2510.060 2538.620 2510.380 2538.940 ;
        RECT 2510.060 2491.020 2510.380 2491.340 ;
        RECT 2508.220 2437.300 2508.540 2437.620 ;
        RECT 2510.060 2437.300 2510.380 2437.620 ;
        RECT 2510.060 2407.380 2510.380 2407.700 ;
        RECT 2510.060 2359.780 2510.380 2360.100 ;
        RECT 2510.060 2359.100 2510.380 2359.420 ;
        RECT 2510.060 2312.860 2510.380 2313.180 ;
        RECT 2508.220 2294.500 2508.540 2294.820 ;
        RECT 2510.060 2263.220 2510.380 2263.540 ;
        RECT 2510.060 2214.260 2510.380 2214.580 ;
        RECT 2510.060 2166.660 2510.380 2166.980 ;
        RECT 2510.060 2142.180 2510.380 2142.500 ;
        RECT 2510.060 2076.900 2510.380 2077.220 ;
        RECT 2510.060 2069.420 2510.380 2069.740 ;
        RECT 2510.060 2021.820 2510.380 2022.140 ;
        RECT 2510.060 1972.860 2510.380 1973.180 ;
        RECT 2510.060 1925.260 2510.380 1925.580 ;
        RECT 2509.140 1804.220 2509.460 1804.540 ;
        RECT 2510.980 1780.420 2511.300 1780.740 ;
        RECT 2510.980 1772.940 2511.300 1773.260 ;
        RECT 2510.980 1725.340 2511.300 1725.660 ;
        RECT 2510.980 1698.140 2511.300 1698.460 ;
        RECT 2510.060 1696.780 2510.380 1697.100 ;
        RECT 2510.060 1676.380 2510.380 1676.700 ;
        RECT 2510.980 1628.780 2511.300 1629.100 ;
        RECT 2509.140 1345.900 2509.460 1346.220 ;
        RECT 2510.060 1345.900 2510.380 1346.220 ;
        RECT 2508.220 1143.940 2508.540 1144.260 ;
        RECT 2509.140 1104.330 2509.460 1104.650 ;
        RECT 2509.140 1034.460 2509.460 1034.780 ;
        RECT 2510.060 1033.780 2510.380 1034.100 ;
        RECT 2510.060 938.580 2510.380 938.900 ;
        RECT 2510.980 937.220 2511.300 937.540 ;
        RECT 2509.140 914.100 2509.460 914.420 ;
        RECT 2510.980 914.100 2511.300 914.420 ;
        RECT 2488.900 512.900 2489.220 513.220 ;
      LAYER met4 ;
        RECT 2508.215 3008.495 2508.545 3008.825 ;
        RECT 2508.230 2946.945 2508.530 3008.495 ;
        RECT 2508.215 2946.615 2508.545 2946.945 ;
        RECT 2509.135 2945.255 2509.465 2945.585 ;
        RECT 2509.150 2939.450 2509.450 2945.255 ;
        RECT 2508.230 2939.150 2509.450 2939.450 ;
        RECT 2508.230 2898.665 2508.530 2939.150 ;
        RECT 2508.215 2898.335 2508.545 2898.665 ;
        RECT 2508.215 2897.655 2508.545 2897.985 ;
        RECT 2508.230 2774.905 2508.530 2897.655 ;
        RECT 2508.215 2774.575 2508.545 2774.905 ;
        RECT 2509.135 2773.895 2509.465 2774.225 ;
        RECT 2509.150 2667.450 2509.450 2773.895 ;
        RECT 2509.150 2667.150 2510.370 2667.450 ;
        RECT 2510.070 2623.945 2510.370 2667.150 ;
        RECT 2510.055 2623.615 2510.385 2623.945 ;
        RECT 2509.135 2611.375 2509.465 2611.705 ;
        RECT 2509.150 2575.650 2509.450 2611.375 ;
        RECT 2509.150 2575.350 2510.370 2575.650 ;
        RECT 2510.070 2538.945 2510.370 2575.350 ;
        RECT 2510.055 2538.615 2510.385 2538.945 ;
        RECT 2510.055 2491.015 2510.385 2491.345 ;
        RECT 2510.070 2490.650 2510.370 2491.015 ;
        RECT 2508.230 2490.350 2510.370 2490.650 ;
        RECT 2508.230 2437.625 2508.530 2490.350 ;
        RECT 2508.215 2437.295 2508.545 2437.625 ;
        RECT 2510.055 2437.295 2510.385 2437.625 ;
        RECT 2510.070 2407.705 2510.370 2437.295 ;
        RECT 2510.055 2407.375 2510.385 2407.705 ;
        RECT 2510.055 2359.775 2510.385 2360.105 ;
        RECT 2510.070 2359.425 2510.370 2359.775 ;
        RECT 2510.055 2359.095 2510.385 2359.425 ;
        RECT 2510.055 2312.855 2510.385 2313.185 ;
        RECT 2510.070 2310.450 2510.370 2312.855 ;
        RECT 2508.230 2310.150 2510.370 2310.450 ;
        RECT 2508.230 2294.825 2508.530 2310.150 ;
        RECT 2508.215 2294.495 2508.545 2294.825 ;
        RECT 2510.055 2263.215 2510.385 2263.545 ;
        RECT 2510.070 2214.585 2510.370 2263.215 ;
        RECT 2510.055 2214.255 2510.385 2214.585 ;
        RECT 2510.055 2166.655 2510.385 2166.985 ;
        RECT 2510.070 2142.505 2510.370 2166.655 ;
        RECT 2510.055 2142.175 2510.385 2142.505 ;
        RECT 2510.055 2076.895 2510.385 2077.225 ;
        RECT 2510.070 2069.745 2510.370 2076.895 ;
        RECT 2510.055 2069.415 2510.385 2069.745 ;
        RECT 2510.055 2021.815 2510.385 2022.145 ;
        RECT 2510.070 1973.185 2510.370 2021.815 ;
        RECT 2510.055 1972.855 2510.385 1973.185 ;
        RECT 2510.055 1925.255 2510.385 1925.585 ;
        RECT 2510.070 1909.250 2510.370 1925.255 ;
        RECT 2509.150 1908.950 2510.370 1909.250 ;
        RECT 2509.150 1804.545 2509.450 1908.950 ;
        RECT 2509.135 1804.215 2509.465 1804.545 ;
        RECT 2510.975 1780.415 2511.305 1780.745 ;
        RECT 2510.990 1773.265 2511.290 1780.415 ;
        RECT 2510.975 1772.935 2511.305 1773.265 ;
        RECT 2510.975 1725.335 2511.305 1725.665 ;
        RECT 2510.990 1698.465 2511.290 1725.335 ;
        RECT 2510.975 1698.135 2511.305 1698.465 ;
        RECT 2510.055 1696.775 2510.385 1697.105 ;
        RECT 2510.070 1676.705 2510.370 1696.775 ;
        RECT 2510.055 1676.375 2510.385 1676.705 ;
        RECT 2510.975 1628.775 2511.305 1629.105 ;
        RECT 2510.990 1599.850 2511.290 1628.775 ;
        RECT 2510.070 1599.550 2511.290 1599.850 ;
        RECT 2510.070 1489.690 2510.370 1599.550 ;
        RECT 2510.070 1489.390 2511.290 1489.690 ;
        RECT 2510.990 1460.450 2511.290 1489.390 ;
        RECT 2509.150 1460.150 2511.290 1460.450 ;
        RECT 2509.150 1346.225 2509.450 1460.150 ;
        RECT 2509.135 1345.895 2509.465 1346.225 ;
        RECT 2510.055 1345.895 2510.385 1346.225 ;
        RECT 2510.070 1276.850 2510.370 1345.895 ;
        RECT 2508.230 1276.550 2510.370 1276.850 ;
        RECT 2508.230 1144.265 2508.530 1276.550 ;
        RECT 2508.215 1143.935 2508.545 1144.265 ;
        RECT 2509.135 1104.325 2509.465 1104.655 ;
        RECT 2509.150 1034.785 2509.450 1104.325 ;
        RECT 2509.135 1034.455 2509.465 1034.785 ;
        RECT 2510.055 1033.775 2510.385 1034.105 ;
        RECT 2510.070 938.905 2510.370 1033.775 ;
        RECT 2510.055 938.575 2510.385 938.905 ;
        RECT 2510.975 937.215 2511.305 937.545 ;
        RECT 2510.990 914.425 2511.290 937.215 ;
        RECT 2509.135 914.095 2509.465 914.425 ;
        RECT 2510.975 914.095 2511.305 914.425 ;
        RECT 2509.150 729.450 2509.450 914.095 ;
        RECT 2509.150 729.150 2510.370 729.450 ;
        RECT 2510.070 685.690 2510.370 729.150 ;
        RECT 2488.470 684.510 2489.650 685.690 ;
        RECT 2509.630 684.510 2510.810 685.690 ;
        RECT 2488.910 513.225 2489.210 684.510 ;
        RECT 2488.895 512.895 2489.225 513.225 ;
      LAYER met5 ;
        RECT 2488.260 684.300 2511.020 685.900 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.570 496.980 1437.890 497.040 ;
        RECT 1441.710 496.980 1442.030 497.040 ;
        RECT 1437.570 496.840 1442.030 496.980 ;
        RECT 1437.570 496.780 1437.890 496.840 ;
        RECT 1441.710 496.780 1442.030 496.840 ;
        RECT 1441.710 75.040 1442.030 75.100 ;
        RECT 1552.570 75.040 1552.890 75.100 ;
        RECT 1441.710 74.900 1552.890 75.040 ;
        RECT 1441.710 74.840 1442.030 74.900 ;
        RECT 1552.570 74.840 1552.890 74.900 ;
      LAYER via ;
        RECT 1437.600 496.780 1437.860 497.040 ;
        RECT 1441.740 496.780 1442.000 497.040 ;
        RECT 1441.740 74.840 1442.000 75.100 ;
        RECT 1552.600 74.840 1552.860 75.100 ;
      LAYER met2 ;
        RECT 1437.730 510.340 1438.010 514.000 ;
        RECT 1437.660 510.000 1438.010 510.340 ;
        RECT 1437.660 497.070 1437.800 510.000 ;
        RECT 1437.600 496.750 1437.860 497.070 ;
        RECT 1441.740 496.750 1442.000 497.070 ;
        RECT 1441.800 75.130 1441.940 496.750 ;
        RECT 1441.740 74.810 1442.000 75.130 ;
        RECT 1552.600 74.810 1552.860 75.130 ;
        RECT 1552.660 17.410 1552.800 74.810 ;
        RECT 1552.660 17.270 1555.100 17.410 ;
        RECT 1554.960 2.400 1555.100 17.270 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2035.820 2519.810 2035.880 ;
        RECT 2541.110 2035.820 2541.430 2035.880 ;
        RECT 2519.490 2035.680 2541.430 2035.820 ;
        RECT 2519.490 2035.620 2519.810 2035.680 ;
        RECT 2541.110 2035.620 2541.430 2035.680 ;
        RECT 1572.810 424.220 1573.130 424.280 ;
        RECT 2541.110 424.220 2541.430 424.280 ;
        RECT 1572.810 424.080 2541.430 424.220 ;
        RECT 1572.810 424.020 1573.130 424.080 ;
        RECT 2541.110 424.020 2541.430 424.080 ;
      LAYER via ;
        RECT 2519.520 2035.620 2519.780 2035.880 ;
        RECT 2541.140 2035.620 2541.400 2035.880 ;
        RECT 1572.840 424.020 1573.100 424.280 ;
        RECT 2541.140 424.020 2541.400 424.280 ;
      LAYER met2 ;
        RECT 2519.510 2037.435 2519.790 2037.805 ;
        RECT 2519.580 2035.910 2519.720 2037.435 ;
        RECT 2519.520 2035.590 2519.780 2035.910 ;
        RECT 2541.140 2035.590 2541.400 2035.910 ;
        RECT 2541.200 424.310 2541.340 2035.590 ;
        RECT 1572.840 423.990 1573.100 424.310 ;
        RECT 2541.140 423.990 2541.400 424.310 ;
        RECT 1572.900 2.400 1573.040 423.990 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2037.480 2519.790 2037.760 ;
      LAYER met3 ;
        RECT 2506.000 2037.770 2510.000 2037.920 ;
        RECT 2519.485 2037.770 2519.815 2037.785 ;
        RECT 2506.000 2037.470 2519.815 2037.770 ;
        RECT 2506.000 2037.320 2510.000 2037.470 ;
        RECT 2519.485 2037.455 2519.815 2037.470 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 3036.780 338.030 3036.840 ;
        RECT 777.930 3036.780 778.250 3036.840 ;
        RECT 337.710 3036.640 778.250 3036.780 ;
        RECT 337.710 3036.580 338.030 3036.640 ;
        RECT 777.930 3036.580 778.250 3036.640 ;
        RECT 337.710 32.200 338.030 32.260 ;
        RECT 1590.290 32.200 1590.610 32.260 ;
        RECT 337.710 32.060 1590.610 32.200 ;
        RECT 337.710 32.000 338.030 32.060 ;
        RECT 1590.290 32.000 1590.610 32.060 ;
      LAYER via ;
        RECT 337.740 3036.580 338.000 3036.840 ;
        RECT 777.960 3036.580 778.220 3036.840 ;
        RECT 337.740 32.000 338.000 32.260 ;
        RECT 1590.320 32.000 1590.580 32.260 ;
      LAYER met2 ;
        RECT 337.740 3036.550 338.000 3036.870 ;
        RECT 777.960 3036.550 778.220 3036.870 ;
        RECT 337.800 32.290 337.940 3036.550 ;
        RECT 778.020 3010.000 778.160 3036.550 ;
        RECT 778.020 3009.340 778.370 3010.000 ;
        RECT 778.090 3006.000 778.370 3009.340 ;
        RECT 337.740 31.970 338.000 32.290 ;
        RECT 1590.320 31.970 1590.580 32.290 ;
        RECT 1590.380 2.400 1590.520 31.970 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1608.230 17.920 1608.550 17.980 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1608.230 17.780 1614.530 17.920 ;
        RECT 1608.230 17.720 1608.550 17.780 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
      LAYER via ;
        RECT 1608.260 17.720 1608.520 17.980 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
      LAYER met2 ;
        RECT 2457.870 3016.635 2458.150 3017.005 ;
        RECT 2589.430 3016.635 2589.710 3017.005 ;
        RECT 2457.940 3010.000 2458.080 3016.635 ;
        RECT 2457.940 3009.340 2458.290 3010.000 ;
        RECT 2458.010 3006.000 2458.290 3009.340 ;
        RECT 2589.500 508.485 2589.640 3016.635 ;
        RECT 1614.230 508.115 1614.510 508.485 ;
        RECT 2589.430 508.115 2589.710 508.485 ;
        RECT 1614.300 18.010 1614.440 508.115 ;
        RECT 1608.260 17.690 1608.520 18.010 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1608.320 2.400 1608.460 17.690 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
      LAYER via2 ;
        RECT 2457.870 3016.680 2458.150 3016.960 ;
        RECT 2589.430 3016.680 2589.710 3016.960 ;
        RECT 1614.230 508.160 1614.510 508.440 ;
        RECT 2589.430 508.160 2589.710 508.440 ;
      LAYER met3 ;
        RECT 2457.845 3016.970 2458.175 3016.985 ;
        RECT 2589.405 3016.970 2589.735 3016.985 ;
        RECT 2457.845 3016.670 2589.735 3016.970 ;
        RECT 2457.845 3016.655 2458.175 3016.670 ;
        RECT 2589.405 3016.655 2589.735 3016.670 ;
        RECT 1614.205 508.450 1614.535 508.465 ;
        RECT 2589.405 508.450 2589.735 508.465 ;
        RECT 1614.205 508.150 2589.735 508.450 ;
        RECT 1614.205 508.135 1614.535 508.150 ;
        RECT 2589.405 508.135 2589.735 508.150 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 710.845 3029.995 711.015 3030.675 ;
        RECT 711.765 3029.995 711.935 3030.675 ;
        RECT 710.845 3029.825 711.935 3029.995 ;
        RECT 717.745 3018.265 717.915 3030.675 ;
      LAYER mcon ;
        RECT 710.845 3030.505 711.015 3030.675 ;
        RECT 711.765 3030.505 711.935 3030.675 ;
        RECT 717.745 3030.505 717.915 3030.675 ;
      LAYER met1 ;
        RECT 410.390 3030.660 410.710 3030.720 ;
        RECT 710.785 3030.660 711.075 3030.705 ;
        RECT 410.390 3030.520 711.075 3030.660 ;
        RECT 410.390 3030.460 410.710 3030.520 ;
        RECT 710.785 3030.475 711.075 3030.520 ;
        RECT 711.705 3030.660 711.995 3030.705 ;
        RECT 717.685 3030.660 717.975 3030.705 ;
        RECT 711.705 3030.520 717.975 3030.660 ;
        RECT 711.705 3030.475 711.995 3030.520 ;
        RECT 717.685 3030.475 717.975 3030.520 ;
        RECT 717.685 3018.420 717.975 3018.465 ;
        RECT 740.210 3018.420 740.530 3018.480 ;
        RECT 717.685 3018.280 740.530 3018.420 ;
        RECT 717.685 3018.235 717.975 3018.280 ;
        RECT 740.210 3018.220 740.530 3018.280 ;
      LAYER via ;
        RECT 410.420 3030.460 410.680 3030.720 ;
        RECT 740.240 3018.220 740.500 3018.480 ;
      LAYER met2 ;
        RECT 410.420 3030.430 410.680 3030.750 ;
        RECT 410.480 776.405 410.620 3030.430 ;
        RECT 740.240 3018.190 740.500 3018.510 ;
        RECT 740.300 3010.000 740.440 3018.190 ;
        RECT 740.300 3009.340 740.650 3010.000 ;
        RECT 740.370 3006.000 740.650 3009.340 ;
        RECT 410.410 776.035 410.690 776.405 ;
        RECT 1626.190 31.435 1626.470 31.805 ;
        RECT 1626.260 2.400 1626.400 31.435 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
      LAYER via2 ;
        RECT 410.410 776.080 410.690 776.360 ;
        RECT 1626.190 31.480 1626.470 31.760 ;
      LAYER met3 ;
        RECT 360.910 776.370 361.290 776.380 ;
        RECT 410.385 776.370 410.715 776.385 ;
        RECT 360.910 776.070 410.715 776.370 ;
        RECT 360.910 776.060 361.290 776.070 ;
        RECT 410.385 776.055 410.715 776.070 ;
        RECT 360.910 31.770 361.290 31.780 ;
        RECT 1626.165 31.770 1626.495 31.785 ;
        RECT 360.910 31.470 1626.495 31.770 ;
        RECT 360.910 31.460 361.290 31.470 ;
        RECT 1626.165 31.455 1626.495 31.470 ;
      LAYER via3 ;
        RECT 360.940 776.060 361.260 776.380 ;
        RECT 360.940 31.460 361.260 31.780 ;
      LAYER met4 ;
        RECT 360.935 776.055 361.265 776.385 ;
        RECT 360.950 31.785 361.250 776.055 ;
        RECT 360.935 31.455 361.265 31.785 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.970 3024.200 1939.290 3024.260 ;
        RECT 2582.050 3024.200 2582.370 3024.260 ;
        RECT 1938.970 3024.060 2582.370 3024.200 ;
        RECT 1938.970 3024.000 1939.290 3024.060 ;
        RECT 2582.050 3024.000 2582.370 3024.060 ;
        RECT 1648.710 486.440 1649.030 486.500 ;
        RECT 2582.050 486.440 2582.370 486.500 ;
        RECT 1648.710 486.300 2582.370 486.440 ;
        RECT 1648.710 486.240 1649.030 486.300 ;
        RECT 2582.050 486.240 2582.370 486.300 ;
        RECT 1644.110 15.880 1644.430 15.940 ;
        RECT 1648.710 15.880 1649.030 15.940 ;
        RECT 1644.110 15.740 1649.030 15.880 ;
        RECT 1644.110 15.680 1644.430 15.740 ;
        RECT 1648.710 15.680 1649.030 15.740 ;
      LAYER via ;
        RECT 1939.000 3024.000 1939.260 3024.260 ;
        RECT 2582.080 3024.000 2582.340 3024.260 ;
        RECT 1648.740 486.240 1649.000 486.500 ;
        RECT 2582.080 486.240 2582.340 486.500 ;
        RECT 1644.140 15.680 1644.400 15.940 ;
        RECT 1648.740 15.680 1649.000 15.940 ;
      LAYER met2 ;
        RECT 1939.000 3023.970 1939.260 3024.290 ;
        RECT 2582.080 3023.970 2582.340 3024.290 ;
        RECT 1939.060 3010.000 1939.200 3023.970 ;
        RECT 1939.060 3009.340 1939.410 3010.000 ;
        RECT 1939.130 3006.000 1939.410 3009.340 ;
        RECT 2582.140 486.530 2582.280 3023.970 ;
        RECT 1648.740 486.210 1649.000 486.530 ;
        RECT 2582.080 486.210 2582.340 486.530 ;
        RECT 1648.800 15.970 1648.940 486.210 ;
        RECT 1644.140 15.650 1644.400 15.970 ;
        RECT 1648.740 15.650 1649.000 15.970 ;
        RECT 1644.200 2.400 1644.340 15.650 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1656.070 38.320 1656.390 38.380 ;
        RECT 1662.050 38.320 1662.370 38.380 ;
        RECT 1656.070 38.180 1662.370 38.320 ;
        RECT 1656.070 38.120 1656.390 38.180 ;
        RECT 1662.050 38.120 1662.370 38.180 ;
      LAYER via ;
        RECT 1656.100 38.120 1656.360 38.380 ;
        RECT 1662.080 38.120 1662.340 38.380 ;
      LAYER met2 ;
        RECT 1656.090 493.835 1656.370 494.205 ;
        RECT 1656.160 38.410 1656.300 493.835 ;
        RECT 1656.100 38.090 1656.360 38.410 ;
        RECT 1662.080 38.090 1662.340 38.410 ;
        RECT 1662.140 2.400 1662.280 38.090 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
      LAYER via2 ;
        RECT 1656.090 493.880 1656.370 494.160 ;
      LAYER met3 ;
        RECT 407.830 2577.690 408.210 2577.700 ;
        RECT 410.000 2577.690 414.000 2577.840 ;
        RECT 407.830 2577.390 414.000 2577.690 ;
        RECT 407.830 2577.380 408.210 2577.390 ;
        RECT 410.000 2577.240 414.000 2577.390 ;
        RECT 407.830 494.170 408.210 494.180 ;
        RECT 1656.065 494.170 1656.395 494.185 ;
        RECT 407.830 493.870 1656.395 494.170 ;
        RECT 407.830 493.860 408.210 493.870 ;
        RECT 1656.065 493.855 1656.395 493.870 ;
      LAYER via3 ;
        RECT 407.860 2577.380 408.180 2577.700 ;
        RECT 407.860 493.860 408.180 494.180 ;
      LAYER met4 ;
        RECT 407.855 2577.375 408.185 2577.705 ;
        RECT 407.870 494.185 408.170 2577.375 ;
        RECT 407.855 493.855 408.185 494.185 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 1621.700 383.570 1621.760 ;
        RECT 393.370 1621.700 393.690 1621.760 ;
        RECT 383.250 1621.560 393.690 1621.700 ;
        RECT 383.250 1621.500 383.570 1621.560 ;
        RECT 393.370 1621.500 393.690 1621.560 ;
        RECT 383.250 451.760 383.570 451.820 ;
        RECT 1676.770 451.760 1677.090 451.820 ;
        RECT 383.250 451.620 1677.090 451.760 ;
        RECT 383.250 451.560 383.570 451.620 ;
        RECT 1676.770 451.560 1677.090 451.620 ;
        RECT 1676.770 62.120 1677.090 62.180 ;
        RECT 1679.530 62.120 1679.850 62.180 ;
        RECT 1676.770 61.980 1679.850 62.120 ;
        RECT 1676.770 61.920 1677.090 61.980 ;
        RECT 1679.530 61.920 1679.850 61.980 ;
      LAYER via ;
        RECT 383.280 1621.500 383.540 1621.760 ;
        RECT 393.400 1621.500 393.660 1621.760 ;
        RECT 383.280 451.560 383.540 451.820 ;
        RECT 1676.800 451.560 1677.060 451.820 ;
        RECT 1676.800 61.920 1677.060 62.180 ;
        RECT 1679.560 61.920 1679.820 62.180 ;
      LAYER met2 ;
        RECT 393.390 1628.075 393.670 1628.445 ;
        RECT 393.460 1621.790 393.600 1628.075 ;
        RECT 383.280 1621.470 383.540 1621.790 ;
        RECT 393.400 1621.470 393.660 1621.790 ;
        RECT 383.340 451.850 383.480 1621.470 ;
        RECT 383.280 451.530 383.540 451.850 ;
        RECT 1676.800 451.530 1677.060 451.850 ;
        RECT 1676.860 62.210 1677.000 451.530 ;
        RECT 1676.800 61.890 1677.060 62.210 ;
        RECT 1679.560 61.890 1679.820 62.210 ;
        RECT 1679.620 2.400 1679.760 61.890 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
      LAYER via2 ;
        RECT 393.390 1628.120 393.670 1628.400 ;
      LAYER met3 ;
        RECT 393.365 1628.410 393.695 1628.425 ;
        RECT 410.000 1628.410 414.000 1628.560 ;
        RECT 393.365 1628.110 414.000 1628.410 ;
        RECT 393.365 1628.095 393.695 1628.110 ;
        RECT 410.000 1627.960 414.000 1628.110 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 16.560 1697.790 16.620 ;
        RECT 1703.910 16.560 1704.230 16.620 ;
        RECT 1697.470 16.420 1704.230 16.560 ;
        RECT 1697.470 16.360 1697.790 16.420 ;
        RECT 1703.910 16.360 1704.230 16.420 ;
      LAYER via ;
        RECT 1697.500 16.360 1697.760 16.620 ;
        RECT 1703.940 16.360 1704.200 16.620 ;
      LAYER met2 ;
        RECT 1703.930 285.755 1704.210 286.125 ;
        RECT 1704.000 16.650 1704.140 285.755 ;
        RECT 1697.500 16.330 1697.760 16.650 ;
        RECT 1703.940 16.330 1704.200 16.650 ;
        RECT 1697.560 2.400 1697.700 16.330 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
      LAYER via2 ;
        RECT 1703.930 285.800 1704.210 286.080 ;
      LAYER met3 ;
        RECT 2506.000 2529.640 2510.000 2530.240 ;
        RECT 2507.310 2528.060 2507.610 2529.640 ;
        RECT 2507.270 2527.740 2507.650 2528.060 ;
        RECT 2499.910 511.850 2500.290 511.860 ;
        RECT 2499.910 511.550 2501.170 511.850 ;
        RECT 2499.910 511.540 2500.290 511.550 ;
        RECT 2500.870 511.180 2501.170 511.550 ;
        RECT 2500.830 510.860 2501.210 511.180 ;
        RECT 2500.830 437.050 2501.210 437.060 ;
        RECT 2503.590 437.050 2503.970 437.060 ;
        RECT 2500.830 436.750 2503.970 437.050 ;
        RECT 2500.830 436.740 2501.210 436.750 ;
        RECT 2503.590 436.740 2503.970 436.750 ;
        RECT 1703.905 286.090 1704.235 286.105 ;
        RECT 2501.750 286.090 2502.130 286.100 ;
        RECT 1703.905 285.790 2502.130 286.090 ;
        RECT 1703.905 285.775 1704.235 285.790 ;
        RECT 2501.750 285.780 2502.130 285.790 ;
      LAYER via3 ;
        RECT 2507.300 2527.740 2507.620 2528.060 ;
        RECT 2499.940 511.540 2500.260 511.860 ;
        RECT 2500.860 510.860 2501.180 511.180 ;
        RECT 2500.860 436.740 2501.180 437.060 ;
        RECT 2503.620 436.740 2503.940 437.060 ;
        RECT 2501.780 285.780 2502.100 286.100 ;
      LAYER met4 ;
        RECT 2507.295 2528.050 2507.625 2528.065 ;
        RECT 2503.630 2527.750 2507.625 2528.050 ;
        RECT 2503.630 2511.050 2503.930 2527.750 ;
        RECT 2507.295 2527.735 2507.625 2527.750 ;
        RECT 2501.790 2510.750 2503.930 2511.050 ;
        RECT 2501.790 2487.250 2502.090 2510.750 ;
        RECT 2500.870 2486.950 2502.090 2487.250 ;
        RECT 2500.870 2426.050 2501.170 2486.950 ;
        RECT 2499.950 2425.750 2501.170 2426.050 ;
        RECT 2499.950 2296.850 2500.250 2425.750 ;
        RECT 2499.950 2296.550 2502.090 2296.850 ;
        RECT 2501.790 2150.650 2502.090 2296.550 ;
        RECT 2500.870 2150.350 2502.090 2150.650 ;
        RECT 2500.870 1943.250 2501.170 2150.350 ;
        RECT 2500.870 1942.950 2502.090 1943.250 ;
        RECT 2501.790 1871.850 2502.090 1942.950 ;
        RECT 2499.950 1871.550 2502.090 1871.850 ;
        RECT 2499.950 1800.450 2500.250 1871.550 ;
        RECT 2499.950 1800.150 2501.170 1800.450 ;
        RECT 2500.870 1684.850 2501.170 1800.150 ;
        RECT 2499.030 1684.550 2501.170 1684.850 ;
        RECT 2499.030 1630.450 2499.330 1684.550 ;
        RECT 2499.030 1630.150 2500.250 1630.450 ;
        RECT 2499.950 1586.250 2500.250 1630.150 ;
        RECT 2499.950 1585.950 2502.090 1586.250 ;
        RECT 2501.790 1491.050 2502.090 1585.950 ;
        RECT 2501.790 1490.750 2503.010 1491.050 ;
        RECT 2502.710 1487.650 2503.010 1490.750 ;
        RECT 2501.790 1487.350 2503.010 1487.650 ;
        RECT 2501.790 1392.450 2502.090 1487.350 ;
        RECT 2499.030 1392.150 2502.090 1392.450 ;
        RECT 2499.030 1266.650 2499.330 1392.150 ;
        RECT 2498.110 1266.350 2499.330 1266.650 ;
        RECT 2498.110 1205.450 2498.410 1266.350 ;
        RECT 2498.110 1205.150 2501.170 1205.450 ;
        RECT 2500.870 987.850 2501.170 1205.150 ;
        RECT 2499.030 987.550 2501.170 987.850 ;
        RECT 2499.030 970.850 2499.330 987.550 ;
        RECT 2499.030 970.550 2501.170 970.850 ;
        RECT 2500.870 923.250 2501.170 970.550 ;
        RECT 2499.950 922.950 2501.170 923.250 ;
        RECT 2499.950 855.250 2500.250 922.950 ;
        RECT 2499.030 854.950 2500.250 855.250 ;
        RECT 2499.030 807.650 2499.330 854.950 ;
        RECT 2499.030 807.350 2500.250 807.650 ;
        RECT 2499.950 726.490 2500.250 807.350 ;
        RECT 2499.510 725.310 2500.690 726.490 ;
        RECT 2499.510 711.710 2500.690 712.890 ;
        RECT 2499.950 685.250 2500.250 711.710 ;
        RECT 2499.030 684.950 2500.250 685.250 ;
        RECT 2499.030 671.650 2499.330 684.950 ;
        RECT 2499.030 671.350 2500.250 671.650 ;
        RECT 2499.950 603.650 2500.250 671.350 ;
        RECT 2499.950 603.350 2502.090 603.650 ;
        RECT 2501.790 579.850 2502.090 603.350 ;
        RECT 2500.870 579.550 2502.090 579.850 ;
        RECT 2500.870 562.850 2501.170 579.550 ;
        RECT 2500.870 562.550 2502.090 562.850 ;
        RECT 2501.790 556.050 2502.090 562.550 ;
        RECT 2499.950 555.750 2502.090 556.050 ;
        RECT 2499.950 511.865 2500.250 555.750 ;
        RECT 2499.935 511.535 2500.265 511.865 ;
        RECT 2500.855 510.855 2501.185 511.185 ;
        RECT 2500.870 437.065 2501.170 510.855 ;
        RECT 2500.855 436.735 2501.185 437.065 ;
        RECT 2503.615 436.735 2503.945 437.065 ;
        RECT 2503.630 338.450 2503.930 436.735 ;
        RECT 2502.710 338.150 2503.930 338.450 ;
        RECT 2502.710 335.050 2503.010 338.150 ;
        RECT 2501.790 334.750 2503.010 335.050 ;
        RECT 2501.790 286.105 2502.090 334.750 ;
        RECT 2501.775 285.775 2502.105 286.105 ;
      LAYER met5 ;
        RECT 2499.300 723.300 2500.900 726.700 ;
        RECT 2498.380 721.700 2500.900 723.300 ;
        RECT 2498.380 713.100 2499.980 721.700 ;
        RECT 2498.380 711.500 2500.900 713.100 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 357.030 495.280 357.350 495.340 ;
        RECT 731.470 495.280 731.790 495.340 ;
        RECT 357.030 495.140 731.790 495.280 ;
        RECT 357.030 495.080 357.350 495.140 ;
        RECT 731.470 495.080 731.790 495.140 ;
        RECT 731.470 20.300 731.790 20.360 ;
        RECT 734.230 20.300 734.550 20.360 ;
        RECT 731.470 20.160 734.550 20.300 ;
        RECT 731.470 20.100 731.790 20.160 ;
        RECT 734.230 20.100 734.550 20.160 ;
      LAYER via ;
        RECT 357.060 495.080 357.320 495.340 ;
        RECT 731.500 495.080 731.760 495.340 ;
        RECT 731.500 20.100 731.760 20.360 ;
        RECT 734.260 20.100 734.520 20.360 ;
      LAYER met2 ;
        RECT 814.290 3006.690 814.570 3006.805 ;
        RECT 814.890 3006.690 815.170 3010.000 ;
        RECT 814.290 3006.550 815.170 3006.690 ;
        RECT 814.290 3006.435 814.570 3006.550 ;
        RECT 814.890 3006.000 815.170 3006.550 ;
        RECT 357.050 2999.635 357.330 3000.005 ;
        RECT 357.120 495.370 357.260 2999.635 ;
        RECT 357.060 495.050 357.320 495.370 ;
        RECT 731.500 495.050 731.760 495.370 ;
        RECT 731.560 20.390 731.700 495.050 ;
        RECT 731.500 20.070 731.760 20.390 ;
        RECT 734.260 20.070 734.520 20.390 ;
        RECT 734.320 2.400 734.460 20.070 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 814.290 3006.480 814.570 3006.760 ;
        RECT 357.050 2999.680 357.330 2999.960 ;
      LAYER met3 ;
        RECT 814.265 3006.780 814.595 3006.785 ;
        RECT 814.265 3006.770 814.850 3006.780 ;
        RECT 814.265 3006.470 815.050 3006.770 ;
        RECT 814.265 3006.460 814.850 3006.470 ;
        RECT 814.265 3006.455 814.595 3006.460 ;
        RECT 357.025 2999.970 357.355 2999.985 ;
        RECT 814.470 2999.970 814.850 2999.980 ;
        RECT 357.025 2999.670 814.850 2999.970 ;
        RECT 357.025 2999.655 357.355 2999.670 ;
        RECT 814.470 2999.660 814.850 2999.670 ;
      LAYER via3 ;
        RECT 814.500 3006.460 814.820 3006.780 ;
        RECT 814.500 2999.660 814.820 2999.980 ;
      LAYER met4 ;
        RECT 814.495 3006.455 814.825 3006.785 ;
        RECT 814.510 2999.985 814.810 3006.455 ;
        RECT 814.495 2999.655 814.825 2999.985 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 377.270 2594.780 377.590 2594.840 ;
        RECT 394.290 2594.780 394.610 2594.840 ;
        RECT 377.270 2594.640 394.610 2594.780 ;
        RECT 377.270 2594.580 377.590 2594.640 ;
        RECT 394.290 2594.580 394.610 2594.640 ;
        RECT 377.270 431.360 377.590 431.420 ;
        RECT 1711.270 431.360 1711.590 431.420 ;
        RECT 377.270 431.220 1711.590 431.360 ;
        RECT 377.270 431.160 377.590 431.220 ;
        RECT 1711.270 431.160 1711.590 431.220 ;
      LAYER via ;
        RECT 377.300 2594.580 377.560 2594.840 ;
        RECT 394.320 2594.580 394.580 2594.840 ;
        RECT 377.300 431.160 377.560 431.420 ;
        RECT 1711.300 431.160 1711.560 431.420 ;
      LAYER met2 ;
        RECT 394.310 2595.035 394.590 2595.405 ;
        RECT 394.380 2594.870 394.520 2595.035 ;
        RECT 377.300 2594.550 377.560 2594.870 ;
        RECT 394.320 2594.550 394.580 2594.870 ;
        RECT 377.360 431.450 377.500 2594.550 ;
        RECT 377.300 431.130 377.560 431.450 ;
        RECT 1711.300 431.130 1711.560 431.450 ;
        RECT 1711.360 17.410 1711.500 431.130 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
      LAYER via2 ;
        RECT 394.310 2595.080 394.590 2595.360 ;
      LAYER met3 ;
        RECT 394.285 2595.370 394.615 2595.385 ;
        RECT 410.000 2595.370 414.000 2595.520 ;
        RECT 394.285 2595.070 414.000 2595.370 ;
        RECT 394.285 2595.055 394.615 2595.070 ;
        RECT 410.000 2594.920 414.000 2595.070 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.230 3036.355 1407.510 3036.725 ;
        RECT 1407.300 3010.000 1407.440 3036.355 ;
        RECT 1407.300 3009.340 1407.650 3010.000 ;
        RECT 1407.370 3006.000 1407.650 3009.340 ;
        RECT 1733.370 46.395 1733.650 46.765 ;
        RECT 1733.440 2.400 1733.580 46.395 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
      LAYER via2 ;
        RECT 1407.230 3036.400 1407.510 3036.680 ;
        RECT 1733.370 46.440 1733.650 46.720 ;
      LAYER met3 ;
        RECT 1407.205 3036.690 1407.535 3036.705 ;
        RECT 2455.750 3036.690 2456.130 3036.700 ;
        RECT 1407.205 3036.390 2456.130 3036.690 ;
        RECT 1407.205 3036.375 1407.535 3036.390 ;
        RECT 2455.750 3036.380 2456.130 3036.390 ;
        RECT 1733.345 46.730 1733.675 46.745 ;
        RECT 2456.670 46.730 2457.050 46.740 ;
        RECT 1733.345 46.430 2457.050 46.730 ;
        RECT 1733.345 46.415 1733.675 46.430 ;
        RECT 2456.670 46.420 2457.050 46.430 ;
      LAYER via3 ;
        RECT 2455.780 3036.380 2456.100 3036.700 ;
        RECT 2456.700 46.420 2457.020 46.740 ;
      LAYER met4 ;
        RECT 2455.775 3036.375 2456.105 3036.705 ;
        RECT 2455.790 3000.650 2456.090 3036.375 ;
        RECT 2455.790 3000.350 2457.930 3000.650 ;
        RECT 2457.630 2973.450 2457.930 3000.350 ;
        RECT 2457.630 2973.150 2458.850 2973.450 ;
        RECT 2458.550 2919.050 2458.850 2973.150 ;
        RECT 2457.630 2918.750 2458.850 2919.050 ;
        RECT 2457.630 2738.850 2457.930 2918.750 ;
        RECT 2457.630 2738.550 2458.850 2738.850 ;
        RECT 2458.550 2711.650 2458.850 2738.550 ;
        RECT 2456.710 2711.350 2458.850 2711.650 ;
        RECT 2456.710 2664.050 2457.010 2711.350 ;
        RECT 2456.710 2663.750 2458.850 2664.050 ;
        RECT 2458.550 2558.650 2458.850 2663.750 ;
        RECT 2456.710 2558.350 2458.850 2558.650 ;
        RECT 2456.710 2541.650 2457.010 2558.350 ;
        RECT 2456.710 2541.350 2458.850 2541.650 ;
        RECT 2458.550 2429.450 2458.850 2541.350 ;
        RECT 2457.630 2429.150 2458.850 2429.450 ;
        RECT 2457.630 2398.850 2457.930 2429.150 ;
        RECT 2454.870 2398.550 2457.930 2398.850 ;
        RECT 2454.870 2378.450 2455.170 2398.550 ;
        RECT 2454.870 2378.150 2458.850 2378.450 ;
        RECT 2458.550 2235.650 2458.850 2378.150 ;
        RECT 2457.630 2235.350 2458.850 2235.650 ;
        RECT 2457.630 2167.650 2457.930 2235.350 ;
        RECT 2457.630 2167.350 2458.850 2167.650 ;
        RECT 2458.550 2028.250 2458.850 2167.350 ;
        RECT 2456.710 2027.950 2458.850 2028.250 ;
        RECT 2456.710 2021.890 2457.010 2027.950 ;
        RECT 2456.270 2020.710 2457.450 2021.890 ;
        RECT 2460.870 2020.710 2462.050 2021.890 ;
        RECT 2461.310 1936.450 2461.610 2020.710 ;
        RECT 2457.630 1936.150 2461.610 1936.450 ;
        RECT 2457.630 1912.650 2457.930 1936.150 ;
        RECT 2455.790 1912.350 2457.930 1912.650 ;
        RECT 2455.790 1909.250 2456.090 1912.350 ;
        RECT 2454.870 1908.950 2456.090 1909.250 ;
        RECT 2454.870 1854.850 2455.170 1908.950 ;
        RECT 2454.870 1854.550 2456.090 1854.850 ;
        RECT 2455.790 1851.450 2456.090 1854.550 ;
        RECT 2455.790 1851.150 2457.930 1851.450 ;
        RECT 2457.630 1824.250 2457.930 1851.150 ;
        RECT 2457.630 1823.950 2458.850 1824.250 ;
        RECT 2458.550 1572.650 2458.850 1823.950 ;
        RECT 2457.630 1572.350 2458.850 1572.650 ;
        RECT 2457.630 1477.450 2457.930 1572.350 ;
        RECT 2457.630 1477.150 2458.850 1477.450 ;
        RECT 2458.550 1324.450 2458.850 1477.150 ;
        RECT 2457.630 1324.150 2458.850 1324.450 ;
        RECT 2457.630 1270.050 2457.930 1324.150 ;
        RECT 2456.710 1269.750 2457.930 1270.050 ;
        RECT 2456.710 1256.450 2457.010 1269.750 ;
        RECT 2456.710 1256.150 2457.930 1256.450 ;
        RECT 2457.630 1161.690 2457.930 1256.150 ;
        RECT 2440.630 1160.510 2441.810 1161.690 ;
        RECT 2457.190 1160.510 2458.370 1161.690 ;
        RECT 2441.070 940.690 2441.370 1160.510 ;
        RECT 2440.630 939.510 2441.810 940.690 ;
        RECT 2456.270 936.110 2457.450 937.290 ;
        RECT 2456.710 46.745 2457.010 936.110 ;
        RECT 2456.695 46.415 2457.025 46.745 ;
      LAYER met5 ;
        RECT 2456.060 2020.500 2462.260 2022.100 ;
        RECT 2440.420 1160.300 2458.580 1161.900 ;
        RECT 2440.420 937.500 2442.020 940.900 ;
        RECT 2440.420 935.900 2457.660 937.500 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.240 25.940 1666.420 26.080 ;
        RECT 1600.410 25.740 1600.730 25.800 ;
        RECT 1655.240 25.740 1655.380 25.940 ;
        RECT 1600.410 25.600 1655.380 25.740 ;
        RECT 1600.410 25.540 1600.730 25.600 ;
        RECT 1666.280 25.400 1666.420 25.940 ;
        RECT 1751.290 25.400 1751.610 25.460 ;
        RECT 1666.280 25.260 1751.610 25.400 ;
        RECT 1751.290 25.200 1751.610 25.260 ;
      LAYER via ;
        RECT 1600.440 25.540 1600.700 25.800 ;
        RECT 1751.320 25.200 1751.580 25.460 ;
      LAYER met2 ;
        RECT 1598.730 510.410 1599.010 514.000 ;
        RECT 1598.730 510.270 1600.640 510.410 ;
        RECT 1598.730 510.000 1599.010 510.270 ;
        RECT 1600.500 25.830 1600.640 510.270 ;
        RECT 1600.440 25.510 1600.700 25.830 ;
        RECT 1751.320 25.170 1751.580 25.490 ;
        RECT 1751.380 2.400 1751.520 25.170 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1470.060 2520.730 1470.120 ;
        RECT 2561.350 1470.060 2561.670 1470.120 ;
        RECT 2520.410 1469.920 2561.670 1470.060 ;
        RECT 2520.410 1469.860 2520.730 1469.920 ;
        RECT 2561.350 1469.860 2561.670 1469.920 ;
        RECT 1772.910 495.620 1773.230 495.680 ;
        RECT 2561.350 495.620 2561.670 495.680 ;
        RECT 1772.910 495.480 2561.670 495.620 ;
        RECT 1772.910 495.420 1773.230 495.480 ;
        RECT 2561.350 495.420 2561.670 495.480 ;
        RECT 1768.770 15.880 1769.090 15.940 ;
        RECT 1772.910 15.880 1773.230 15.940 ;
        RECT 1768.770 15.740 1773.230 15.880 ;
        RECT 1768.770 15.680 1769.090 15.740 ;
        RECT 1772.910 15.680 1773.230 15.740 ;
      LAYER via ;
        RECT 2520.440 1469.860 2520.700 1470.120 ;
        RECT 2561.380 1469.860 2561.640 1470.120 ;
        RECT 1772.940 495.420 1773.200 495.680 ;
        RECT 2561.380 495.420 2561.640 495.680 ;
        RECT 1768.800 15.680 1769.060 15.940 ;
        RECT 1772.940 15.680 1773.200 15.940 ;
      LAYER met2 ;
        RECT 2520.430 1471.675 2520.710 1472.045 ;
        RECT 2520.500 1470.150 2520.640 1471.675 ;
        RECT 2520.440 1469.830 2520.700 1470.150 ;
        RECT 2561.380 1469.830 2561.640 1470.150 ;
        RECT 2561.440 495.710 2561.580 1469.830 ;
        RECT 1772.940 495.390 1773.200 495.710 ;
        RECT 2561.380 495.390 2561.640 495.710 ;
        RECT 1773.000 15.970 1773.140 495.390 ;
        RECT 1768.800 15.650 1769.060 15.970 ;
        RECT 1772.940 15.650 1773.200 15.970 ;
        RECT 1768.860 2.400 1769.000 15.650 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1471.720 2520.710 1472.000 ;
      LAYER met3 ;
        RECT 2506.000 1472.010 2510.000 1472.160 ;
        RECT 2520.405 1472.010 2520.735 1472.025 ;
        RECT 2506.000 1471.710 2520.735 1472.010 ;
        RECT 2506.000 1471.560 2510.000 1471.710 ;
        RECT 2520.405 1471.695 2520.735 1471.710 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.250 252.180 1786.570 252.240 ;
        RECT 2076.970 252.180 2077.290 252.240 ;
        RECT 1786.250 252.040 2077.290 252.180 ;
        RECT 1786.250 251.980 1786.570 252.040 ;
        RECT 2076.970 251.980 2077.290 252.040 ;
      LAYER via ;
        RECT 1786.280 251.980 1786.540 252.240 ;
        RECT 2077.000 251.980 2077.260 252.240 ;
      LAYER met2 ;
        RECT 2079.890 510.410 2080.170 514.000 ;
        RECT 2077.060 510.270 2080.170 510.410 ;
        RECT 2077.060 252.270 2077.200 510.270 ;
        RECT 2079.890 510.000 2080.170 510.270 ;
        RECT 1786.280 251.950 1786.540 252.270 ;
        RECT 2077.000 251.950 2077.260 252.270 ;
        RECT 1786.340 7.890 1786.480 251.950 ;
        RECT 1786.340 7.750 1786.940 7.890 ;
        RECT 1786.800 2.400 1786.940 7.750 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.690 496.640 919.010 496.700 ;
        RECT 924.210 496.640 924.530 496.700 ;
        RECT 918.690 496.500 924.530 496.640 ;
        RECT 918.690 496.440 919.010 496.500 ;
        RECT 924.210 496.440 924.530 496.500 ;
        RECT 924.210 382.740 924.530 382.800 ;
        RECT 1800.970 382.740 1801.290 382.800 ;
        RECT 924.210 382.600 1801.290 382.740 ;
        RECT 924.210 382.540 924.530 382.600 ;
        RECT 1800.970 382.540 1801.290 382.600 ;
      LAYER via ;
        RECT 918.720 496.440 918.980 496.700 ;
        RECT 924.240 496.440 924.500 496.700 ;
        RECT 924.240 382.540 924.500 382.800 ;
        RECT 1801.000 382.540 1801.260 382.800 ;
      LAYER met2 ;
        RECT 918.850 510.340 919.130 514.000 ;
        RECT 918.780 510.000 919.130 510.340 ;
        RECT 918.780 496.730 918.920 510.000 ;
        RECT 918.720 496.410 918.980 496.730 ;
        RECT 924.240 496.410 924.500 496.730 ;
        RECT 924.300 382.830 924.440 496.410 ;
        RECT 924.240 382.510 924.500 382.830 ;
        RECT 1801.000 382.510 1801.260 382.830 ;
        RECT 1801.060 17.410 1801.200 382.510 ;
        RECT 1801.060 17.270 1804.880 17.410 ;
        RECT 1804.740 2.400 1804.880 17.270 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2284.890 3030.320 2285.210 3030.380 ;
        RECT 2588.950 3030.320 2589.270 3030.380 ;
        RECT 2284.890 3030.180 2589.270 3030.320 ;
        RECT 2284.890 3030.120 2285.210 3030.180 ;
        RECT 2588.950 3030.120 2589.270 3030.180 ;
        RECT 1828.110 487.120 1828.430 487.180 ;
        RECT 2588.950 487.120 2589.270 487.180 ;
        RECT 1828.110 486.980 2589.270 487.120 ;
        RECT 1828.110 486.920 1828.430 486.980 ;
        RECT 2588.950 486.920 2589.270 486.980 ;
        RECT 1822.590 16.900 1822.910 16.960 ;
        RECT 1828.110 16.900 1828.430 16.960 ;
        RECT 1822.590 16.760 1828.430 16.900 ;
        RECT 1822.590 16.700 1822.910 16.760 ;
        RECT 1828.110 16.700 1828.430 16.760 ;
      LAYER via ;
        RECT 2284.920 3030.120 2285.180 3030.380 ;
        RECT 2588.980 3030.120 2589.240 3030.380 ;
        RECT 1828.140 486.920 1828.400 487.180 ;
        RECT 2588.980 486.920 2589.240 487.180 ;
        RECT 1822.620 16.700 1822.880 16.960 ;
        RECT 1828.140 16.700 1828.400 16.960 ;
      LAYER met2 ;
        RECT 2284.920 3030.090 2285.180 3030.410 ;
        RECT 2588.980 3030.090 2589.240 3030.410 ;
        RECT 2284.980 3010.000 2285.120 3030.090 ;
        RECT 2284.980 3009.340 2285.330 3010.000 ;
        RECT 2285.050 3006.000 2285.330 3009.340 ;
        RECT 2589.040 487.210 2589.180 3030.090 ;
        RECT 1828.140 486.890 1828.400 487.210 ;
        RECT 2588.980 486.890 2589.240 487.210 ;
        RECT 1828.200 16.990 1828.340 486.890 ;
        RECT 1822.620 16.670 1822.880 16.990 ;
        RECT 1828.140 16.670 1828.400 16.990 ;
        RECT 1822.680 2.400 1822.820 16.670 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.710 2084.100 384.030 2084.160 ;
        RECT 393.370 2084.100 393.690 2084.160 ;
        RECT 383.710 2083.960 393.690 2084.100 ;
        RECT 383.710 2083.900 384.030 2083.960 ;
        RECT 393.370 2083.900 393.690 2083.960 ;
        RECT 383.710 203.900 384.030 203.960 ;
        RECT 1835.470 203.900 1835.790 203.960 ;
        RECT 383.710 203.760 1835.790 203.900 ;
        RECT 383.710 203.700 384.030 203.760 ;
        RECT 1835.470 203.700 1835.790 203.760 ;
      LAYER via ;
        RECT 383.740 2083.900 384.000 2084.160 ;
        RECT 393.400 2083.900 393.660 2084.160 ;
        RECT 383.740 203.700 384.000 203.960 ;
        RECT 1835.500 203.700 1835.760 203.960 ;
      LAYER met2 ;
        RECT 383.740 2083.870 384.000 2084.190 ;
        RECT 393.400 2084.045 393.660 2084.190 ;
        RECT 383.800 203.990 383.940 2083.870 ;
        RECT 393.390 2083.675 393.670 2084.045 ;
        RECT 383.740 203.670 384.000 203.990 ;
        RECT 1835.500 203.670 1835.760 203.990 ;
        RECT 1835.560 17.410 1835.700 203.670 ;
        RECT 1835.560 17.270 1840.300 17.410 ;
        RECT 1840.160 2.400 1840.300 17.270 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
      LAYER via2 ;
        RECT 393.390 2083.720 393.670 2084.000 ;
      LAYER met3 ;
        RECT 393.365 2084.010 393.695 2084.025 ;
        RECT 410.000 2084.010 414.000 2084.160 ;
        RECT 393.365 2083.710 414.000 2084.010 ;
        RECT 393.365 2083.695 393.695 2083.710 ;
        RECT 410.000 2083.560 414.000 2083.710 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 315.630 1932.120 315.950 1932.180 ;
        RECT 393.370 1932.120 393.690 1932.180 ;
        RECT 315.630 1931.980 393.690 1932.120 ;
        RECT 315.630 1931.920 315.950 1931.980 ;
        RECT 393.370 1931.920 393.690 1931.980 ;
        RECT 315.630 74.360 315.950 74.420 ;
        RECT 1856.170 74.360 1856.490 74.420 ;
        RECT 315.630 74.220 1856.490 74.360 ;
        RECT 315.630 74.160 315.950 74.220 ;
        RECT 1856.170 74.160 1856.490 74.220 ;
      LAYER via ;
        RECT 315.660 1931.920 315.920 1932.180 ;
        RECT 393.400 1931.920 393.660 1932.180 ;
        RECT 315.660 74.160 315.920 74.420 ;
        RECT 1856.200 74.160 1856.460 74.420 ;
      LAYER met2 ;
        RECT 393.390 1938.155 393.670 1938.525 ;
        RECT 393.460 1932.210 393.600 1938.155 ;
        RECT 315.660 1931.890 315.920 1932.210 ;
        RECT 393.400 1931.890 393.660 1932.210 ;
        RECT 315.720 74.450 315.860 1931.890 ;
        RECT 315.660 74.130 315.920 74.450 ;
        RECT 1856.200 74.130 1856.460 74.450 ;
        RECT 1856.260 17.410 1856.400 74.130 ;
        RECT 1856.260 17.270 1858.240 17.410 ;
        RECT 1858.100 2.400 1858.240 17.270 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
      LAYER via2 ;
        RECT 393.390 1938.200 393.670 1938.480 ;
      LAYER met3 ;
        RECT 393.365 1938.490 393.695 1938.505 ;
        RECT 410.000 1938.490 414.000 1938.640 ;
        RECT 393.365 1938.190 414.000 1938.490 ;
        RECT 393.365 1938.175 393.695 1938.190 ;
        RECT 410.000 1938.040 414.000 1938.190 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 19.280 1876.730 19.340 ;
        RECT 2031.890 19.280 2032.210 19.340 ;
        RECT 1876.410 19.140 2032.210 19.280 ;
        RECT 1876.410 19.080 1876.730 19.140 ;
        RECT 2031.890 19.080 2032.210 19.140 ;
      LAYER via ;
        RECT 1876.440 19.080 1876.700 19.340 ;
        RECT 2031.920 19.080 2032.180 19.340 ;
      LAYER met2 ;
        RECT 2521.350 931.075 2521.630 931.445 ;
        RECT 2521.420 926.685 2521.560 931.075 ;
        RECT 2521.350 926.315 2521.630 926.685 ;
        RECT 2520.890 882.795 2521.170 883.165 ;
        RECT 2520.960 877.045 2521.100 882.795 ;
        RECT 2520.890 876.675 2521.170 877.045 ;
        RECT 2031.910 495.195 2032.190 495.565 ;
        RECT 2031.980 19.370 2032.120 495.195 ;
        RECT 1876.440 19.050 1876.700 19.370 ;
        RECT 2031.920 19.050 2032.180 19.370 ;
        RECT 1876.500 9.930 1876.640 19.050 ;
        RECT 1876.040 9.790 1876.640 9.930 ;
        RECT 1876.040 2.400 1876.180 9.790 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
      LAYER via2 ;
        RECT 2521.350 931.120 2521.630 931.400 ;
        RECT 2521.350 926.360 2521.630 926.640 ;
        RECT 2520.890 882.840 2521.170 883.120 ;
        RECT 2520.890 876.720 2521.170 877.000 ;
        RECT 2031.910 495.240 2032.190 495.520 ;
      LAYER met3 ;
        RECT 2506.000 2657.930 2510.000 2658.080 ;
        RECT 2521.070 2657.930 2521.450 2657.940 ;
        RECT 2506.000 2657.630 2521.450 2657.930 ;
        RECT 2506.000 2657.480 2510.000 2657.630 ;
        RECT 2521.070 2657.620 2521.450 2657.630 ;
        RECT 2521.325 931.420 2521.655 931.425 ;
        RECT 2521.070 931.410 2521.655 931.420 ;
        RECT 2521.070 931.110 2521.880 931.410 ;
        RECT 2521.070 931.100 2521.655 931.110 ;
        RECT 2521.325 931.095 2521.655 931.100 ;
        RECT 2521.325 926.660 2521.655 926.665 ;
        RECT 2521.070 926.650 2521.655 926.660 ;
        RECT 2520.870 926.350 2521.655 926.650 ;
        RECT 2521.070 926.340 2521.655 926.350 ;
        RECT 2521.325 926.335 2521.655 926.340 ;
        RECT 2520.865 883.140 2521.195 883.145 ;
        RECT 2520.865 883.130 2521.450 883.140 ;
        RECT 2520.640 882.830 2521.450 883.130 ;
        RECT 2520.865 882.820 2521.450 882.830 ;
        RECT 2520.865 882.815 2521.195 882.820 ;
        RECT 2520.865 877.020 2521.195 877.025 ;
        RECT 2520.865 877.010 2521.450 877.020 ;
        RECT 2520.640 876.710 2521.450 877.010 ;
        RECT 2520.865 876.700 2521.450 876.710 ;
        RECT 2520.865 876.695 2521.195 876.700 ;
        RECT 2031.885 495.530 2032.215 495.545 ;
        RECT 2521.070 495.530 2521.450 495.540 ;
        RECT 2031.885 495.230 2521.450 495.530 ;
        RECT 2031.885 495.215 2032.215 495.230 ;
        RECT 2521.070 495.220 2521.450 495.230 ;
      LAYER via3 ;
        RECT 2521.100 2657.620 2521.420 2657.940 ;
        RECT 2521.100 931.100 2521.420 931.420 ;
        RECT 2521.100 926.340 2521.420 926.660 ;
        RECT 2521.100 882.820 2521.420 883.140 ;
        RECT 2521.100 876.700 2521.420 877.020 ;
        RECT 2521.100 495.220 2521.420 495.540 ;
      LAYER met4 ;
        RECT 2521.095 2657.615 2521.425 2657.945 ;
        RECT 2521.110 931.425 2521.410 2657.615 ;
        RECT 2521.095 931.095 2521.425 931.425 ;
        RECT 2521.095 926.335 2521.425 926.665 ;
        RECT 2521.110 883.145 2521.410 926.335 ;
        RECT 2521.095 882.815 2521.425 883.145 ;
        RECT 2521.095 876.695 2521.425 877.025 ;
        RECT 2521.110 495.545 2521.410 876.695 ;
        RECT 2521.095 495.215 2521.425 495.545 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 349.670 1187.180 349.990 1187.240 ;
        RECT 393.370 1187.180 393.690 1187.240 ;
        RECT 349.670 1187.040 393.690 1187.180 ;
        RECT 349.670 1186.980 349.990 1187.040 ;
        RECT 393.370 1186.980 393.690 1187.040 ;
        RECT 349.670 19.960 349.990 20.020 ;
        RECT 752.170 19.960 752.490 20.020 ;
        RECT 349.670 19.820 752.490 19.960 ;
        RECT 349.670 19.760 349.990 19.820 ;
        RECT 752.170 19.760 752.490 19.820 ;
      LAYER via ;
        RECT 349.700 1186.980 349.960 1187.240 ;
        RECT 393.400 1186.980 393.660 1187.240 ;
        RECT 349.700 19.760 349.960 20.020 ;
        RECT 752.200 19.760 752.460 20.020 ;
      LAYER met2 ;
        RECT 393.390 1188.795 393.670 1189.165 ;
        RECT 393.460 1187.270 393.600 1188.795 ;
        RECT 349.700 1186.950 349.960 1187.270 ;
        RECT 393.400 1186.950 393.660 1187.270 ;
        RECT 349.760 20.050 349.900 1186.950 ;
        RECT 349.700 19.730 349.960 20.050 ;
        RECT 752.200 19.730 752.460 20.050 ;
        RECT 752.260 2.400 752.400 19.730 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 393.390 1188.840 393.670 1189.120 ;
      LAYER met3 ;
        RECT 393.365 1189.130 393.695 1189.145 ;
        RECT 410.000 1189.130 414.000 1189.280 ;
        RECT 393.365 1188.830 414.000 1189.130 ;
        RECT 393.365 1188.815 393.695 1188.830 ;
        RECT 410.000 1188.680 414.000 1188.830 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 384.170 2629.120 384.490 2629.180 ;
        RECT 393.370 2629.120 393.690 2629.180 ;
        RECT 384.170 2628.980 393.690 2629.120 ;
        RECT 384.170 2628.920 384.490 2628.980 ;
        RECT 393.370 2628.920 393.690 2628.980 ;
        RECT 384.170 396.680 384.490 396.740 ;
        RECT 1890.670 396.680 1890.990 396.740 ;
        RECT 384.170 396.540 1890.990 396.680 ;
        RECT 384.170 396.480 384.490 396.540 ;
        RECT 1890.670 396.480 1890.990 396.540 ;
      LAYER via ;
        RECT 384.200 2628.920 384.460 2629.180 ;
        RECT 393.400 2628.920 393.660 2629.180 ;
        RECT 384.200 396.480 384.460 396.740 ;
        RECT 1890.700 396.480 1890.960 396.740 ;
      LAYER met2 ;
        RECT 393.390 2631.755 393.670 2632.125 ;
        RECT 393.460 2629.210 393.600 2631.755 ;
        RECT 384.200 2628.890 384.460 2629.210 ;
        RECT 393.400 2628.890 393.660 2629.210 ;
        RECT 384.260 396.770 384.400 2628.890 ;
        RECT 384.200 396.450 384.460 396.770 ;
        RECT 1890.700 396.450 1890.960 396.770 ;
        RECT 1890.760 17.410 1890.900 396.450 ;
        RECT 1890.760 17.270 1894.120 17.410 ;
        RECT 1893.980 2.400 1894.120 17.270 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
      LAYER via2 ;
        RECT 393.390 2631.800 393.670 2632.080 ;
      LAYER met3 ;
        RECT 393.365 2632.090 393.695 2632.105 ;
        RECT 410.000 2632.090 414.000 2632.240 ;
        RECT 393.365 2631.790 414.000 2632.090 ;
        RECT 393.365 2631.775 393.695 2631.790 ;
        RECT 410.000 2631.640 414.000 2631.790 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1864.450 3036.780 1864.770 3036.840 ;
        RECT 2608.270 3036.780 2608.590 3036.840 ;
        RECT 1864.450 3036.640 2608.590 3036.780 ;
        RECT 1864.450 3036.580 1864.770 3036.640 ;
        RECT 2608.270 3036.580 2608.590 3036.640 ;
        RECT 1911.830 44.780 1912.150 44.840 ;
        RECT 2608.270 44.780 2608.590 44.840 ;
        RECT 1911.830 44.640 2608.590 44.780 ;
        RECT 1911.830 44.580 1912.150 44.640 ;
        RECT 2608.270 44.580 2608.590 44.640 ;
      LAYER via ;
        RECT 1864.480 3036.580 1864.740 3036.840 ;
        RECT 2608.300 3036.580 2608.560 3036.840 ;
        RECT 1911.860 44.580 1912.120 44.840 ;
        RECT 2608.300 44.580 2608.560 44.840 ;
      LAYER met2 ;
        RECT 1864.480 3036.550 1864.740 3036.870 ;
        RECT 2608.300 3036.550 2608.560 3036.870 ;
        RECT 1864.540 3010.000 1864.680 3036.550 ;
        RECT 1864.540 3009.340 1864.890 3010.000 ;
        RECT 1864.610 3006.000 1864.890 3009.340 ;
        RECT 2608.360 44.870 2608.500 3036.550 ;
        RECT 1911.860 44.550 1912.120 44.870 ;
        RECT 2608.300 44.550 2608.560 44.870 ;
        RECT 1911.920 2.400 1912.060 44.550 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2223.250 3025.220 2223.570 3025.280 ;
        RECT 2608.730 3025.220 2609.050 3025.280 ;
        RECT 2223.250 3025.080 2609.050 3025.220 ;
        RECT 2223.250 3025.020 2223.570 3025.080 ;
        RECT 2608.730 3025.020 2609.050 3025.080 ;
        RECT 1931.610 468.080 1931.930 468.140 ;
        RECT 2608.730 468.080 2609.050 468.140 ;
        RECT 1931.610 467.940 2609.050 468.080 ;
        RECT 1931.610 467.880 1931.930 467.940 ;
        RECT 2608.730 467.880 2609.050 467.940 ;
        RECT 1929.310 16.900 1929.630 16.960 ;
        RECT 1931.610 16.900 1931.930 16.960 ;
        RECT 1929.310 16.760 1931.930 16.900 ;
        RECT 1929.310 16.700 1929.630 16.760 ;
        RECT 1931.610 16.700 1931.930 16.760 ;
      LAYER via ;
        RECT 2223.280 3025.020 2223.540 3025.280 ;
        RECT 2608.760 3025.020 2609.020 3025.280 ;
        RECT 1931.640 467.880 1931.900 468.140 ;
        RECT 2608.760 467.880 2609.020 468.140 ;
        RECT 1929.340 16.700 1929.600 16.960 ;
        RECT 1931.640 16.700 1931.900 16.960 ;
      LAYER met2 ;
        RECT 2223.280 3024.990 2223.540 3025.310 ;
        RECT 2608.760 3024.990 2609.020 3025.310 ;
        RECT 2223.340 3010.000 2223.480 3024.990 ;
        RECT 2223.340 3009.340 2223.690 3010.000 ;
        RECT 2223.410 3006.000 2223.690 3009.340 ;
        RECT 2608.820 468.170 2608.960 3024.990 ;
        RECT 1931.640 467.850 1931.900 468.170 ;
        RECT 2608.760 467.850 2609.020 468.170 ;
        RECT 1931.700 16.990 1931.840 467.850 ;
        RECT 1929.340 16.670 1929.600 16.990 ;
        RECT 1931.640 16.670 1931.900 16.990 ;
        RECT 1929.400 2.400 1929.540 16.670 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1945.945 48.365 1946.115 96.475 ;
      LAYER mcon ;
        RECT 1945.945 96.305 1946.115 96.475 ;
      LAYER met1 ;
        RECT 1945.870 96.460 1946.190 96.520 ;
        RECT 1945.675 96.320 1946.190 96.460 ;
        RECT 1945.870 96.260 1946.190 96.320 ;
        RECT 1945.885 48.520 1946.175 48.565 ;
        RECT 1947.250 48.520 1947.570 48.580 ;
        RECT 1945.885 48.380 1947.570 48.520 ;
        RECT 1945.885 48.335 1946.175 48.380 ;
        RECT 1947.250 48.320 1947.570 48.380 ;
      LAYER via ;
        RECT 1945.900 96.260 1946.160 96.520 ;
        RECT 1947.280 48.320 1947.540 48.580 ;
      LAYER met2 ;
        RECT 1945.890 265.355 1946.170 265.725 ;
        RECT 1945.960 96.550 1946.100 265.355 ;
        RECT 1945.900 96.230 1946.160 96.550 ;
        RECT 1947.280 48.290 1947.540 48.610 ;
        RECT 1947.340 2.400 1947.480 48.290 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1945.890 265.400 1946.170 265.680 ;
      LAYER met3 ;
        RECT 410.000 2722.760 414.000 2723.360 ;
        RECT 371.030 2719.130 371.410 2719.140 ;
        RECT 410.630 2719.130 410.930 2722.760 ;
        RECT 371.030 2718.830 410.930 2719.130 ;
        RECT 371.030 2718.820 371.410 2718.830 ;
        RECT 371.030 265.690 371.410 265.700 ;
        RECT 1945.865 265.690 1946.195 265.705 ;
        RECT 371.030 265.390 1946.195 265.690 ;
        RECT 371.030 265.380 371.410 265.390 ;
        RECT 1945.865 265.375 1946.195 265.390 ;
      LAYER via3 ;
        RECT 371.060 2718.820 371.380 2719.140 ;
        RECT 371.060 265.380 371.380 265.700 ;
      LAYER met4 ;
        RECT 371.055 2718.815 371.385 2719.145 ;
        RECT 371.070 265.705 371.370 2718.815 ;
        RECT 371.055 265.375 371.385 265.705 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1965.265 2.805 1965.435 14.195 ;
      LAYER mcon ;
        RECT 1965.265 14.025 1965.435 14.195 ;
      LAYER met1 ;
        RECT 1966.110 473.180 1966.430 473.240 ;
        RECT 2527.770 473.180 2528.090 473.240 ;
        RECT 1966.110 473.040 2528.090 473.180 ;
        RECT 1966.110 472.980 1966.430 473.040 ;
        RECT 2527.770 472.980 2528.090 473.040 ;
        RECT 1965.205 14.180 1965.495 14.225 ;
        RECT 1966.110 14.180 1966.430 14.240 ;
        RECT 1965.205 14.040 1966.430 14.180 ;
        RECT 1965.205 13.995 1965.495 14.040 ;
        RECT 1966.110 13.980 1966.430 14.040 ;
        RECT 1965.190 2.960 1965.510 3.020 ;
        RECT 1964.995 2.820 1965.510 2.960 ;
        RECT 1965.190 2.760 1965.510 2.820 ;
      LAYER via ;
        RECT 1966.140 472.980 1966.400 473.240 ;
        RECT 2527.800 472.980 2528.060 473.240 ;
        RECT 1966.140 13.980 1966.400 14.240 ;
        RECT 1965.220 2.760 1965.480 3.020 ;
      LAYER met2 ;
        RECT 2527.790 1270.395 2528.070 1270.765 ;
        RECT 2527.860 473.270 2528.000 1270.395 ;
        RECT 1966.140 472.950 1966.400 473.270 ;
        RECT 2527.800 472.950 2528.060 473.270 ;
        RECT 1966.200 14.270 1966.340 472.950 ;
        RECT 1966.140 13.950 1966.400 14.270 ;
        RECT 1965.220 2.730 1965.480 3.050 ;
        RECT 1965.280 2.400 1965.420 2.730 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 2527.790 1270.440 2528.070 1270.720 ;
      LAYER met3 ;
        RECT 2506.000 1270.730 2510.000 1270.880 ;
        RECT 2527.765 1270.730 2528.095 1270.745 ;
        RECT 2506.000 1270.430 2528.095 1270.730 ;
        RECT 2506.000 1270.280 2510.000 1270.430 ;
        RECT 2527.765 1270.415 2528.095 1270.430 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 410.620 1055.630 410.680 ;
        RECT 1980.370 410.620 1980.690 410.680 ;
        RECT 1055.310 410.480 1980.690 410.620 ;
        RECT 1055.310 410.420 1055.630 410.480 ;
        RECT 1980.370 410.420 1980.690 410.480 ;
        RECT 1980.370 2.960 1980.690 3.020 ;
        RECT 1983.130 2.960 1983.450 3.020 ;
        RECT 1980.370 2.820 1983.450 2.960 ;
        RECT 1980.370 2.760 1980.690 2.820 ;
        RECT 1983.130 2.760 1983.450 2.820 ;
      LAYER via ;
        RECT 1055.340 410.420 1055.600 410.680 ;
        RECT 1980.400 410.420 1980.660 410.680 ;
        RECT 1980.400 2.760 1980.660 3.020 ;
        RECT 1983.160 2.760 1983.420 3.020 ;
      LAYER met2 ;
        RECT 1055.010 511.770 1055.290 514.000 ;
        RECT 1055.010 511.630 1056.000 511.770 ;
        RECT 1055.010 510.000 1055.290 511.630 ;
        RECT 1055.860 483.210 1056.000 511.630 ;
        RECT 1055.400 483.070 1056.000 483.210 ;
        RECT 1055.400 410.710 1055.540 483.070 ;
        RECT 1055.340 410.390 1055.600 410.710 ;
        RECT 1980.400 410.390 1980.660 410.710 ;
        RECT 1980.460 3.050 1980.600 410.390 ;
        RECT 1980.400 2.730 1980.660 3.050 ;
        RECT 1983.160 2.730 1983.420 3.050 ;
        RECT 1983.220 2.400 1983.360 2.730 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1339.130 502.420 1339.450 502.480 ;
        RECT 1345.110 502.420 1345.430 502.480 ;
        RECT 1339.130 502.280 1345.430 502.420 ;
        RECT 1339.130 502.220 1339.450 502.280 ;
        RECT 1345.110 502.220 1345.430 502.280 ;
        RECT 1345.110 114.140 1345.430 114.200 ;
        RECT 2001.070 114.140 2001.390 114.200 ;
        RECT 1345.110 114.000 2001.390 114.140 ;
        RECT 1345.110 113.940 1345.430 114.000 ;
        RECT 2001.070 113.940 2001.390 114.000 ;
      LAYER via ;
        RECT 1339.160 502.220 1339.420 502.480 ;
        RECT 1345.140 502.220 1345.400 502.480 ;
        RECT 1345.140 113.940 1345.400 114.200 ;
        RECT 2001.100 113.940 2001.360 114.200 ;
      LAYER met2 ;
        RECT 1339.290 510.340 1339.570 514.000 ;
        RECT 1339.220 510.000 1339.570 510.340 ;
        RECT 1339.220 502.510 1339.360 510.000 ;
        RECT 1339.160 502.190 1339.420 502.510 ;
        RECT 1345.140 502.190 1345.400 502.510 ;
        RECT 1345.200 114.230 1345.340 502.190 ;
        RECT 1345.140 113.910 1345.400 114.230 ;
        RECT 2001.100 113.910 2001.360 114.230 ;
        RECT 2001.160 2.400 2001.300 113.910 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.370 3016.720 876.690 3016.780 ;
        RECT 1593.970 3016.720 1594.290 3016.780 ;
        RECT 876.370 3016.580 1594.290 3016.720 ;
        RECT 876.370 3016.520 876.690 3016.580 ;
        RECT 1593.970 3016.520 1594.290 3016.580 ;
      LAYER via ;
        RECT 876.400 3016.520 876.660 3016.780 ;
        RECT 1594.000 3016.520 1594.260 3016.780 ;
      LAYER met2 ;
        RECT 876.400 3016.490 876.660 3016.810 ;
        RECT 1594.000 3016.490 1594.260 3016.810 ;
        RECT 876.460 3010.000 876.600 3016.490 ;
        RECT 1594.060 3011.565 1594.200 3016.490 ;
        RECT 1593.990 3011.195 1594.270 3011.565 ;
        RECT 876.460 3009.340 876.810 3010.000 ;
        RECT 876.530 3006.000 876.810 3009.340 ;
        RECT 2018.570 32.115 2018.850 32.485 ;
        RECT 2018.640 2.400 2018.780 32.115 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 1593.990 3011.240 1594.270 3011.520 ;
        RECT 2018.570 32.160 2018.850 32.440 ;
      LAYER met3 ;
        RECT 1593.965 3011.530 1594.295 3011.545 ;
        RECT 2463.110 3011.530 2463.490 3011.540 ;
        RECT 1593.965 3011.230 2463.490 3011.530 ;
        RECT 1593.965 3011.215 1594.295 3011.230 ;
        RECT 2463.110 3011.220 2463.490 3011.230 ;
        RECT 2018.545 32.450 2018.875 32.465 ;
        RECT 2463.110 32.450 2463.490 32.460 ;
        RECT 2018.545 32.150 2463.490 32.450 ;
        RECT 2018.545 32.135 2018.875 32.150 ;
        RECT 2463.110 32.140 2463.490 32.150 ;
      LAYER via3 ;
        RECT 2463.140 3011.220 2463.460 3011.540 ;
        RECT 2463.140 32.140 2463.460 32.460 ;
      LAYER met4 ;
        RECT 2463.135 3011.215 2463.465 3011.545 ;
        RECT 2463.150 32.465 2463.450 3011.215 ;
        RECT 2463.135 32.135 2463.465 32.465 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1493.710 3024.115 1493.990 3024.485 ;
        RECT 1493.780 3010.000 1493.920 3024.115 ;
        RECT 1493.780 3009.340 1494.130 3010.000 ;
        RECT 1493.850 3006.000 1494.130 3009.340 ;
        RECT 2036.510 31.435 2036.790 31.805 ;
        RECT 2036.580 2.400 2036.720 31.435 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
      LAYER via2 ;
        RECT 1493.710 3024.160 1493.990 3024.440 ;
        RECT 2036.510 31.480 2036.790 31.760 ;
      LAYER met3 ;
        RECT 1493.685 3024.450 1494.015 3024.465 ;
        RECT 2459.430 3024.450 2459.810 3024.460 ;
        RECT 1493.685 3024.150 2459.810 3024.450 ;
        RECT 1493.685 3024.135 1494.015 3024.150 ;
        RECT 2459.430 3024.140 2459.810 3024.150 ;
        RECT 2036.485 31.770 2036.815 31.785 ;
        RECT 2484.270 31.770 2484.650 31.780 ;
        RECT 2036.485 31.470 2484.650 31.770 ;
        RECT 2036.485 31.455 2036.815 31.470 ;
        RECT 2484.270 31.460 2484.650 31.470 ;
      LAYER via3 ;
        RECT 2459.460 3024.140 2459.780 3024.460 ;
        RECT 2484.300 31.460 2484.620 31.780 ;
      LAYER met4 ;
        RECT 2459.455 3024.135 2459.785 3024.465 ;
        RECT 2459.470 2551.850 2459.770 3024.135 ;
        RECT 2457.630 2551.550 2459.770 2551.850 ;
        RECT 2457.630 2545.050 2457.930 2551.550 ;
        RECT 2457.630 2544.750 2459.770 2545.050 ;
        RECT 2459.470 2181.250 2459.770 2544.750 ;
        RECT 2459.470 2180.950 2461.610 2181.250 ;
        RECT 2461.310 2174.450 2461.610 2180.950 ;
        RECT 2459.470 2174.150 2461.610 2174.450 ;
        RECT 2459.470 1950.050 2459.770 2174.150 ;
        RECT 2454.870 1949.750 2459.770 1950.050 ;
        RECT 2454.870 1933.490 2455.170 1949.750 ;
        RECT 2454.430 1932.310 2455.610 1933.490 ;
        RECT 2459.030 1932.310 2460.210 1933.490 ;
        RECT 2459.470 940.690 2459.770 1932.310 ;
        RECT 2459.030 939.510 2460.210 940.690 ;
        RECT 2483.870 939.510 2485.050 940.690 ;
        RECT 2484.310 31.785 2484.610 939.510 ;
        RECT 2484.295 31.455 2484.625 31.785 ;
      LAYER met5 ;
        RECT 2454.220 1932.100 2460.420 1933.700 ;
        RECT 2458.820 939.300 2485.260 940.900 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2055.885 434.945 2056.055 468.435 ;
        RECT 2055.885 338.045 2056.055 385.815 ;
        RECT 2055.885 241.485 2056.055 289.595 ;
        RECT 2055.885 48.705 2056.055 96.475 ;
        RECT 2054.505 2.805 2054.675 48.195 ;
      LAYER mcon ;
        RECT 2055.885 468.265 2056.055 468.435 ;
        RECT 2055.885 385.645 2056.055 385.815 ;
        RECT 2055.885 289.425 2056.055 289.595 ;
        RECT 2055.885 96.305 2056.055 96.475 ;
        RECT 2054.505 48.025 2054.675 48.195 ;
      LAYER met1 ;
        RECT 2519.490 2145.980 2519.810 2146.040 ;
        RECT 2610.570 2145.980 2610.890 2146.040 ;
        RECT 2519.490 2145.840 2610.890 2145.980 ;
        RECT 2519.490 2145.780 2519.810 2145.840 ;
        RECT 2610.570 2145.780 2610.890 2145.840 ;
        RECT 2055.825 468.420 2056.115 468.465 ;
        RECT 2610.570 468.420 2610.890 468.480 ;
        RECT 2055.825 468.280 2610.890 468.420 ;
        RECT 2055.825 468.235 2056.115 468.280 ;
        RECT 2610.570 468.220 2610.890 468.280 ;
        RECT 2055.810 435.100 2056.130 435.160 ;
        RECT 2055.615 434.960 2056.130 435.100 ;
        RECT 2055.810 434.900 2056.130 434.960 ;
        RECT 2055.810 385.800 2056.130 385.860 ;
        RECT 2055.615 385.660 2056.130 385.800 ;
        RECT 2055.810 385.600 2056.130 385.660 ;
        RECT 2055.810 338.200 2056.130 338.260 ;
        RECT 2055.615 338.060 2056.130 338.200 ;
        RECT 2055.810 338.000 2056.130 338.060 ;
        RECT 2055.810 289.580 2056.130 289.640 ;
        RECT 2055.615 289.440 2056.130 289.580 ;
        RECT 2055.810 289.380 2056.130 289.440 ;
        RECT 2055.810 241.640 2056.130 241.700 ;
        RECT 2055.615 241.500 2056.130 241.640 ;
        RECT 2055.810 241.440 2056.130 241.500 ;
        RECT 2055.810 144.740 2056.130 144.800 ;
        RECT 2056.730 144.740 2057.050 144.800 ;
        RECT 2055.810 144.600 2057.050 144.740 ;
        RECT 2055.810 144.540 2056.130 144.600 ;
        RECT 2056.730 144.540 2057.050 144.600 ;
        RECT 2055.810 96.460 2056.130 96.520 ;
        RECT 2055.615 96.320 2056.130 96.460 ;
        RECT 2055.810 96.260 2056.130 96.320 ;
        RECT 2055.810 48.860 2056.130 48.920 ;
        RECT 2055.615 48.720 2056.130 48.860 ;
        RECT 2055.810 48.660 2056.130 48.720 ;
        RECT 2054.445 48.180 2054.735 48.225 ;
        RECT 2055.810 48.180 2056.130 48.240 ;
        RECT 2054.445 48.040 2056.130 48.180 ;
        RECT 2054.445 47.995 2054.735 48.040 ;
        RECT 2055.810 47.980 2056.130 48.040 ;
        RECT 2054.430 2.960 2054.750 3.020 ;
        RECT 2054.235 2.820 2054.750 2.960 ;
        RECT 2054.430 2.760 2054.750 2.820 ;
      LAYER via ;
        RECT 2519.520 2145.780 2519.780 2146.040 ;
        RECT 2610.600 2145.780 2610.860 2146.040 ;
        RECT 2610.600 468.220 2610.860 468.480 ;
        RECT 2055.840 434.900 2056.100 435.160 ;
        RECT 2055.840 385.600 2056.100 385.860 ;
        RECT 2055.840 338.000 2056.100 338.260 ;
        RECT 2055.840 289.380 2056.100 289.640 ;
        RECT 2055.840 241.440 2056.100 241.700 ;
        RECT 2055.840 144.540 2056.100 144.800 ;
        RECT 2056.760 144.540 2057.020 144.800 ;
        RECT 2055.840 96.260 2056.100 96.520 ;
        RECT 2055.840 48.660 2056.100 48.920 ;
        RECT 2055.840 47.980 2056.100 48.240 ;
        RECT 2054.460 2.760 2054.720 3.020 ;
      LAYER met2 ;
        RECT 2519.510 2146.235 2519.790 2146.605 ;
        RECT 2519.580 2146.070 2519.720 2146.235 ;
        RECT 2519.520 2145.750 2519.780 2146.070 ;
        RECT 2610.600 2145.750 2610.860 2146.070 ;
        RECT 2610.660 468.510 2610.800 2145.750 ;
        RECT 2610.600 468.190 2610.860 468.510 ;
        RECT 2055.840 434.870 2056.100 435.190 ;
        RECT 2055.900 385.890 2056.040 434.870 ;
        RECT 2055.840 385.570 2056.100 385.890 ;
        RECT 2055.840 337.970 2056.100 338.290 ;
        RECT 2055.900 289.670 2056.040 337.970 ;
        RECT 2055.840 289.350 2056.100 289.670 ;
        RECT 2055.840 241.410 2056.100 241.730 ;
        RECT 2055.900 144.830 2056.040 241.410 ;
        RECT 2055.840 144.510 2056.100 144.830 ;
        RECT 2056.760 144.510 2057.020 144.830 ;
        RECT 2056.820 97.085 2056.960 144.510 ;
        RECT 2055.830 96.715 2056.110 97.085 ;
        RECT 2056.750 96.715 2057.030 97.085 ;
        RECT 2055.900 96.550 2056.040 96.715 ;
        RECT 2055.840 96.230 2056.100 96.550 ;
        RECT 2055.840 48.630 2056.100 48.950 ;
        RECT 2055.900 48.270 2056.040 48.630 ;
        RECT 2055.840 47.950 2056.100 48.270 ;
        RECT 2054.460 2.730 2054.720 3.050 ;
        RECT 2054.520 2.400 2054.660 2.730 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2146.280 2519.790 2146.560 ;
        RECT 2055.830 96.760 2056.110 97.040 ;
        RECT 2056.750 96.760 2057.030 97.040 ;
      LAYER met3 ;
        RECT 2506.000 2146.570 2510.000 2146.720 ;
        RECT 2519.485 2146.570 2519.815 2146.585 ;
        RECT 2506.000 2146.270 2519.815 2146.570 ;
        RECT 2506.000 2146.120 2510.000 2146.270 ;
        RECT 2519.485 2146.255 2519.815 2146.270 ;
        RECT 2055.805 97.050 2056.135 97.065 ;
        RECT 2056.725 97.050 2057.055 97.065 ;
        RECT 2055.805 96.750 2057.055 97.050 ;
        RECT 2055.805 96.735 2056.135 96.750 ;
        RECT 2056.725 96.735 2057.055 96.750 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 414.605 2507.925 414.775 2539.375 ;
        RECT 414.605 2346.085 414.775 2374.815 ;
        RECT 414.605 2208.385 414.775 2242.895 ;
        RECT 414.145 1873.825 414.315 1931.455 ;
        RECT 414.605 1684.105 414.775 1712.495 ;
        RECT 414.605 1472.965 414.775 1497.615 ;
        RECT 414.605 1297.185 414.775 1369.095 ;
        RECT 414.145 1087.065 414.315 1097.775 ;
        RECT 414.145 1037.425 414.315 1049.835 ;
        RECT 414.605 789.905 414.775 976.395 ;
        RECT 414.145 718.505 414.315 726.155 ;
      LAYER mcon ;
        RECT 414.605 2539.205 414.775 2539.375 ;
        RECT 414.605 2374.645 414.775 2374.815 ;
        RECT 414.605 2242.725 414.775 2242.895 ;
        RECT 414.145 1931.285 414.315 1931.455 ;
        RECT 414.605 1712.325 414.775 1712.495 ;
        RECT 414.605 1497.445 414.775 1497.615 ;
        RECT 414.605 1368.925 414.775 1369.095 ;
        RECT 414.145 1097.605 414.315 1097.775 ;
        RECT 414.145 1049.665 414.315 1049.835 ;
        RECT 414.605 976.225 414.775 976.395 ;
        RECT 414.145 725.985 414.315 726.155 ;
      LAYER met1 ;
        RECT 416.370 3025.560 416.690 3025.620 ;
        RECT 728.250 3025.560 728.570 3025.620 ;
        RECT 416.370 3025.420 728.570 3025.560 ;
        RECT 416.370 3025.360 416.690 3025.420 ;
        RECT 728.250 3025.360 728.570 3025.420 ;
        RECT 414.530 2539.360 414.850 2539.420 ;
        RECT 414.335 2539.220 414.850 2539.360 ;
        RECT 414.530 2539.160 414.850 2539.220 ;
        RECT 414.530 2508.080 414.850 2508.140 ;
        RECT 414.335 2507.940 414.850 2508.080 ;
        RECT 414.530 2507.880 414.850 2507.940 ;
        RECT 414.545 2374.800 414.835 2374.845 ;
        RECT 414.990 2374.800 415.310 2374.860 ;
        RECT 414.545 2374.660 415.310 2374.800 ;
        RECT 414.545 2374.615 414.835 2374.660 ;
        RECT 414.990 2374.600 415.310 2374.660 ;
        RECT 414.545 2346.240 414.835 2346.285 ;
        RECT 414.990 2346.240 415.310 2346.300 ;
        RECT 414.545 2346.100 415.310 2346.240 ;
        RECT 414.545 2346.055 414.835 2346.100 ;
        RECT 414.990 2346.040 415.310 2346.100 ;
        RECT 414.530 2242.880 414.850 2242.940 ;
        RECT 414.335 2242.740 414.850 2242.880 ;
        RECT 414.530 2242.680 414.850 2242.740 ;
        RECT 414.530 2208.540 414.850 2208.600 ;
        RECT 414.335 2208.400 414.850 2208.540 ;
        RECT 414.530 2208.340 414.850 2208.400 ;
        RECT 414.070 2201.060 414.390 2201.120 ;
        RECT 414.530 2201.060 414.850 2201.120 ;
        RECT 414.070 2200.920 414.850 2201.060 ;
        RECT 414.070 2200.860 414.390 2200.920 ;
        RECT 414.530 2200.860 414.850 2200.920 ;
        RECT 414.070 2152.780 414.390 2152.840 ;
        RECT 414.990 2152.780 415.310 2152.840 ;
        RECT 414.070 2152.640 415.310 2152.780 ;
        RECT 414.070 2152.580 414.390 2152.640 ;
        RECT 414.990 2152.580 415.310 2152.640 ;
        RECT 414.085 1931.440 414.375 1931.485 ;
        RECT 414.530 1931.440 414.850 1931.500 ;
        RECT 414.085 1931.300 414.850 1931.440 ;
        RECT 414.085 1931.255 414.375 1931.300 ;
        RECT 414.530 1931.240 414.850 1931.300 ;
        RECT 414.070 1873.980 414.390 1874.040 ;
        RECT 413.875 1873.840 414.390 1873.980 ;
        RECT 414.070 1873.780 414.390 1873.840 ;
        RECT 414.530 1712.480 414.850 1712.540 ;
        RECT 414.335 1712.340 414.850 1712.480 ;
        RECT 414.530 1712.280 414.850 1712.340 ;
        RECT 414.530 1684.260 414.850 1684.320 ;
        RECT 414.335 1684.120 414.850 1684.260 ;
        RECT 414.530 1684.060 414.850 1684.120 ;
        RECT 414.070 1594.160 414.390 1594.220 ;
        RECT 414.530 1594.160 414.850 1594.220 ;
        RECT 414.070 1594.020 414.850 1594.160 ;
        RECT 414.070 1593.960 414.390 1594.020 ;
        RECT 414.530 1593.960 414.850 1594.020 ;
        RECT 414.530 1497.600 414.850 1497.660 ;
        RECT 414.335 1497.460 414.850 1497.600 ;
        RECT 414.530 1497.400 414.850 1497.460 ;
        RECT 414.530 1473.120 414.850 1473.180 ;
        RECT 414.335 1472.980 414.850 1473.120 ;
        RECT 414.530 1472.920 414.850 1472.980 ;
        RECT 414.530 1369.080 414.850 1369.140 ;
        RECT 414.335 1368.940 414.850 1369.080 ;
        RECT 414.530 1368.880 414.850 1368.940 ;
        RECT 414.530 1297.340 414.850 1297.400 ;
        RECT 414.335 1297.200 414.850 1297.340 ;
        RECT 414.530 1297.140 414.850 1297.200 ;
        RECT 414.070 1297.000 414.390 1297.060 ;
        RECT 414.070 1296.860 414.760 1297.000 ;
        RECT 414.070 1296.800 414.390 1296.860 ;
        RECT 414.620 1296.040 414.760 1296.860 ;
        RECT 414.530 1295.780 414.850 1296.040 ;
        RECT 414.085 1097.760 414.375 1097.805 ;
        RECT 414.530 1097.760 414.850 1097.820 ;
        RECT 414.085 1097.620 414.850 1097.760 ;
        RECT 414.085 1097.575 414.375 1097.620 ;
        RECT 414.530 1097.560 414.850 1097.620 ;
        RECT 414.085 1087.220 414.375 1087.265 ;
        RECT 414.990 1087.220 415.310 1087.280 ;
        RECT 414.085 1087.080 415.310 1087.220 ;
        RECT 414.085 1087.035 414.375 1087.080 ;
        RECT 414.990 1087.020 415.310 1087.080 ;
        RECT 414.085 1049.820 414.375 1049.865 ;
        RECT 414.530 1049.820 414.850 1049.880 ;
        RECT 414.085 1049.680 414.850 1049.820 ;
        RECT 414.085 1049.635 414.375 1049.680 ;
        RECT 414.530 1049.620 414.850 1049.680 ;
        RECT 414.085 1037.580 414.375 1037.625 ;
        RECT 414.530 1037.580 414.850 1037.640 ;
        RECT 414.085 1037.440 414.850 1037.580 ;
        RECT 414.085 1037.395 414.375 1037.440 ;
        RECT 414.530 1037.380 414.850 1037.440 ;
        RECT 414.530 976.380 414.850 976.440 ;
        RECT 414.335 976.240 414.850 976.380 ;
        RECT 414.530 976.180 414.850 976.240 ;
        RECT 414.530 790.060 414.850 790.120 ;
        RECT 414.335 789.920 414.850 790.060 ;
        RECT 414.530 789.860 414.850 789.920 ;
        RECT 414.085 726.140 414.375 726.185 ;
        RECT 414.530 726.140 414.850 726.200 ;
        RECT 414.085 726.000 414.850 726.140 ;
        RECT 414.085 725.955 414.375 726.000 ;
        RECT 414.530 725.940 414.850 726.000 ;
        RECT 414.085 718.660 414.375 718.705 ;
        RECT 414.530 718.660 414.850 718.720 ;
        RECT 414.085 718.520 414.850 718.660 ;
        RECT 414.085 718.475 414.375 718.520 ;
        RECT 414.530 718.460 414.850 718.520 ;
        RECT 355.650 700.300 355.970 700.360 ;
        RECT 414.530 700.300 414.850 700.360 ;
        RECT 355.650 700.160 414.850 700.300 ;
        RECT 355.650 700.100 355.970 700.160 ;
        RECT 414.530 700.100 414.850 700.160 ;
        RECT 355.650 34.240 355.970 34.300 ;
        RECT 769.650 34.240 769.970 34.300 ;
        RECT 355.650 34.100 769.970 34.240 ;
        RECT 355.650 34.040 355.970 34.100 ;
        RECT 769.650 34.040 769.970 34.100 ;
      LAYER via ;
        RECT 416.400 3025.360 416.660 3025.620 ;
        RECT 728.280 3025.360 728.540 3025.620 ;
        RECT 414.560 2539.160 414.820 2539.420 ;
        RECT 414.560 2507.880 414.820 2508.140 ;
        RECT 415.020 2374.600 415.280 2374.860 ;
        RECT 415.020 2346.040 415.280 2346.300 ;
        RECT 414.560 2242.680 414.820 2242.940 ;
        RECT 414.560 2208.340 414.820 2208.600 ;
        RECT 414.100 2200.860 414.360 2201.120 ;
        RECT 414.560 2200.860 414.820 2201.120 ;
        RECT 414.100 2152.580 414.360 2152.840 ;
        RECT 415.020 2152.580 415.280 2152.840 ;
        RECT 414.560 1931.240 414.820 1931.500 ;
        RECT 414.100 1873.780 414.360 1874.040 ;
        RECT 414.560 1712.280 414.820 1712.540 ;
        RECT 414.560 1684.060 414.820 1684.320 ;
        RECT 414.100 1593.960 414.360 1594.220 ;
        RECT 414.560 1593.960 414.820 1594.220 ;
        RECT 414.560 1497.400 414.820 1497.660 ;
        RECT 414.560 1472.920 414.820 1473.180 ;
        RECT 414.560 1368.880 414.820 1369.140 ;
        RECT 414.560 1297.140 414.820 1297.400 ;
        RECT 414.100 1296.800 414.360 1297.060 ;
        RECT 414.560 1295.780 414.820 1296.040 ;
        RECT 414.560 1097.560 414.820 1097.820 ;
        RECT 415.020 1087.020 415.280 1087.280 ;
        RECT 414.560 1049.620 414.820 1049.880 ;
        RECT 414.560 1037.380 414.820 1037.640 ;
        RECT 414.560 976.180 414.820 976.440 ;
        RECT 414.560 789.860 414.820 790.120 ;
        RECT 414.560 725.940 414.820 726.200 ;
        RECT 414.560 718.460 414.820 718.720 ;
        RECT 355.680 700.100 355.940 700.360 ;
        RECT 414.560 700.100 414.820 700.360 ;
        RECT 355.680 34.040 355.940 34.300 ;
        RECT 769.680 34.040 769.940 34.300 ;
      LAYER met2 ;
        RECT 416.400 3025.330 416.660 3025.650 ;
        RECT 728.280 3025.330 728.540 3025.650 ;
        RECT 416.460 2984.250 416.600 3025.330 ;
        RECT 728.340 3010.000 728.480 3025.330 ;
        RECT 728.340 3009.340 728.690 3010.000 ;
        RECT 728.410 3006.000 728.690 3009.340 ;
        RECT 416.460 2984.110 417.520 2984.250 ;
        RECT 417.380 2959.770 417.520 2984.110 ;
        RECT 416.920 2959.630 417.520 2959.770 ;
        RECT 416.920 2922.370 417.060 2959.630 ;
        RECT 416.460 2922.230 417.060 2922.370 ;
        RECT 416.460 2897.890 416.600 2922.230 ;
        RECT 415.540 2897.750 416.600 2897.890 ;
        RECT 415.540 2849.780 415.680 2897.750 ;
        RECT 415.540 2849.640 417.060 2849.780 ;
        RECT 416.920 2815.610 417.060 2849.640 ;
        RECT 416.460 2815.470 417.060 2815.610 ;
        RECT 416.460 2767.330 416.600 2815.470 ;
        RECT 416.460 2767.190 417.060 2767.330 ;
        RECT 416.920 2719.050 417.060 2767.190 ;
        RECT 416.460 2718.910 417.060 2719.050 ;
        RECT 416.460 2670.770 416.600 2718.910 ;
        RECT 416.460 2670.630 417.060 2670.770 ;
        RECT 416.920 2622.490 417.060 2670.630 ;
        RECT 416.460 2622.350 417.060 2622.490 ;
        RECT 416.460 2574.210 416.600 2622.350 ;
        RECT 416.460 2574.070 417.060 2574.210 ;
        RECT 414.560 2539.360 414.820 2539.450 ;
        RECT 416.920 2539.360 417.060 2574.070 ;
        RECT 414.560 2539.220 417.060 2539.360 ;
        RECT 414.560 2539.130 414.820 2539.220 ;
        RECT 414.560 2507.850 414.820 2508.170 ;
        RECT 414.620 2507.570 414.760 2507.850 ;
        RECT 414.620 2507.430 417.980 2507.570 ;
        RECT 417.840 2442.970 417.980 2507.430 ;
        RECT 417.840 2442.830 418.440 2442.970 ;
        RECT 418.300 2374.970 418.440 2442.830 ;
        RECT 415.080 2374.890 418.440 2374.970 ;
        RECT 415.020 2374.830 418.440 2374.890 ;
        RECT 415.020 2374.570 415.280 2374.830 ;
        RECT 415.020 2346.010 415.280 2346.330 ;
        RECT 415.080 2318.530 415.220 2346.010 ;
        RECT 415.080 2318.390 416.600 2318.530 ;
        RECT 416.460 2294.050 416.600 2318.390 ;
        RECT 416.000 2293.910 416.600 2294.050 ;
        RECT 416.000 2260.050 416.140 2293.910 ;
        RECT 416.000 2259.910 416.600 2260.050 ;
        RECT 414.560 2242.880 414.820 2242.970 ;
        RECT 416.460 2242.880 416.600 2259.910 ;
        RECT 414.560 2242.740 416.600 2242.880 ;
        RECT 414.560 2242.650 414.820 2242.740 ;
        RECT 414.560 2208.310 414.820 2208.630 ;
        RECT 414.620 2201.150 414.760 2208.310 ;
        RECT 414.100 2200.830 414.360 2201.150 ;
        RECT 414.560 2200.830 414.820 2201.150 ;
        RECT 414.160 2159.410 414.300 2200.830 ;
        RECT 414.160 2159.270 415.220 2159.410 ;
        RECT 415.080 2152.870 415.220 2159.270 ;
        RECT 414.100 2152.550 414.360 2152.870 ;
        RECT 415.020 2152.550 415.280 2152.870 ;
        RECT 414.160 2107.050 414.300 2152.550 ;
        RECT 414.160 2106.910 416.600 2107.050 ;
        RECT 416.460 2098.210 416.600 2106.910 ;
        RECT 416.000 2098.070 416.600 2098.210 ;
        RECT 416.000 2092.090 416.140 2098.070 ;
        RECT 416.000 2091.950 416.600 2092.090 ;
        RECT 416.460 2086.650 416.600 2091.950 ;
        RECT 414.620 2086.510 416.600 2086.650 ;
        RECT 414.620 2039.730 414.760 2086.510 ;
        RECT 414.620 2039.590 415.680 2039.730 ;
        RECT 415.540 2028.680 415.680 2039.590 ;
        RECT 415.540 2028.540 416.600 2028.680 ;
        RECT 416.460 2021.370 416.600 2028.540 ;
        RECT 416.000 2021.230 416.600 2021.370 ;
        RECT 416.000 1968.330 416.140 2021.230 ;
        RECT 415.080 1968.190 416.140 1968.330 ;
        RECT 415.080 1966.970 415.220 1968.190 ;
        RECT 415.080 1966.830 415.680 1966.970 ;
        RECT 415.540 1943.170 415.680 1966.830 ;
        RECT 415.540 1943.030 416.600 1943.170 ;
        RECT 416.460 1931.610 416.600 1943.030 ;
        RECT 414.620 1931.530 416.600 1931.610 ;
        RECT 414.560 1931.470 416.600 1931.530 ;
        RECT 414.560 1931.210 414.820 1931.470 ;
        RECT 414.100 1873.810 414.360 1874.070 ;
        RECT 414.100 1873.750 415.220 1873.810 ;
        RECT 414.160 1873.670 415.220 1873.750 ;
        RECT 415.080 1873.130 415.220 1873.670 ;
        RECT 415.080 1872.990 415.680 1873.130 ;
        RECT 415.540 1835.730 415.680 1872.990 ;
        RECT 415.540 1835.590 416.600 1835.730 ;
        RECT 416.460 1834.370 416.600 1835.590 ;
        RECT 415.540 1834.230 416.600 1834.370 ;
        RECT 415.540 1731.690 415.680 1834.230 ;
        RECT 415.540 1731.550 416.140 1731.690 ;
        RECT 416.000 1712.650 416.140 1731.550 ;
        RECT 414.620 1712.570 416.140 1712.650 ;
        RECT 414.560 1712.510 416.140 1712.570 ;
        RECT 414.560 1712.250 414.820 1712.510 ;
        RECT 414.560 1684.090 414.820 1684.350 ;
        RECT 414.560 1684.030 415.220 1684.090 ;
        RECT 414.620 1683.950 415.220 1684.030 ;
        RECT 415.080 1642.610 415.220 1683.950 ;
        RECT 415.080 1642.470 416.600 1642.610 ;
        RECT 416.460 1618.810 416.600 1642.470 ;
        RECT 414.620 1618.670 416.600 1618.810 ;
        RECT 414.620 1594.250 414.760 1618.670 ;
        RECT 414.100 1593.930 414.360 1594.250 ;
        RECT 414.560 1593.930 414.820 1594.250 ;
        RECT 414.160 1546.050 414.300 1593.930 ;
        RECT 414.160 1545.910 416.600 1546.050 ;
        RECT 416.460 1512.050 416.600 1545.910 ;
        RECT 415.080 1511.910 416.600 1512.050 ;
        RECT 414.560 1497.600 414.820 1497.690 ;
        RECT 415.080 1497.600 415.220 1511.910 ;
        RECT 414.560 1497.460 415.220 1497.600 ;
        RECT 414.560 1497.370 414.820 1497.460 ;
        RECT 414.560 1472.890 414.820 1473.210 ;
        RECT 414.620 1471.930 414.760 1472.890 ;
        RECT 414.620 1471.790 417.520 1471.930 ;
        RECT 417.380 1369.250 417.520 1471.790 ;
        RECT 414.620 1369.170 417.520 1369.250 ;
        RECT 414.560 1369.110 417.520 1369.170 ;
        RECT 414.560 1368.850 414.820 1369.110 ;
        RECT 414.620 1297.430 414.760 1297.585 ;
        RECT 414.560 1297.170 414.820 1297.430 ;
        RECT 414.160 1297.110 414.820 1297.170 ;
        RECT 414.160 1297.090 414.760 1297.110 ;
        RECT 414.100 1297.030 414.760 1297.090 ;
        RECT 414.100 1296.770 414.360 1297.030 ;
        RECT 414.560 1295.750 414.820 1296.070 ;
        RECT 414.620 1230.530 414.760 1295.750 ;
        RECT 414.620 1230.390 416.140 1230.530 ;
        RECT 416.000 1160.490 416.140 1230.390 ;
        RECT 416.000 1160.350 416.600 1160.490 ;
        RECT 416.460 1159.810 416.600 1160.350 ;
        RECT 416.460 1159.670 417.520 1159.810 ;
        RECT 417.380 1097.930 417.520 1159.670 ;
        RECT 414.620 1097.850 417.520 1097.930 ;
        RECT 414.560 1097.790 417.520 1097.850 ;
        RECT 414.560 1097.530 414.820 1097.790 ;
        RECT 415.020 1087.050 415.280 1087.310 ;
        RECT 415.020 1086.990 418.440 1087.050 ;
        RECT 415.080 1086.910 418.440 1086.990 ;
        RECT 418.300 1053.730 418.440 1086.910 ;
        RECT 415.540 1053.590 418.440 1053.730 ;
        RECT 415.540 1053.050 415.680 1053.590 ;
        RECT 414.620 1052.910 415.680 1053.050 ;
        RECT 414.620 1049.910 414.760 1052.910 ;
        RECT 414.560 1049.590 414.820 1049.910 ;
        RECT 414.560 1037.350 414.820 1037.670 ;
        RECT 414.620 976.470 414.760 1037.350 ;
        RECT 414.560 976.150 414.820 976.470 ;
        RECT 414.560 789.830 414.820 790.150 ;
        RECT 414.620 776.120 414.760 789.830 ;
        RECT 414.620 775.980 417.980 776.120 ;
        RECT 417.840 745.690 417.980 775.980 ;
        RECT 417.380 745.550 417.980 745.690 ;
        RECT 417.380 743.650 417.520 745.550 ;
        RECT 416.000 743.510 417.520 743.650 ;
        RECT 416.000 740.930 416.140 743.510 ;
        RECT 414.620 740.790 416.140 740.930 ;
        RECT 414.620 726.230 414.760 740.790 ;
        RECT 414.560 725.910 414.820 726.230 ;
        RECT 414.560 718.490 414.820 718.750 ;
        RECT 414.560 718.430 415.680 718.490 ;
        RECT 414.620 718.350 415.680 718.430 ;
        RECT 355.680 700.070 355.940 700.390 ;
        RECT 414.560 700.300 414.820 700.390 ;
        RECT 415.540 700.300 415.680 718.350 ;
        RECT 414.560 700.160 415.680 700.300 ;
        RECT 414.560 700.070 414.820 700.160 ;
        RECT 355.740 34.330 355.880 700.070 ;
        RECT 355.680 34.010 355.940 34.330 ;
        RECT 769.680 34.010 769.940 34.330 ;
        RECT 769.740 2.400 769.880 34.010 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2070.070 96.460 2070.390 96.520 ;
        RECT 2072.370 96.460 2072.690 96.520 ;
        RECT 2070.070 96.320 2072.690 96.460 ;
        RECT 2070.070 96.260 2070.390 96.320 ;
        RECT 2072.370 96.260 2072.690 96.320 ;
      LAYER via ;
        RECT 2070.100 96.260 2070.360 96.520 ;
        RECT 2072.400 96.260 2072.660 96.520 ;
      LAYER met2 ;
        RECT 2049.390 175.595 2049.670 175.965 ;
        RECT 2049.460 146.045 2049.600 175.595 ;
        RECT 2049.390 145.675 2049.670 146.045 ;
        RECT 2070.090 144.995 2070.370 145.365 ;
        RECT 2070.160 96.550 2070.300 144.995 ;
        RECT 2070.100 96.230 2070.360 96.550 ;
        RECT 2072.400 96.230 2072.660 96.550 ;
        RECT 2072.460 2.400 2072.600 96.230 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 2049.390 175.640 2049.670 175.920 ;
        RECT 2049.390 145.720 2049.670 146.000 ;
        RECT 2070.090 145.040 2070.370 145.320 ;
      LAYER met3 ;
        RECT 371.950 2705.530 372.330 2705.540 ;
        RECT 410.000 2705.530 414.000 2705.680 ;
        RECT 371.950 2705.230 414.000 2705.530 ;
        RECT 371.950 2705.220 372.330 2705.230 ;
        RECT 410.000 2705.080 414.000 2705.230 ;
        RECT 371.950 175.930 372.330 175.940 ;
        RECT 2049.365 175.930 2049.695 175.945 ;
        RECT 371.950 175.630 2049.695 175.930 ;
        RECT 371.950 175.620 372.330 175.630 ;
        RECT 2049.365 175.615 2049.695 175.630 ;
        RECT 2049.365 146.010 2049.695 146.025 ;
        RECT 2049.365 145.710 2070.380 146.010 ;
        RECT 2049.365 145.695 2049.695 145.710 ;
        RECT 2070.080 145.345 2070.380 145.710 ;
        RECT 2070.065 145.015 2070.395 145.345 ;
      LAYER via3 ;
        RECT 371.980 2705.220 372.300 2705.540 ;
        RECT 371.980 175.620 372.300 175.940 ;
      LAYER met4 ;
        RECT 371.975 2705.215 372.305 2705.545 ;
        RECT 371.990 175.945 372.290 2705.215 ;
        RECT 371.975 175.615 372.305 175.945 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 322.990 3019.440 323.310 3019.500 ;
        RECT 493.650 3019.440 493.970 3019.500 ;
        RECT 322.990 3019.300 493.970 3019.440 ;
        RECT 322.990 3019.240 323.310 3019.300 ;
        RECT 493.650 3019.240 493.970 3019.300 ;
        RECT 322.990 73.340 323.310 73.400 ;
        RECT 2083.870 73.340 2084.190 73.400 ;
        RECT 322.990 73.200 2084.190 73.340 ;
        RECT 322.990 73.140 323.310 73.200 ;
        RECT 2083.870 73.140 2084.190 73.200 ;
        RECT 2083.870 38.320 2084.190 38.380 ;
        RECT 2089.850 38.320 2090.170 38.380 ;
        RECT 2083.870 38.180 2090.170 38.320 ;
        RECT 2083.870 38.120 2084.190 38.180 ;
        RECT 2089.850 38.120 2090.170 38.180 ;
      LAYER via ;
        RECT 323.020 3019.240 323.280 3019.500 ;
        RECT 493.680 3019.240 493.940 3019.500 ;
        RECT 323.020 73.140 323.280 73.400 ;
        RECT 2083.900 73.140 2084.160 73.400 ;
        RECT 2083.900 38.120 2084.160 38.380 ;
        RECT 2089.880 38.120 2090.140 38.380 ;
      LAYER met2 ;
        RECT 323.020 3019.210 323.280 3019.530 ;
        RECT 493.680 3019.210 493.940 3019.530 ;
        RECT 323.080 73.430 323.220 3019.210 ;
        RECT 493.740 3010.000 493.880 3019.210 ;
        RECT 493.740 3009.340 494.090 3010.000 ;
        RECT 493.810 3006.000 494.090 3009.340 ;
        RECT 323.020 73.110 323.280 73.430 ;
        RECT 2083.900 73.110 2084.160 73.430 ;
        RECT 2083.960 38.410 2084.100 73.110 ;
        RECT 2083.900 38.090 2084.160 38.410 ;
        RECT 2089.880 38.090 2090.140 38.410 ;
        RECT 2089.940 2.400 2090.080 38.090 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2107.790 16.900 2108.110 16.960 ;
        RECT 2111.010 16.900 2111.330 16.960 ;
        RECT 2107.790 16.760 2111.330 16.900 ;
        RECT 2107.790 16.700 2108.110 16.760 ;
        RECT 2111.010 16.700 2111.330 16.760 ;
      LAYER via ;
        RECT 2107.820 16.700 2108.080 16.960 ;
        RECT 2111.040 16.700 2111.300 16.960 ;
      LAYER met2 ;
        RECT 2502.490 438.075 2502.770 438.445 ;
        RECT 2502.560 410.565 2502.700 438.075 ;
        RECT 2111.030 410.195 2111.310 410.565 ;
        RECT 2502.490 410.195 2502.770 410.565 ;
        RECT 2111.100 16.990 2111.240 410.195 ;
        RECT 2107.820 16.670 2108.080 16.990 ;
        RECT 2111.040 16.670 2111.300 16.990 ;
        RECT 2107.880 2.400 2108.020 16.670 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 2502.490 438.120 2502.770 438.400 ;
        RECT 2111.030 410.240 2111.310 410.520 ;
        RECT 2502.490 410.240 2502.770 410.520 ;
      LAYER met3 ;
        RECT 2506.000 995.560 2510.000 996.160 ;
        RECT 2507.310 994.660 2507.610 995.560 ;
        RECT 2507.270 994.340 2507.650 994.660 ;
        RECT 2502.465 438.420 2502.795 438.425 ;
        RECT 2502.465 438.410 2503.050 438.420 ;
        RECT 2502.240 438.110 2503.050 438.410 ;
        RECT 2502.465 438.100 2503.050 438.110 ;
        RECT 2502.465 438.095 2502.795 438.100 ;
        RECT 2111.005 410.530 2111.335 410.545 ;
        RECT 2502.465 410.530 2502.795 410.545 ;
        RECT 2111.005 410.230 2502.795 410.530 ;
        RECT 2111.005 410.215 2111.335 410.230 ;
        RECT 2502.465 410.215 2502.795 410.230 ;
      LAYER via3 ;
        RECT 2507.300 994.340 2507.620 994.660 ;
        RECT 2502.700 438.100 2503.020 438.420 ;
      LAYER met4 ;
        RECT 2507.295 994.650 2507.625 994.665 ;
        RECT 2503.630 994.350 2507.625 994.650 ;
        RECT 2503.630 947.050 2503.930 994.350 ;
        RECT 2507.295 994.335 2507.625 994.350 ;
        RECT 2501.790 946.750 2503.930 947.050 ;
        RECT 2501.790 814.890 2502.090 946.750 ;
        RECT 2501.350 813.710 2502.530 814.890 ;
        RECT 2501.350 806.910 2502.530 808.090 ;
        RECT 2501.790 732.850 2502.090 806.910 ;
        RECT 2501.790 732.550 2503.930 732.850 ;
        RECT 2503.630 624.050 2503.930 732.550 ;
        RECT 2501.790 623.750 2503.930 624.050 ;
        RECT 2501.790 613.850 2502.090 623.750 ;
        RECT 2501.790 613.550 2503.010 613.850 ;
        RECT 2502.710 438.425 2503.010 613.550 ;
        RECT 2502.695 438.095 2503.025 438.425 ;
      LAYER met5 ;
        RECT 2501.140 806.700 2502.740 815.100 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.550 3030.915 1679.830 3031.285 ;
        RECT 1679.620 3010.000 1679.760 3030.915 ;
        RECT 1679.620 3009.340 1679.970 3010.000 ;
        RECT 1679.690 3006.000 1679.970 3009.340 ;
        RECT 2125.750 32.795 2126.030 33.165 ;
        RECT 2125.820 2.400 2125.960 32.795 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
      LAYER via2 ;
        RECT 1679.550 3030.960 1679.830 3031.240 ;
        RECT 2125.750 32.840 2126.030 33.120 ;
      LAYER met3 ;
        RECT 1679.525 3031.250 1679.855 3031.265 ;
        RECT 2539.470 3031.250 2539.850 3031.260 ;
        RECT 1679.525 3030.950 2539.850 3031.250 ;
        RECT 1679.525 3030.935 1679.855 3030.950 ;
        RECT 2539.470 3030.940 2539.850 3030.950 ;
        RECT 2125.725 33.130 2126.055 33.145 ;
        RECT 2539.470 33.130 2539.850 33.140 ;
        RECT 2125.725 32.830 2539.850 33.130 ;
        RECT 2125.725 32.815 2126.055 32.830 ;
        RECT 2539.470 32.820 2539.850 32.830 ;
      LAYER via3 ;
        RECT 2539.500 3030.940 2539.820 3031.260 ;
        RECT 2539.500 32.820 2539.820 33.140 ;
      LAYER met4 ;
        RECT 2539.495 3030.935 2539.825 3031.265 ;
        RECT 2539.510 33.145 2539.810 3030.935 ;
        RECT 2539.495 32.815 2539.825 33.145 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 369.450 1042.000 369.770 1042.060 ;
        RECT 393.370 1042.000 393.690 1042.060 ;
        RECT 369.450 1041.860 393.690 1042.000 ;
        RECT 369.450 1041.800 369.770 1041.860 ;
        RECT 393.370 1041.800 393.690 1041.860 ;
        RECT 369.450 73.000 369.770 73.060 ;
        RECT 2139.070 73.000 2139.390 73.060 ;
        RECT 369.450 72.860 2139.390 73.000 ;
        RECT 369.450 72.800 369.770 72.860 ;
        RECT 2139.070 72.800 2139.390 72.860 ;
      LAYER via ;
        RECT 369.480 1041.800 369.740 1042.060 ;
        RECT 393.400 1041.800 393.660 1042.060 ;
        RECT 369.480 72.800 369.740 73.060 ;
        RECT 2139.100 72.800 2139.360 73.060 ;
      LAYER met2 ;
        RECT 393.390 1043.275 393.670 1043.645 ;
        RECT 393.460 1042.090 393.600 1043.275 ;
        RECT 369.480 1041.770 369.740 1042.090 ;
        RECT 393.400 1041.770 393.660 1042.090 ;
        RECT 369.540 73.090 369.680 1041.770 ;
        RECT 369.480 72.770 369.740 73.090 ;
        RECT 2139.100 72.770 2139.360 73.090 ;
        RECT 2139.160 16.730 2139.300 72.770 ;
        RECT 2139.160 16.590 2143.900 16.730 ;
        RECT 2143.760 2.400 2143.900 16.590 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
      LAYER via2 ;
        RECT 393.390 1043.320 393.670 1043.600 ;
      LAYER met3 ;
        RECT 393.365 1043.610 393.695 1043.625 ;
        RECT 410.000 1043.610 414.000 1043.760 ;
        RECT 393.365 1043.310 414.000 1043.610 ;
        RECT 393.365 1043.295 393.695 1043.310 ;
        RECT 410.000 1043.160 414.000 1043.310 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1304.480 2520.730 1304.540 ;
        RECT 2535.590 1304.480 2535.910 1304.540 ;
        RECT 2520.410 1304.340 2535.910 1304.480 ;
        RECT 2520.410 1304.280 2520.730 1304.340 ;
        RECT 2535.590 1304.280 2535.910 1304.340 ;
        RECT 2166.210 468.760 2166.530 468.820 ;
        RECT 2535.590 468.760 2535.910 468.820 ;
        RECT 2166.210 468.620 2535.910 468.760 ;
        RECT 2166.210 468.560 2166.530 468.620 ;
        RECT 2535.590 468.560 2535.910 468.620 ;
        RECT 2161.610 30.160 2161.930 30.220 ;
        RECT 2166.210 30.160 2166.530 30.220 ;
        RECT 2161.610 30.020 2166.530 30.160 ;
        RECT 2161.610 29.960 2161.930 30.020 ;
        RECT 2166.210 29.960 2166.530 30.020 ;
      LAYER via ;
        RECT 2520.440 1304.280 2520.700 1304.540 ;
        RECT 2535.620 1304.280 2535.880 1304.540 ;
        RECT 2166.240 468.560 2166.500 468.820 ;
        RECT 2535.620 468.560 2535.880 468.820 ;
        RECT 2161.640 29.960 2161.900 30.220 ;
        RECT 2166.240 29.960 2166.500 30.220 ;
      LAYER met2 ;
        RECT 2520.430 1307.115 2520.710 1307.485 ;
        RECT 2520.500 1304.570 2520.640 1307.115 ;
        RECT 2520.440 1304.250 2520.700 1304.570 ;
        RECT 2535.620 1304.250 2535.880 1304.570 ;
        RECT 2535.680 468.850 2535.820 1304.250 ;
        RECT 2166.240 468.530 2166.500 468.850 ;
        RECT 2535.620 468.530 2535.880 468.850 ;
        RECT 2166.300 30.250 2166.440 468.530 ;
        RECT 2161.640 29.930 2161.900 30.250 ;
        RECT 2166.240 29.930 2166.500 30.250 ;
        RECT 2161.700 2.400 2161.840 29.930 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1307.160 2520.710 1307.440 ;
      LAYER met3 ;
        RECT 2506.000 1307.450 2510.000 1307.600 ;
        RECT 2520.405 1307.450 2520.735 1307.465 ;
        RECT 2506.000 1307.150 2520.735 1307.450 ;
        RECT 2506.000 1307.000 2510.000 1307.150 ;
        RECT 2520.405 1307.135 2520.735 1307.150 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2491.080 2519.810 2491.140 ;
        RECT 2539.730 2491.080 2540.050 2491.140 ;
        RECT 2519.490 2490.940 2540.050 2491.080 ;
        RECT 2519.490 2490.880 2519.810 2490.940 ;
        RECT 2539.730 2490.880 2540.050 2490.940 ;
        RECT 2180.010 459.580 2180.330 459.640 ;
        RECT 2539.730 459.580 2540.050 459.640 ;
        RECT 2180.010 459.440 2540.050 459.580 ;
        RECT 2180.010 459.380 2180.330 459.440 ;
        RECT 2539.730 459.380 2540.050 459.440 ;
      LAYER via ;
        RECT 2519.520 2490.880 2519.780 2491.140 ;
        RECT 2539.760 2490.880 2540.020 2491.140 ;
        RECT 2180.040 459.380 2180.300 459.640 ;
        RECT 2539.760 459.380 2540.020 459.640 ;
      LAYER met2 ;
        RECT 2519.510 2494.395 2519.790 2494.765 ;
        RECT 2519.580 2491.170 2519.720 2494.395 ;
        RECT 2519.520 2490.850 2519.780 2491.170 ;
        RECT 2539.760 2490.850 2540.020 2491.170 ;
        RECT 2539.820 459.670 2539.960 2490.850 ;
        RECT 2180.040 459.350 2180.300 459.670 ;
        RECT 2539.760 459.350 2540.020 459.670 ;
        RECT 2180.100 16.730 2180.240 459.350 ;
        RECT 2179.180 16.590 2180.240 16.730 ;
        RECT 2179.180 2.400 2179.320 16.590 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2494.440 2519.790 2494.720 ;
      LAYER met3 ;
        RECT 2506.000 2494.730 2510.000 2494.880 ;
        RECT 2519.485 2494.730 2519.815 2494.745 ;
        RECT 2506.000 2494.430 2519.815 2494.730 ;
        RECT 2506.000 2494.280 2510.000 2494.430 ;
        RECT 2519.485 2494.415 2519.815 2494.430 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.810 3016.720 2470.130 3016.780 ;
        RECT 2581.590 3016.720 2581.910 3016.780 ;
        RECT 2469.810 3016.580 2581.910 3016.720 ;
        RECT 2469.810 3016.520 2470.130 3016.580 ;
        RECT 2581.590 3016.520 2581.910 3016.580 ;
        RECT 2200.710 482.020 2201.030 482.080 ;
        RECT 2581.590 482.020 2581.910 482.080 ;
        RECT 2200.710 481.880 2581.910 482.020 ;
        RECT 2200.710 481.820 2201.030 481.880 ;
        RECT 2581.590 481.820 2581.910 481.880 ;
        RECT 2197.030 16.900 2197.350 16.960 ;
        RECT 2200.710 16.900 2201.030 16.960 ;
        RECT 2197.030 16.760 2201.030 16.900 ;
        RECT 2197.030 16.700 2197.350 16.760 ;
        RECT 2200.710 16.700 2201.030 16.760 ;
      LAYER via ;
        RECT 2469.840 3016.520 2470.100 3016.780 ;
        RECT 2581.620 3016.520 2581.880 3016.780 ;
        RECT 2200.740 481.820 2201.000 482.080 ;
        RECT 2581.620 481.820 2581.880 482.080 ;
        RECT 2197.060 16.700 2197.320 16.960 ;
        RECT 2200.740 16.700 2201.000 16.960 ;
      LAYER met2 ;
        RECT 2469.840 3016.490 2470.100 3016.810 ;
        RECT 2581.620 3016.490 2581.880 3016.810 ;
        RECT 2469.900 3010.000 2470.040 3016.490 ;
        RECT 2469.900 3009.340 2470.250 3010.000 ;
        RECT 2469.970 3006.000 2470.250 3009.340 ;
        RECT 2581.680 482.110 2581.820 3016.490 ;
        RECT 2200.740 481.790 2201.000 482.110 ;
        RECT 2581.620 481.790 2581.880 482.110 ;
        RECT 2200.800 16.990 2200.940 481.790 ;
        RECT 2197.060 16.670 2197.320 16.990 ;
        RECT 2200.740 16.670 2201.000 16.990 ;
        RECT 2197.120 2.400 2197.260 16.670 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2514.890 527.580 2515.210 527.640 ;
        RECT 2522.250 527.580 2522.570 527.640 ;
        RECT 2514.890 527.440 2522.570 527.580 ;
        RECT 2514.890 527.380 2515.210 527.440 ;
        RECT 2522.250 527.380 2522.570 527.440 ;
        RECT 2214.970 19.280 2215.290 19.340 ;
        RECT 2514.890 19.280 2515.210 19.340 ;
        RECT 2214.970 19.140 2515.210 19.280 ;
        RECT 2214.970 19.080 2215.290 19.140 ;
        RECT 2514.890 19.080 2515.210 19.140 ;
      LAYER via ;
        RECT 2514.920 527.380 2515.180 527.640 ;
        RECT 2522.280 527.380 2522.540 527.640 ;
        RECT 2215.000 19.080 2215.260 19.340 ;
        RECT 2514.920 19.080 2515.180 19.340 ;
      LAYER met2 ;
        RECT 2522.270 813.435 2522.550 813.805 ;
        RECT 2522.340 527.670 2522.480 813.435 ;
        RECT 2514.920 527.350 2515.180 527.670 ;
        RECT 2522.280 527.350 2522.540 527.670 ;
        RECT 2514.980 19.370 2515.120 527.350 ;
        RECT 2215.000 19.050 2215.260 19.370 ;
        RECT 2514.920 19.050 2515.180 19.370 ;
        RECT 2215.060 2.400 2215.200 19.050 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
      LAYER via2 ;
        RECT 2522.270 813.480 2522.550 813.760 ;
      LAYER met3 ;
        RECT 2506.000 813.770 2510.000 813.920 ;
        RECT 2522.245 813.770 2522.575 813.785 ;
        RECT 2506.000 813.470 2522.575 813.770 ;
        RECT 2506.000 813.320 2510.000 813.470 ;
        RECT 2522.245 813.455 2522.575 813.470 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 370.370 2242.880 370.690 2242.940 ;
        RECT 393.370 2242.880 393.690 2242.940 ;
        RECT 370.370 2242.740 393.690 2242.880 ;
        RECT 370.370 2242.680 370.690 2242.740 ;
        RECT 393.370 2242.680 393.690 2242.740 ;
        RECT 370.370 348.400 370.690 348.460 ;
        RECT 2228.770 348.400 2229.090 348.460 ;
        RECT 370.370 348.260 2229.090 348.400 ;
        RECT 370.370 348.200 370.690 348.260 ;
        RECT 2228.770 348.200 2229.090 348.260 ;
        RECT 2228.770 11.120 2229.090 11.180 ;
        RECT 2232.910 11.120 2233.230 11.180 ;
        RECT 2228.770 10.980 2233.230 11.120 ;
        RECT 2228.770 10.920 2229.090 10.980 ;
        RECT 2232.910 10.920 2233.230 10.980 ;
      LAYER via ;
        RECT 370.400 2242.680 370.660 2242.940 ;
        RECT 393.400 2242.680 393.660 2242.940 ;
        RECT 370.400 348.200 370.660 348.460 ;
        RECT 2228.800 348.200 2229.060 348.460 ;
        RECT 2228.800 10.920 2229.060 11.180 ;
        RECT 2232.940 10.920 2233.200 11.180 ;
      LAYER met2 ;
        RECT 393.390 2248.235 393.670 2248.605 ;
        RECT 393.460 2242.970 393.600 2248.235 ;
        RECT 370.400 2242.650 370.660 2242.970 ;
        RECT 393.400 2242.650 393.660 2242.970 ;
        RECT 370.460 348.490 370.600 2242.650 ;
        RECT 370.400 348.170 370.660 348.490 ;
        RECT 2228.800 348.170 2229.060 348.490 ;
        RECT 2228.860 11.210 2229.000 348.170 ;
        RECT 2228.800 10.890 2229.060 11.210 ;
        RECT 2232.940 10.890 2233.200 11.210 ;
        RECT 2233.000 2.400 2233.140 10.890 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 393.390 2248.280 393.670 2248.560 ;
      LAYER met3 ;
        RECT 393.365 2248.570 393.695 2248.585 ;
        RECT 410.000 2248.570 414.000 2248.720 ;
        RECT 393.365 2248.270 414.000 2248.570 ;
        RECT 393.365 2248.255 393.695 2248.270 ;
        RECT 410.000 2248.120 414.000 2248.270 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 73.680 793.430 73.740 ;
        RECT 2518.570 73.680 2518.890 73.740 ;
        RECT 793.110 73.540 2518.890 73.680 ;
        RECT 793.110 73.480 793.430 73.540 ;
        RECT 2518.570 73.480 2518.890 73.540 ;
        RECT 787.590 20.300 787.910 20.360 ;
        RECT 793.110 20.300 793.430 20.360 ;
        RECT 787.590 20.160 793.430 20.300 ;
        RECT 787.590 20.100 787.910 20.160 ;
        RECT 793.110 20.100 793.430 20.160 ;
      LAYER via ;
        RECT 793.140 73.480 793.400 73.740 ;
        RECT 2518.600 73.480 2518.860 73.740 ;
        RECT 787.620 20.100 787.880 20.360 ;
        RECT 793.140 20.100 793.400 20.360 ;
      LAYER met2 ;
        RECT 2518.590 739.995 2518.870 740.365 ;
        RECT 2518.660 73.770 2518.800 739.995 ;
        RECT 793.140 73.450 793.400 73.770 ;
        RECT 2518.600 73.450 2518.860 73.770 ;
        RECT 793.200 20.390 793.340 73.450 ;
        RECT 787.620 20.070 787.880 20.390 ;
        RECT 793.140 20.070 793.400 20.390 ;
        RECT 787.680 2.400 787.820 20.070 ;
        RECT 787.470 -4.800 788.030 2.400 ;
      LAYER via2 ;
        RECT 2518.590 740.040 2518.870 740.320 ;
      LAYER met3 ;
        RECT 2506.000 740.330 2510.000 740.480 ;
        RECT 2518.565 740.330 2518.895 740.345 ;
        RECT 2506.000 740.030 2518.895 740.330 ;
        RECT 2506.000 739.880 2510.000 740.030 ;
        RECT 2518.565 740.015 2518.895 740.030 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.290 3006.690 1247.570 3010.000 ;
        RECT 1248.530 3006.690 1248.810 3006.805 ;
        RECT 1247.290 3006.550 1248.810 3006.690 ;
        RECT 1247.290 3006.000 1247.570 3006.550 ;
        RECT 1248.530 3006.435 1248.810 3006.550 ;
        RECT 2250.870 17.835 2251.150 18.205 ;
        RECT 2250.940 2.400 2251.080 17.835 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
      LAYER via2 ;
        RECT 1248.530 3006.480 1248.810 3006.760 ;
        RECT 2250.870 17.880 2251.150 18.160 ;
      LAYER met3 ;
        RECT 1248.505 3006.770 1248.835 3006.785 ;
        RECT 1293.790 3006.770 1294.170 3006.780 ;
        RECT 1248.505 3006.470 1294.170 3006.770 ;
        RECT 1248.505 3006.455 1248.835 3006.470 ;
        RECT 1293.790 3006.460 1294.170 3006.470 ;
        RECT 1293.790 3003.370 1294.170 3003.380 ;
        RECT 2476.910 3003.370 2477.290 3003.380 ;
        RECT 1293.790 3003.070 2477.290 3003.370 ;
        RECT 1293.790 3003.060 1294.170 3003.070 ;
        RECT 2476.910 3003.060 2477.290 3003.070 ;
        RECT 2250.845 18.170 2251.175 18.185 ;
        RECT 2459.430 18.170 2459.810 18.180 ;
        RECT 2250.845 17.870 2459.810 18.170 ;
        RECT 2250.845 17.855 2251.175 17.870 ;
        RECT 2459.430 17.860 2459.810 17.870 ;
      LAYER via3 ;
        RECT 1293.820 3006.460 1294.140 3006.780 ;
        RECT 1293.820 3003.060 1294.140 3003.380 ;
        RECT 2476.940 3003.060 2477.260 3003.380 ;
        RECT 2459.460 17.860 2459.780 18.180 ;
      LAYER met4 ;
        RECT 1293.815 3006.455 1294.145 3006.785 ;
        RECT 1293.830 3003.385 1294.130 3006.455 ;
        RECT 1293.815 3003.055 1294.145 3003.385 ;
        RECT 2476.935 3003.055 2477.265 3003.385 ;
        RECT 2476.950 2993.850 2477.250 3003.055 ;
        RECT 2476.030 2993.550 2477.250 2993.850 ;
        RECT 2476.030 2946.930 2476.330 2993.550 ;
        RECT 2476.030 2946.630 2477.250 2946.930 ;
        RECT 2476.950 2939.450 2477.250 2946.630 ;
        RECT 2475.110 2939.150 2477.250 2939.450 ;
        RECT 2475.110 2891.850 2475.410 2939.150 ;
        RECT 2475.110 2891.550 2478.170 2891.850 ;
        RECT 2477.870 2851.050 2478.170 2891.550 ;
        RECT 2476.950 2850.750 2478.170 2851.050 ;
        RECT 2476.950 2745.650 2477.250 2850.750 ;
        RECT 2476.950 2745.350 2478.170 2745.650 ;
        RECT 2477.870 2698.050 2478.170 2745.350 ;
        RECT 2476.950 2697.750 2478.170 2698.050 ;
        RECT 2476.950 2262.850 2477.250 2697.750 ;
        RECT 2476.950 2262.550 2479.090 2262.850 ;
        RECT 2478.790 2215.250 2479.090 2262.550 ;
        RECT 2476.950 2214.950 2479.090 2215.250 ;
        RECT 2476.950 2120.050 2477.250 2214.950 ;
        RECT 2476.950 2119.750 2479.090 2120.050 ;
        RECT 2478.790 2077.210 2479.090 2119.750 ;
        RECT 2476.950 2076.910 2479.090 2077.210 ;
        RECT 2476.950 2069.050 2477.250 2076.910 ;
        RECT 2476.030 2068.750 2477.250 2069.050 ;
        RECT 2476.030 2021.890 2476.330 2068.750 ;
        RECT 2465.470 2020.710 2466.650 2021.890 ;
        RECT 2475.590 2020.710 2476.770 2021.890 ;
        RECT 2465.910 1974.290 2466.210 2020.710 ;
        RECT 2465.470 1973.110 2466.650 1974.290 ;
        RECT 2476.510 1973.110 2477.690 1974.290 ;
        RECT 2476.950 1810.650 2477.250 1973.110 ;
        RECT 2476.030 1810.350 2477.250 1810.650 ;
        RECT 2476.030 1773.250 2476.330 1810.350 ;
        RECT 2476.030 1772.950 2477.250 1773.250 ;
        RECT 2476.950 1735.850 2477.250 1772.950 ;
        RECT 2475.110 1735.550 2477.250 1735.850 ;
        RECT 2475.110 1715.890 2475.410 1735.550 ;
        RECT 2474.670 1714.710 2475.850 1715.890 ;
        RECT 2481.110 1714.710 2482.290 1715.890 ;
        RECT 2481.550 1671.250 2481.850 1714.710 ;
        RECT 2480.630 1670.950 2481.850 1671.250 ;
        RECT 2480.630 1667.850 2480.930 1670.950 ;
        RECT 2477.870 1667.550 2480.930 1667.850 ;
        RECT 2477.870 1637.250 2478.170 1667.550 ;
        RECT 2476.950 1636.950 2478.170 1637.250 ;
        RECT 2476.950 1501.250 2477.250 1636.950 ;
        RECT 2476.950 1500.950 2479.090 1501.250 ;
        RECT 2478.790 1453.650 2479.090 1500.950 ;
        RECT 2476.950 1453.350 2479.090 1453.650 ;
        RECT 2476.950 920.290 2477.250 1453.350 ;
        RECT 2459.030 919.110 2460.210 920.290 ;
        RECT 2476.510 919.110 2477.690 920.290 ;
        RECT 2459.470 18.185 2459.770 919.110 ;
        RECT 2459.455 17.855 2459.785 18.185 ;
      LAYER met5 ;
        RECT 2465.260 2020.500 2476.980 2022.100 ;
        RECT 2465.260 1972.900 2477.900 1974.500 ;
        RECT 2474.460 1714.500 2482.500 1716.100 ;
        RECT 2458.820 918.900 2477.900 920.500 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 508.200 2270.030 508.260 ;
        RECT 2528.230 508.200 2528.550 508.260 ;
        RECT 2269.710 508.060 2528.550 508.200 ;
        RECT 2269.710 508.000 2270.030 508.060 ;
        RECT 2528.230 508.000 2528.550 508.060 ;
        RECT 2268.330 14.180 2268.650 14.240 ;
        RECT 2269.710 14.180 2270.030 14.240 ;
        RECT 2268.330 14.040 2270.030 14.180 ;
        RECT 2268.330 13.980 2268.650 14.040 ;
        RECT 2269.710 13.980 2270.030 14.040 ;
      LAYER via ;
        RECT 2269.740 508.000 2270.000 508.260 ;
        RECT 2528.260 508.000 2528.520 508.260 ;
        RECT 2268.360 13.980 2268.620 14.240 ;
        RECT 2269.740 13.980 2270.000 14.240 ;
      LAYER met2 ;
        RECT 2528.250 904.555 2528.530 904.925 ;
        RECT 2528.320 508.290 2528.460 904.555 ;
        RECT 2269.740 507.970 2270.000 508.290 ;
        RECT 2528.260 507.970 2528.520 508.290 ;
        RECT 2269.800 14.270 2269.940 507.970 ;
        RECT 2268.360 13.950 2268.620 14.270 ;
        RECT 2269.740 13.950 2270.000 14.270 ;
        RECT 2268.420 2.400 2268.560 13.950 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
      LAYER via2 ;
        RECT 2528.250 904.600 2528.530 904.880 ;
      LAYER met3 ;
        RECT 2506.000 904.890 2510.000 905.040 ;
        RECT 2528.225 904.890 2528.555 904.905 ;
        RECT 2506.000 904.590 2528.555 904.890 ;
        RECT 2506.000 904.440 2510.000 904.590 ;
        RECT 2528.225 904.575 2528.555 904.590 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 868.550 99.860 868.870 99.920 ;
        RECT 2283.970 99.860 2284.290 99.920 ;
        RECT 868.550 99.720 2284.290 99.860 ;
        RECT 868.550 99.660 868.870 99.720 ;
        RECT 2283.970 99.660 2284.290 99.720 ;
      LAYER via ;
        RECT 868.580 99.660 868.840 99.920 ;
        RECT 2284.000 99.660 2284.260 99.920 ;
      LAYER met2 ;
        RECT 869.170 510.410 869.450 514.000 ;
        RECT 868.640 510.270 869.450 510.410 ;
        RECT 868.640 99.950 868.780 510.270 ;
        RECT 869.170 510.000 869.450 510.270 ;
        RECT 868.580 99.630 868.840 99.950 ;
        RECT 2284.000 99.630 2284.260 99.950 ;
        RECT 2284.060 16.730 2284.200 99.630 ;
        RECT 2284.060 16.590 2286.500 16.730 ;
        RECT 2286.360 2.400 2286.500 16.590 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 288.950 1676.780 289.270 1676.840 ;
        RECT 393.370 1676.780 393.690 1676.840 ;
        RECT 288.950 1676.640 393.690 1676.780 ;
        RECT 288.950 1676.580 289.270 1676.640 ;
        RECT 393.370 1676.580 393.690 1676.640 ;
        RECT 288.950 72.660 289.270 72.720 ;
        RECT 2297.770 72.660 2298.090 72.720 ;
        RECT 288.950 72.520 2298.090 72.660 ;
        RECT 288.950 72.460 289.270 72.520 ;
        RECT 2297.770 72.460 2298.090 72.520 ;
        RECT 2297.770 16.900 2298.090 16.960 ;
        RECT 2304.210 16.900 2304.530 16.960 ;
        RECT 2297.770 16.760 2304.530 16.900 ;
        RECT 2297.770 16.700 2298.090 16.760 ;
        RECT 2304.210 16.700 2304.530 16.760 ;
      LAYER via ;
        RECT 288.980 1676.580 289.240 1676.840 ;
        RECT 393.400 1676.580 393.660 1676.840 ;
        RECT 288.980 72.460 289.240 72.720 ;
        RECT 2297.800 72.460 2298.060 72.720 ;
        RECT 2297.800 16.700 2298.060 16.960 ;
        RECT 2304.240 16.700 2304.500 16.960 ;
      LAYER met2 ;
        RECT 393.390 1682.475 393.670 1682.845 ;
        RECT 393.460 1676.870 393.600 1682.475 ;
        RECT 288.980 1676.550 289.240 1676.870 ;
        RECT 393.400 1676.550 393.660 1676.870 ;
        RECT 289.040 72.750 289.180 1676.550 ;
        RECT 288.980 72.430 289.240 72.750 ;
        RECT 2297.800 72.430 2298.060 72.750 ;
        RECT 2297.860 16.990 2298.000 72.430 ;
        RECT 2297.800 16.670 2298.060 16.990 ;
        RECT 2304.240 16.670 2304.500 16.990 ;
        RECT 2304.300 2.400 2304.440 16.670 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 393.390 1682.520 393.670 1682.800 ;
      LAYER met3 ;
        RECT 393.365 1682.810 393.695 1682.825 ;
        RECT 410.000 1682.810 414.000 1682.960 ;
        RECT 393.365 1682.510 414.000 1682.810 ;
        RECT 393.365 1682.495 393.695 1682.510 ;
        RECT 410.000 1682.360 414.000 1682.510 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2075.290 3006.690 2075.570 3010.000 ;
        RECT 2076.990 3006.690 2077.270 3006.805 ;
        RECT 2075.290 3006.550 2077.270 3006.690 ;
        RECT 2075.290 3006.000 2075.570 3006.550 ;
        RECT 2076.990 3006.435 2077.270 3006.550 ;
        RECT 2322.170 19.195 2322.450 19.565 ;
        RECT 2322.240 2.400 2322.380 19.195 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 2076.990 3006.480 2077.270 3006.760 ;
        RECT 2322.170 19.240 2322.450 19.520 ;
      LAYER met3 ;
        RECT 2076.965 3006.770 2077.295 3006.785 ;
        RECT 2076.965 3006.470 2079.810 3006.770 ;
        RECT 2076.965 3006.455 2077.295 3006.470 ;
        RECT 2079.510 3004.050 2079.810 3006.470 ;
        RECT 2491.630 3004.050 2492.010 3004.060 ;
        RECT 2079.510 3003.750 2492.010 3004.050 ;
        RECT 2491.630 3003.740 2492.010 3003.750 ;
        RECT 2322.145 19.530 2322.475 19.545 ;
        RECT 2451.150 19.530 2451.530 19.540 ;
        RECT 2322.145 19.230 2451.530 19.530 ;
        RECT 2322.145 19.215 2322.475 19.230 ;
        RECT 2451.150 19.220 2451.530 19.230 ;
      LAYER via3 ;
        RECT 2491.660 3003.740 2491.980 3004.060 ;
        RECT 2451.180 19.220 2451.500 19.540 ;
      LAYER met4 ;
        RECT 2491.655 3003.735 2491.985 3004.065 ;
        RECT 2491.670 2291.410 2491.970 3003.735 ;
        RECT 2491.670 2291.110 2496.570 2291.410 ;
        RECT 2496.270 2266.250 2496.570 2291.110 ;
        RECT 2491.670 2265.950 2496.570 2266.250 ;
        RECT 2491.670 1212.690 2491.970 2265.950 ;
        RECT 2491.230 1211.510 2492.410 1212.690 ;
        RECT 2450.750 1204.710 2451.930 1205.890 ;
        RECT 2451.190 19.545 2451.490 1204.710 ;
        RECT 2451.175 19.215 2451.505 19.545 ;
      LAYER met5 ;
        RECT 2491.020 1211.300 2493.540 1212.900 ;
        RECT 2491.940 1206.100 2493.540 1211.300 ;
        RECT 2450.540 1204.500 2493.540 1206.100 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2277.530 501.400 2277.850 501.460 ;
        RECT 2283.510 501.400 2283.830 501.460 ;
        RECT 2277.530 501.260 2283.830 501.400 ;
        RECT 2277.530 501.200 2277.850 501.260 ;
        RECT 2283.510 501.200 2283.830 501.260 ;
        RECT 2283.510 24.720 2283.830 24.780 ;
        RECT 2339.630 24.720 2339.950 24.780 ;
        RECT 2283.510 24.580 2339.950 24.720 ;
        RECT 2283.510 24.520 2283.830 24.580 ;
        RECT 2339.630 24.520 2339.950 24.580 ;
      LAYER via ;
        RECT 2277.560 501.200 2277.820 501.460 ;
        RECT 2283.540 501.200 2283.800 501.460 ;
        RECT 2283.540 24.520 2283.800 24.780 ;
        RECT 2339.660 24.520 2339.920 24.780 ;
      LAYER met2 ;
        RECT 2277.690 510.340 2277.970 514.000 ;
        RECT 2277.620 510.000 2277.970 510.340 ;
        RECT 2277.620 501.490 2277.760 510.000 ;
        RECT 2277.560 501.170 2277.820 501.490 ;
        RECT 2283.540 501.170 2283.800 501.490 ;
        RECT 2283.600 24.810 2283.740 501.170 ;
        RECT 2283.540 24.490 2283.800 24.810 ;
        RECT 2339.660 24.490 2339.920 24.810 ;
        RECT 2339.720 2.400 2339.860 24.490 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1790.850 3023.520 1791.170 3023.580 ;
        RECT 2519.030 3023.520 2519.350 3023.580 ;
        RECT 1790.850 3023.380 2519.350 3023.520 ;
        RECT 1790.850 3023.320 1791.170 3023.380 ;
        RECT 2519.030 3023.320 2519.350 3023.380 ;
      LAYER via ;
        RECT 1790.880 3023.320 1791.140 3023.580 ;
        RECT 2519.060 3023.320 2519.320 3023.580 ;
      LAYER met2 ;
        RECT 1790.880 3023.290 1791.140 3023.610 ;
        RECT 2519.060 3023.290 2519.320 3023.610 ;
        RECT 1790.940 3010.000 1791.080 3023.290 ;
        RECT 1790.940 3009.340 1791.290 3010.000 ;
        RECT 1791.010 3006.000 1791.290 3009.340 ;
        RECT 2519.120 906.285 2519.260 3023.290 ;
        RECT 2519.050 905.915 2519.330 906.285 ;
        RECT 2357.590 33.475 2357.870 33.845 ;
        RECT 2357.660 2.400 2357.800 33.475 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
      LAYER via2 ;
        RECT 2519.050 905.960 2519.330 906.240 ;
        RECT 2357.590 33.520 2357.870 33.800 ;
      LAYER met3 ;
        RECT 2516.470 906.250 2516.850 906.260 ;
        RECT 2519.025 906.250 2519.355 906.265 ;
        RECT 2516.470 905.950 2519.355 906.250 ;
        RECT 2516.470 905.940 2516.850 905.950 ;
        RECT 2519.025 905.935 2519.355 905.950 ;
        RECT 2357.565 33.810 2357.895 33.825 ;
        RECT 2477.830 33.810 2478.210 33.820 ;
        RECT 2357.565 33.510 2478.210 33.810 ;
        RECT 2357.565 33.495 2357.895 33.510 ;
        RECT 2477.830 33.500 2478.210 33.510 ;
      LAYER via3 ;
        RECT 2516.500 905.940 2516.820 906.260 ;
        RECT 2477.860 33.500 2478.180 33.820 ;
      LAYER met4 ;
        RECT 2516.070 905.510 2517.250 906.690 ;
        RECT 2477.430 902.110 2478.610 903.290 ;
        RECT 2477.870 33.825 2478.170 902.110 ;
        RECT 2477.855 33.495 2478.185 33.825 ;
      LAYER met5 ;
        RECT 2477.220 905.300 2517.460 906.900 ;
        RECT 2477.220 901.900 2478.820 905.300 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2228.385 33.405 2228.555 47.855 ;
      LAYER mcon ;
        RECT 2228.385 47.685 2228.555 47.855 ;
      LAYER met1 ;
        RECT 2227.850 289.920 2228.170 289.980 ;
        RECT 2228.310 289.920 2228.630 289.980 ;
        RECT 2227.850 289.780 2228.630 289.920 ;
        RECT 2227.850 289.720 2228.170 289.780 ;
        RECT 2228.310 289.720 2228.630 289.780 ;
        RECT 2227.850 193.360 2228.170 193.420 ;
        RECT 2228.310 193.360 2228.630 193.420 ;
        RECT 2227.850 193.220 2228.630 193.360 ;
        RECT 2227.850 193.160 2228.170 193.220 ;
        RECT 2228.310 193.160 2228.630 193.220 ;
        RECT 2227.850 96.800 2228.170 96.860 ;
        RECT 2228.310 96.800 2228.630 96.860 ;
        RECT 2227.850 96.660 2228.630 96.800 ;
        RECT 2227.850 96.600 2228.170 96.660 ;
        RECT 2228.310 96.600 2228.630 96.660 ;
        RECT 2228.310 47.840 2228.630 47.900 ;
        RECT 2228.115 47.700 2228.630 47.840 ;
        RECT 2228.310 47.640 2228.630 47.700 ;
        RECT 2228.325 33.560 2228.615 33.605 ;
        RECT 2375.510 33.560 2375.830 33.620 ;
        RECT 2228.325 33.420 2375.830 33.560 ;
        RECT 2228.325 33.375 2228.615 33.420 ;
        RECT 2375.510 33.360 2375.830 33.420 ;
      LAYER via ;
        RECT 2227.880 289.720 2228.140 289.980 ;
        RECT 2228.340 289.720 2228.600 289.980 ;
        RECT 2227.880 193.160 2228.140 193.420 ;
        RECT 2228.340 193.160 2228.600 193.420 ;
        RECT 2227.880 96.600 2228.140 96.860 ;
        RECT 2228.340 96.600 2228.600 96.860 ;
        RECT 2228.340 47.640 2228.600 47.900 ;
        RECT 2375.540 33.360 2375.800 33.620 ;
      LAYER met2 ;
        RECT 2228.010 510.410 2228.290 514.000 ;
        RECT 2227.480 510.270 2228.290 510.410 ;
        RECT 2227.480 483.325 2227.620 510.270 ;
        RECT 2228.010 510.000 2228.290 510.270 ;
        RECT 2227.410 482.955 2227.690 483.325 ;
        RECT 2228.330 482.955 2228.610 483.325 ;
        RECT 2228.400 337.690 2228.540 482.955 ;
        RECT 2227.940 337.550 2228.540 337.690 ;
        RECT 2227.940 290.010 2228.080 337.550 ;
        RECT 2227.880 289.690 2228.140 290.010 ;
        RECT 2228.340 289.690 2228.600 290.010 ;
        RECT 2228.400 241.130 2228.540 289.690 ;
        RECT 2227.940 240.990 2228.540 241.130 ;
        RECT 2227.940 193.450 2228.080 240.990 ;
        RECT 2227.880 193.130 2228.140 193.450 ;
        RECT 2228.340 193.130 2228.600 193.450 ;
        RECT 2228.400 144.570 2228.540 193.130 ;
        RECT 2227.940 144.430 2228.540 144.570 ;
        RECT 2227.940 96.890 2228.080 144.430 ;
        RECT 2227.880 96.570 2228.140 96.890 ;
        RECT 2228.340 96.570 2228.600 96.890 ;
        RECT 2228.400 47.930 2228.540 96.570 ;
        RECT 2228.340 47.610 2228.600 47.930 ;
        RECT 2375.540 33.330 2375.800 33.650 ;
        RECT 2375.600 2.400 2375.740 33.330 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
      LAYER via2 ;
        RECT 2227.410 483.000 2227.690 483.280 ;
        RECT 2228.330 483.000 2228.610 483.280 ;
      LAYER met3 ;
        RECT 2227.385 483.290 2227.715 483.305 ;
        RECT 2228.305 483.290 2228.635 483.305 ;
        RECT 2227.385 482.990 2228.635 483.290 ;
        RECT 2227.385 482.975 2227.715 482.990 ;
        RECT 2228.305 482.975 2228.635 482.990 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2393.910 500.380 2394.230 500.440 ;
        RECT 2528.690 500.380 2529.010 500.440 ;
        RECT 2393.910 500.240 2529.010 500.380 ;
        RECT 2393.910 500.180 2394.230 500.240 ;
        RECT 2528.690 500.180 2529.010 500.240 ;
      LAYER via ;
        RECT 2393.940 500.180 2394.200 500.440 ;
        RECT 2528.720 500.180 2528.980 500.440 ;
      LAYER met2 ;
        RECT 2528.710 648.875 2528.990 649.245 ;
        RECT 2528.780 500.470 2528.920 648.875 ;
        RECT 2393.940 500.150 2394.200 500.470 ;
        RECT 2528.720 500.150 2528.980 500.470 ;
        RECT 2394.000 17.410 2394.140 500.150 ;
        RECT 2393.540 17.270 2394.140 17.410 ;
        RECT 2393.540 2.400 2393.680 17.270 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 2528.710 648.920 2528.990 649.200 ;
      LAYER met3 ;
        RECT 2506.000 649.210 2510.000 649.360 ;
        RECT 2528.685 649.210 2529.015 649.225 ;
        RECT 2506.000 648.910 2529.015 649.210 ;
        RECT 2506.000 648.760 2510.000 648.910 ;
        RECT 2528.685 648.895 2529.015 648.910 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2408.190 389.115 2408.470 389.485 ;
        RECT 2408.260 16.730 2408.400 389.115 ;
        RECT 2408.260 16.590 2411.620 16.730 ;
        RECT 2411.480 2.400 2411.620 16.590 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 2408.190 389.160 2408.470 389.440 ;
      LAYER met3 ;
        RECT 410.000 2120.280 414.000 2120.880 ;
        RECT 370.110 2118.690 370.490 2118.700 ;
        RECT 410.630 2118.690 410.930 2120.280 ;
        RECT 370.110 2118.390 410.930 2118.690 ;
        RECT 370.110 2118.380 370.490 2118.390 ;
        RECT 370.110 389.450 370.490 389.460 ;
        RECT 2408.165 389.450 2408.495 389.465 ;
        RECT 370.110 389.150 2408.495 389.450 ;
        RECT 370.110 389.140 370.490 389.150 ;
        RECT 2408.165 389.135 2408.495 389.150 ;
      LAYER via3 ;
        RECT 370.140 2118.380 370.460 2118.700 ;
        RECT 370.140 389.140 370.460 389.460 ;
      LAYER met4 ;
        RECT 370.135 2118.375 370.465 2118.705 ;
        RECT 370.150 389.465 370.450 2118.375 ;
        RECT 370.135 389.135 370.465 389.465 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1782.645 483.225 1782.815 501.415 ;
        RECT 1783.565 351.305 1783.735 385.815 ;
        RECT 1783.105 241.485 1783.275 289.595 ;
      LAYER mcon ;
        RECT 1782.645 501.245 1782.815 501.415 ;
        RECT 1783.565 385.645 1783.735 385.815 ;
        RECT 1783.105 289.425 1783.275 289.595 ;
      LAYER met1 ;
        RECT 1782.585 501.400 1782.875 501.445 ;
        RECT 1881.930 501.400 1882.250 501.460 ;
        RECT 1782.585 501.260 1882.250 501.400 ;
        RECT 1782.585 501.215 1782.875 501.260 ;
        RECT 1881.930 501.200 1882.250 501.260 ;
        RECT 1782.570 483.380 1782.890 483.440 ;
        RECT 1782.375 483.240 1782.890 483.380 ;
        RECT 1782.570 483.180 1782.890 483.240 ;
        RECT 1782.570 448.500 1782.890 448.760 ;
        RECT 1782.660 448.020 1782.800 448.500 ;
        RECT 1783.030 448.020 1783.350 448.080 ;
        RECT 1782.660 447.880 1783.350 448.020 ;
        RECT 1783.030 447.820 1783.350 447.880 ;
        RECT 1783.030 400.220 1783.350 400.480 ;
        RECT 1783.120 399.740 1783.260 400.220 ;
        RECT 1783.490 399.740 1783.810 399.800 ;
        RECT 1783.120 399.600 1783.810 399.740 ;
        RECT 1783.490 399.540 1783.810 399.600 ;
        RECT 1783.490 385.800 1783.810 385.860 ;
        RECT 1783.295 385.660 1783.810 385.800 ;
        RECT 1783.490 385.600 1783.810 385.660 ;
        RECT 1783.505 351.460 1783.795 351.505 ;
        RECT 1783.950 351.460 1784.270 351.520 ;
        RECT 1783.505 351.320 1784.270 351.460 ;
        RECT 1783.505 351.275 1783.795 351.320 ;
        RECT 1783.950 351.260 1784.270 351.320 ;
        RECT 1783.030 289.580 1783.350 289.640 ;
        RECT 1782.835 289.440 1783.350 289.580 ;
        RECT 1783.030 289.380 1783.350 289.440 ;
        RECT 1783.045 241.640 1783.335 241.685 ;
        RECT 1783.490 241.640 1783.810 241.700 ;
        RECT 1783.045 241.500 1783.810 241.640 ;
        RECT 1783.045 241.455 1783.335 241.500 ;
        RECT 1783.490 241.440 1783.810 241.500 ;
        RECT 806.910 190.300 807.230 190.360 ;
        RECT 1784.410 190.300 1784.730 190.360 ;
        RECT 806.910 190.160 1784.730 190.300 ;
        RECT 806.910 190.100 807.230 190.160 ;
        RECT 1784.410 190.100 1784.730 190.160 ;
        RECT 805.530 14.180 805.850 14.240 ;
        RECT 806.910 14.180 807.230 14.240 ;
        RECT 805.530 14.040 807.230 14.180 ;
        RECT 805.530 13.980 805.850 14.040 ;
        RECT 806.910 13.980 807.230 14.040 ;
      LAYER via ;
        RECT 1881.960 501.200 1882.220 501.460 ;
        RECT 1782.600 483.180 1782.860 483.440 ;
        RECT 1782.600 448.500 1782.860 448.760 ;
        RECT 1783.060 447.820 1783.320 448.080 ;
        RECT 1783.060 400.220 1783.320 400.480 ;
        RECT 1783.520 399.540 1783.780 399.800 ;
        RECT 1783.520 385.600 1783.780 385.860 ;
        RECT 1783.980 351.260 1784.240 351.520 ;
        RECT 1783.060 289.380 1783.320 289.640 ;
        RECT 1783.520 241.440 1783.780 241.700 ;
        RECT 806.940 190.100 807.200 190.360 ;
        RECT 1784.440 190.100 1784.700 190.360 ;
        RECT 805.560 13.980 805.820 14.240 ;
        RECT 806.940 13.980 807.200 14.240 ;
      LAYER met2 ;
        RECT 1882.090 510.340 1882.370 514.000 ;
        RECT 1882.020 510.000 1882.370 510.340 ;
        RECT 1882.020 501.490 1882.160 510.000 ;
        RECT 1881.960 501.170 1882.220 501.490 ;
        RECT 1782.600 483.150 1782.860 483.470 ;
        RECT 1782.660 448.790 1782.800 483.150 ;
        RECT 1782.600 448.470 1782.860 448.790 ;
        RECT 1783.060 447.790 1783.320 448.110 ;
        RECT 1783.120 400.510 1783.260 447.790 ;
        RECT 1783.060 400.190 1783.320 400.510 ;
        RECT 1783.520 399.510 1783.780 399.830 ;
        RECT 1783.580 385.890 1783.720 399.510 ;
        RECT 1783.520 385.570 1783.780 385.890 ;
        RECT 1783.980 351.230 1784.240 351.550 ;
        RECT 1784.040 303.690 1784.180 351.230 ;
        RECT 1783.120 303.550 1784.180 303.690 ;
        RECT 1783.120 289.670 1783.260 303.550 ;
        RECT 1783.060 289.350 1783.320 289.670 ;
        RECT 1783.520 241.410 1783.780 241.730 ;
        RECT 1783.580 207.130 1783.720 241.410 ;
        RECT 1783.580 206.990 1784.640 207.130 ;
        RECT 1784.500 190.390 1784.640 206.990 ;
        RECT 806.940 190.070 807.200 190.390 ;
        RECT 1784.440 190.070 1784.700 190.390 ;
        RECT 807.000 14.270 807.140 190.070 ;
        RECT 805.560 13.950 805.820 14.270 ;
        RECT 806.940 13.950 807.200 14.270 ;
        RECT 805.620 2.400 805.760 13.950 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.150 3010.600 45.470 3010.660 ;
        RECT 604.970 3010.600 605.290 3010.660 ;
        RECT 45.150 3010.460 605.290 3010.600 ;
        RECT 45.150 3010.400 45.470 3010.460 ;
        RECT 604.970 3010.400 605.290 3010.460 ;
        RECT 2.830 20.300 3.150 20.360 ;
        RECT 45.150 20.300 45.470 20.360 ;
        RECT 2.830 20.160 45.470 20.300 ;
        RECT 2.830 20.100 3.150 20.160 ;
        RECT 45.150 20.100 45.470 20.160 ;
      LAYER via ;
        RECT 45.180 3010.400 45.440 3010.660 ;
        RECT 605.000 3010.400 605.260 3010.660 ;
        RECT 2.860 20.100 3.120 20.360 ;
        RECT 45.180 20.100 45.440 20.360 ;
      LAYER met2 ;
        RECT 45.180 3010.370 45.440 3010.690 ;
        RECT 605.000 3010.370 605.260 3010.690 ;
        RECT 45.240 20.390 45.380 3010.370 ;
        RECT 605.060 3010.000 605.200 3010.370 ;
        RECT 605.060 3009.340 605.410 3010.000 ;
        RECT 605.130 3006.000 605.410 3009.340 ;
        RECT 2.860 20.070 3.120 20.390 ;
        RECT 45.180 20.070 45.440 20.390 ;
        RECT 2.920 2.400 3.060 20.070 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 30.965 2996.165 31.135 2998.035 ;
        RECT 48.445 2997.185 48.615 2998.035 ;
        RECT 96.285 2997.185 96.455 2998.375 ;
        RECT 110.085 2998.205 110.715 2998.375 ;
        RECT 158.845 2997.525 159.015 2998.375 ;
        RECT 193.345 2998.205 193.515 2999.055 ;
        RECT 241.185 2997.865 241.355 2999.055 ;
        RECT 255.445 2997.525 255.615 2998.375 ;
      LAYER mcon ;
        RECT 193.345 2998.885 193.515 2999.055 ;
        RECT 96.285 2998.205 96.455 2998.375 ;
        RECT 110.545 2998.205 110.715 2998.375 ;
        RECT 158.845 2998.205 159.015 2998.375 ;
        RECT 241.185 2998.885 241.355 2999.055 ;
        RECT 30.965 2997.865 31.135 2998.035 ;
        RECT 48.445 2997.865 48.615 2998.035 ;
        RECT 255.445 2998.205 255.615 2998.375 ;
      LAYER met1 ;
        RECT 417.290 3005.500 417.610 3005.560 ;
        RECT 418.210 3005.500 418.530 3005.560 ;
        RECT 417.290 3005.360 418.530 3005.500 ;
        RECT 417.290 3005.300 417.610 3005.360 ;
        RECT 418.210 3005.300 418.530 3005.360 ;
        RECT 417.290 3000.060 417.610 3000.120 ;
        RECT 375.980 2999.920 417.610 3000.060 ;
        RECT 193.285 2999.040 193.575 2999.085 ;
        RECT 241.125 2999.040 241.415 2999.085 ;
        RECT 193.285 2998.900 241.415 2999.040 ;
        RECT 193.285 2998.855 193.575 2998.900 ;
        RECT 241.125 2998.855 241.415 2998.900 ;
        RECT 302.840 2998.560 314.020 2998.700 ;
        RECT 96.225 2998.360 96.515 2998.405 ;
        RECT 110.025 2998.360 110.315 2998.405 ;
        RECT 96.225 2998.220 110.315 2998.360 ;
        RECT 96.225 2998.175 96.515 2998.220 ;
        RECT 110.025 2998.175 110.315 2998.220 ;
        RECT 110.485 2998.360 110.775 2998.405 ;
        RECT 158.785 2998.360 159.075 2998.405 ;
        RECT 193.285 2998.360 193.575 2998.405 ;
        RECT 110.485 2998.220 116.680 2998.360 ;
        RECT 110.485 2998.175 110.775 2998.220 ;
        RECT 30.905 2998.020 31.195 2998.065 ;
        RECT 48.385 2998.020 48.675 2998.065 ;
        RECT 30.905 2997.880 48.675 2998.020 ;
        RECT 116.540 2998.020 116.680 2998.220 ;
        RECT 158.785 2998.220 193.575 2998.360 ;
        RECT 158.785 2998.175 159.075 2998.220 ;
        RECT 193.285 2998.175 193.575 2998.220 ;
        RECT 255.385 2998.360 255.675 2998.405 ;
        RECT 302.840 2998.360 302.980 2998.560 ;
        RECT 255.385 2998.220 302.980 2998.360 ;
        RECT 255.385 2998.175 255.675 2998.220 ;
        RECT 241.125 2998.020 241.415 2998.065 ;
        RECT 313.880 2998.020 314.020 2998.560 ;
        RECT 375.980 2998.020 376.120 2999.920 ;
        RECT 417.290 2999.860 417.610 2999.920 ;
        RECT 116.540 2997.880 158.540 2998.020 ;
        RECT 30.905 2997.835 31.195 2997.880 ;
        RECT 48.385 2997.835 48.675 2997.880 ;
        RECT 158.400 2997.680 158.540 2997.880 ;
        RECT 241.125 2997.880 255.140 2998.020 ;
        RECT 313.880 2997.880 376.120 2998.020 ;
        RECT 241.125 2997.835 241.415 2997.880 ;
        RECT 158.785 2997.680 159.075 2997.725 ;
        RECT 158.400 2997.540 159.075 2997.680 ;
        RECT 255.000 2997.680 255.140 2997.880 ;
        RECT 255.385 2997.680 255.675 2997.725 ;
        RECT 255.000 2997.540 255.675 2997.680 ;
        RECT 158.785 2997.495 159.075 2997.540 ;
        RECT 255.385 2997.495 255.675 2997.540 ;
        RECT 48.385 2997.340 48.675 2997.385 ;
        RECT 96.225 2997.340 96.515 2997.385 ;
        RECT 48.385 2997.200 96.515 2997.340 ;
        RECT 48.385 2997.155 48.675 2997.200 ;
        RECT 96.225 2997.155 96.515 2997.200 ;
        RECT 13.410 2996.320 13.730 2996.380 ;
        RECT 30.905 2996.320 31.195 2996.365 ;
        RECT 13.410 2996.180 31.195 2996.320 ;
        RECT 13.410 2996.120 13.730 2996.180 ;
        RECT 30.905 2996.135 31.195 2996.180 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 417.320 3005.300 417.580 3005.560 ;
        RECT 418.240 3005.300 418.500 3005.560 ;
        RECT 417.320 2999.860 417.580 3000.120 ;
        RECT 13.440 2996.120 13.700 2996.380 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 419.290 3006.690 419.570 3010.000 ;
        RECT 418.300 3006.550 419.570 3006.690 ;
        RECT 418.300 3005.590 418.440 3006.550 ;
        RECT 419.290 3006.000 419.570 3006.550 ;
        RECT 417.320 3005.270 417.580 3005.590 ;
        RECT 418.240 3005.270 418.500 3005.590 ;
        RECT 417.380 3000.150 417.520 3005.270 ;
        RECT 417.320 2999.830 417.580 3000.150 ;
        RECT 13.440 2996.090 13.700 2996.410 ;
        RECT 13.500 17.670 13.640 2996.090 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.240 14.650 17.300 ;
        RECT 65.390 17.240 65.710 17.300 ;
        RECT 14.330 17.100 65.710 17.240 ;
        RECT 14.330 17.040 14.650 17.100 ;
        RECT 65.390 17.040 65.710 17.100 ;
      LAYER via ;
        RECT 14.360 17.040 14.620 17.300 ;
        RECT 65.420 17.040 65.680 17.300 ;
      LAYER met2 ;
        RECT 1530.050 3006.690 1530.330 3006.805 ;
        RECT 1531.570 3006.690 1531.850 3010.000 ;
        RECT 1530.050 3006.550 1531.850 3006.690 ;
        RECT 1530.050 3006.435 1530.330 3006.550 ;
        RECT 1531.570 3006.000 1531.850 3006.550 ;
        RECT 65.410 3002.355 65.690 3002.725 ;
        RECT 65.480 17.330 65.620 3002.355 ;
        RECT 14.360 17.010 14.620 17.330 ;
        RECT 65.420 17.010 65.680 17.330 ;
        RECT 14.420 2.400 14.560 17.010 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 1530.050 3006.480 1530.330 3006.760 ;
        RECT 65.410 3002.400 65.690 3002.680 ;
      LAYER met3 ;
        RECT 1507.230 3006.770 1507.610 3006.780 ;
        RECT 1530.025 3006.770 1530.355 3006.785 ;
        RECT 1507.230 3006.470 1530.355 3006.770 ;
        RECT 1507.230 3006.460 1507.610 3006.470 ;
        RECT 1530.025 3006.455 1530.355 3006.470 ;
        RECT 65.385 3002.690 65.715 3002.705 ;
        RECT 1507.230 3002.690 1507.610 3002.700 ;
        RECT 65.385 3002.390 1507.610 3002.690 ;
        RECT 65.385 3002.375 65.715 3002.390 ;
        RECT 1507.230 3002.380 1507.610 3002.390 ;
      LAYER via3 ;
        RECT 1507.260 3006.460 1507.580 3006.780 ;
        RECT 1507.260 3002.380 1507.580 3002.700 ;
      LAYER met4 ;
        RECT 1507.255 3006.455 1507.585 3006.785 ;
        RECT 1507.270 3002.705 1507.570 3006.455 ;
        RECT 1507.255 3002.375 1507.585 3002.705 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 529.145 3001.605 529.315 3006.535 ;
      LAYER mcon ;
        RECT 529.145 3006.365 529.315 3006.535 ;
      LAYER met1 ;
        RECT 529.070 3006.520 529.390 3006.580 ;
        RECT 528.875 3006.380 529.390 3006.520 ;
        RECT 529.070 3006.320 529.390 3006.380 ;
        RECT 79.190 3001.760 79.510 3001.820 ;
        RECT 529.085 3001.760 529.375 3001.805 ;
        RECT 79.190 3001.620 529.375 3001.760 ;
        RECT 79.190 3001.560 79.510 3001.620 ;
        RECT 529.085 3001.575 529.375 3001.620 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 79.190 17.920 79.510 17.980 ;
        RECT 38.250 17.780 79.510 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 79.190 17.720 79.510 17.780 ;
      LAYER via ;
        RECT 529.100 3006.320 529.360 3006.580 ;
        RECT 79.220 3001.560 79.480 3001.820 ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 79.220 17.720 79.480 17.980 ;
      LAYER met2 ;
        RECT 530.610 3006.690 530.890 3010.000 ;
        RECT 529.160 3006.610 530.890 3006.690 ;
        RECT 529.100 3006.550 530.890 3006.610 ;
        RECT 529.100 3006.290 529.360 3006.550 ;
        RECT 530.610 3006.000 530.890 3006.550 ;
        RECT 79.220 3001.530 79.480 3001.850 ;
        RECT 79.280 18.010 79.420 3001.530 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 79.220 17.690 79.480 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.470 3011.620 524.790 3011.680 ;
        RECT 2321.690 3011.620 2322.010 3011.680 ;
        RECT 524.470 3011.480 2322.010 3011.620 ;
        RECT 524.470 3011.420 524.790 3011.480 ;
        RECT 2321.690 3011.420 2322.010 3011.480 ;
      LAYER via ;
        RECT 524.500 3011.420 524.760 3011.680 ;
        RECT 2321.720 3011.420 2321.980 3011.680 ;
      LAYER met2 ;
        RECT 524.500 3011.390 524.760 3011.710 ;
        RECT 2321.720 3011.390 2321.980 3011.710 ;
        RECT 524.560 3009.525 524.700 3011.390 ;
        RECT 2321.780 3010.000 2321.920 3011.390 ;
        RECT 241.130 3009.155 241.410 3009.525 ;
        RECT 524.490 3009.155 524.770 3009.525 ;
        RECT 2321.780 3009.340 2322.130 3010.000 ;
        RECT 241.200 17.410 241.340 3009.155 ;
        RECT 2321.850 3006.000 2322.130 3009.340 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 241.130 3009.200 241.410 3009.480 ;
        RECT 524.490 3009.200 524.770 3009.480 ;
      LAYER met3 ;
        RECT 241.105 3009.490 241.435 3009.505 ;
        RECT 524.465 3009.490 524.795 3009.505 ;
        RECT 241.105 3009.190 524.795 3009.490 ;
        RECT 241.105 3009.175 241.435 3009.190 ;
        RECT 524.465 3009.175 524.795 3009.190 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 17.580 258.450 17.640 ;
        RECT 261.810 17.580 262.130 17.640 ;
        RECT 258.130 17.440 262.130 17.580 ;
        RECT 258.130 17.380 258.450 17.440 ;
        RECT 261.810 17.380 262.130 17.440 ;
      LAYER via ;
        RECT 258.160 17.380 258.420 17.640 ;
        RECT 261.840 17.380 262.100 17.640 ;
      LAYER met2 ;
        RECT 261.830 3008.475 262.110 3008.845 ;
        RECT 1838.250 3008.730 1838.530 3008.845 ;
        RECT 1839.770 3008.730 1840.050 3010.000 ;
        RECT 1838.250 3008.590 1840.050 3008.730 ;
        RECT 1838.250 3008.475 1838.530 3008.590 ;
        RECT 261.900 17.670 262.040 3008.475 ;
        RECT 1839.770 3006.000 1840.050 3008.590 ;
        RECT 258.160 17.350 258.420 17.670 ;
        RECT 261.840 17.350 262.100 17.670 ;
        RECT 258.220 2.400 258.360 17.350 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 261.830 3008.520 262.110 3008.800 ;
        RECT 1838.250 3008.520 1838.530 3008.800 ;
      LAYER met3 ;
        RECT 261.805 3008.810 262.135 3008.825 ;
        RECT 1838.225 3008.810 1838.555 3008.825 ;
        RECT 261.805 3008.510 1838.555 3008.810 ;
        RECT 261.805 3008.495 262.135 3008.510 ;
        RECT 1838.225 3008.495 1838.555 3008.510 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2495.590 503.355 2495.870 503.725 ;
        RECT 2495.660 338.485 2495.800 503.355 ;
        RECT 2495.590 338.115 2495.870 338.485 ;
        RECT 2496.050 334.715 2496.330 335.085 ;
        RECT 2496.120 300.405 2496.260 334.715 ;
        RECT 2496.050 300.035 2496.330 300.405 ;
        RECT 2496.050 275.555 2496.330 275.925 ;
        RECT 2496.120 229.005 2496.260 275.555 ;
        RECT 2496.050 228.635 2496.330 229.005 ;
        RECT 2496.050 227.275 2496.330 227.645 ;
        RECT 2496.120 203.845 2496.260 227.275 ;
        RECT 2496.050 203.475 2496.330 203.845 ;
        RECT 276.090 23.955 276.370 24.325 ;
        RECT 276.160 2.400 276.300 23.955 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 2495.590 503.400 2495.870 503.680 ;
        RECT 2495.590 338.160 2495.870 338.440 ;
        RECT 2496.050 334.760 2496.330 335.040 ;
        RECT 2496.050 300.080 2496.330 300.360 ;
        RECT 2496.050 275.600 2496.330 275.880 ;
        RECT 2496.050 228.680 2496.330 228.960 ;
        RECT 2496.050 227.320 2496.330 227.600 ;
        RECT 2496.050 203.520 2496.330 203.800 ;
        RECT 276.090 24.000 276.370 24.280 ;
      LAYER met3 ;
        RECT 2506.000 1196.840 2510.000 1197.440 ;
        RECT 2509.150 1194.570 2509.450 1196.840 ;
        RECT 2510.030 1194.570 2510.410 1194.580 ;
        RECT 2509.150 1194.270 2510.410 1194.570 ;
        RECT 2510.030 1194.260 2510.410 1194.270 ;
        RECT 2494.390 503.690 2494.770 503.700 ;
        RECT 2495.565 503.690 2495.895 503.705 ;
        RECT 2494.390 503.390 2495.895 503.690 ;
        RECT 2494.390 503.380 2494.770 503.390 ;
        RECT 2495.565 503.375 2495.895 503.390 ;
        RECT 2495.565 338.460 2495.895 338.465 ;
        RECT 2495.310 338.450 2495.895 338.460 ;
        RECT 2495.110 338.150 2495.895 338.450 ;
        RECT 2495.310 338.140 2495.895 338.150 ;
        RECT 2495.565 338.135 2495.895 338.140 ;
        RECT 2495.310 335.050 2495.690 335.060 ;
        RECT 2496.025 335.050 2496.355 335.065 ;
        RECT 2495.310 334.750 2496.355 335.050 ;
        RECT 2495.310 334.740 2495.690 334.750 ;
        RECT 2496.025 334.735 2496.355 334.750 ;
        RECT 2496.025 300.380 2496.355 300.385 ;
        RECT 2496.025 300.370 2496.610 300.380 ;
        RECT 2495.800 300.070 2496.610 300.370 ;
        RECT 2496.025 300.060 2496.610 300.070 ;
        RECT 2496.025 300.055 2496.355 300.060 ;
        RECT 2496.025 275.900 2496.355 275.905 ;
        RECT 2496.025 275.890 2496.610 275.900 ;
        RECT 2495.800 275.590 2496.610 275.890 ;
        RECT 2496.025 275.580 2496.610 275.590 ;
        RECT 2496.025 275.575 2496.355 275.580 ;
        RECT 2496.025 228.980 2496.355 228.985 ;
        RECT 2496.025 228.970 2496.610 228.980 ;
        RECT 2496.025 228.670 2496.810 228.970 ;
        RECT 2496.025 228.660 2496.610 228.670 ;
        RECT 2496.025 228.655 2496.355 228.660 ;
        RECT 2496.025 227.620 2496.355 227.625 ;
        RECT 2496.025 227.610 2496.610 227.620 ;
        RECT 2495.800 227.310 2496.610 227.610 ;
        RECT 2496.025 227.300 2496.610 227.310 ;
        RECT 2496.025 227.295 2496.355 227.300 ;
        RECT 2496.025 203.820 2496.355 203.825 ;
        RECT 2496.025 203.810 2496.610 203.820 ;
        RECT 2496.025 203.510 2496.810 203.810 ;
        RECT 2496.025 203.500 2496.610 203.510 ;
        RECT 2496.025 203.495 2496.355 203.500 ;
        RECT 276.065 24.290 276.395 24.305 ;
        RECT 2496.230 24.290 2496.610 24.300 ;
        RECT 276.065 23.990 2496.610 24.290 ;
        RECT 276.065 23.975 276.395 23.990 ;
        RECT 2496.230 23.980 2496.610 23.990 ;
      LAYER via3 ;
        RECT 2510.060 1194.260 2510.380 1194.580 ;
        RECT 2494.420 503.380 2494.740 503.700 ;
        RECT 2495.340 338.140 2495.660 338.460 ;
        RECT 2495.340 334.740 2495.660 335.060 ;
        RECT 2496.260 300.060 2496.580 300.380 ;
        RECT 2496.260 275.580 2496.580 275.900 ;
        RECT 2496.260 228.660 2496.580 228.980 ;
        RECT 2496.260 227.300 2496.580 227.620 ;
        RECT 2496.260 203.500 2496.580 203.820 ;
        RECT 2496.260 23.980 2496.580 24.300 ;
      LAYER met4 ;
        RECT 2510.055 1194.255 2510.385 1194.585 ;
        RECT 2510.070 1175.290 2510.370 1194.255 ;
        RECT 2494.910 1174.110 2496.090 1175.290 ;
        RECT 2509.630 1174.110 2510.810 1175.290 ;
        RECT 2495.350 1052.450 2495.650 1174.110 ;
        RECT 2495.350 1052.150 2496.570 1052.450 ;
        RECT 2496.270 1049.050 2496.570 1052.150 ;
        RECT 2494.430 1048.750 2496.570 1049.050 ;
        RECT 2494.430 855.250 2494.730 1048.750 ;
        RECT 2494.430 854.950 2495.650 855.250 ;
        RECT 2495.350 811.490 2495.650 854.950 ;
        RECT 2494.910 810.310 2496.090 811.490 ;
        RECT 2493.990 806.910 2495.170 808.090 ;
        RECT 2494.430 774.330 2494.730 806.910 ;
        RECT 2494.430 774.030 2495.650 774.330 ;
        RECT 2495.350 770.250 2495.650 774.030 ;
        RECT 2493.510 769.950 2495.650 770.250 ;
        RECT 2493.510 756.650 2493.810 769.950 ;
        RECT 2493.510 756.350 2494.730 756.650 ;
        RECT 2494.430 740.090 2494.730 756.350 ;
        RECT 2488.470 738.910 2489.650 740.090 ;
        RECT 2493.990 738.910 2495.170 740.090 ;
        RECT 2488.910 719.690 2489.210 738.910 ;
        RECT 2495.350 722.350 2498.410 722.650 ;
        RECT 2495.350 719.690 2495.650 722.350 ;
        RECT 2488.470 718.510 2489.650 719.690 ;
        RECT 2494.910 718.510 2496.090 719.690 ;
        RECT 2498.110 719.250 2498.410 722.350 ;
        RECT 2498.110 718.950 2502.090 719.250 ;
        RECT 2501.790 671.650 2502.090 718.950 ;
        RECT 2500.870 671.350 2502.090 671.650 ;
        RECT 2500.870 654.650 2501.170 671.350 ;
        RECT 2500.870 654.350 2502.090 654.650 ;
        RECT 2501.790 634.690 2502.090 654.350 ;
        RECT 2495.830 633.510 2497.010 634.690 ;
        RECT 2501.350 633.510 2502.530 634.690 ;
        RECT 2496.270 579.850 2496.570 633.510 ;
        RECT 2494.430 579.550 2496.570 579.850 ;
        RECT 2494.430 503.705 2494.730 579.550 ;
        RECT 2494.415 503.375 2494.745 503.705 ;
        RECT 2495.335 338.135 2495.665 338.465 ;
        RECT 2495.350 335.065 2495.650 338.135 ;
        RECT 2495.335 334.735 2495.665 335.065 ;
        RECT 2496.255 300.055 2496.585 300.385 ;
        RECT 2496.270 275.905 2496.570 300.055 ;
        RECT 2496.255 275.575 2496.585 275.905 ;
        RECT 2496.255 228.655 2496.585 228.985 ;
        RECT 2496.270 227.625 2496.570 228.655 ;
        RECT 2496.255 227.295 2496.585 227.625 ;
        RECT 2496.255 203.495 2496.585 203.825 ;
        RECT 2496.270 158.250 2496.570 203.495 ;
        RECT 2495.350 157.950 2496.570 158.250 ;
        RECT 2495.350 110.650 2495.650 157.950 ;
        RECT 2494.430 110.350 2495.650 110.650 ;
        RECT 2494.430 107.250 2494.730 110.350 ;
        RECT 2494.430 106.950 2496.570 107.250 ;
        RECT 2496.270 24.305 2496.570 106.950 ;
        RECT 2496.255 23.975 2496.585 24.305 ;
      LAYER met5 ;
        RECT 2494.700 1173.900 2511.020 1175.500 ;
        RECT 2493.780 810.100 2496.300 811.700 ;
        RECT 2493.780 806.700 2495.380 810.100 ;
        RECT 2488.260 738.700 2495.380 740.300 ;
        RECT 2488.260 718.300 2496.300 719.900 ;
        RECT 2495.620 633.300 2502.740 634.900 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.310 79.800 296.630 79.860 ;
        RECT 1166.170 79.800 1166.490 79.860 ;
        RECT 296.310 79.660 1166.490 79.800 ;
        RECT 296.310 79.600 296.630 79.660 ;
        RECT 1166.170 79.600 1166.490 79.660 ;
        RECT 294.010 17.240 294.330 17.300 ;
        RECT 296.310 17.240 296.630 17.300 ;
        RECT 294.010 17.100 296.630 17.240 ;
        RECT 294.010 17.040 294.330 17.100 ;
        RECT 296.310 17.040 296.630 17.100 ;
      LAYER via ;
        RECT 296.340 79.600 296.600 79.860 ;
        RECT 1166.200 79.600 1166.460 79.860 ;
        RECT 294.040 17.040 294.300 17.300 ;
        RECT 296.340 17.040 296.600 17.300 ;
      LAYER met2 ;
        RECT 1166.330 510.340 1166.610 514.000 ;
        RECT 1166.260 510.000 1166.610 510.340 ;
        RECT 1166.260 79.890 1166.400 510.000 ;
        RECT 296.340 79.570 296.600 79.890 ;
        RECT 1166.200 79.570 1166.460 79.890 ;
        RECT 296.400 17.330 296.540 79.570 ;
        RECT 294.040 17.010 294.300 17.330 ;
        RECT 296.340 17.010 296.600 17.330 ;
        RECT 294.100 2.400 294.240 17.010 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 315.170 1663.180 315.490 1663.240 ;
        RECT 393.370 1663.180 393.690 1663.240 ;
        RECT 315.170 1663.040 393.690 1663.180 ;
        RECT 315.170 1662.980 315.490 1663.040 ;
        RECT 393.370 1662.980 393.690 1663.040 ;
        RECT 311.950 17.580 312.270 17.640 ;
        RECT 315.170 17.580 315.490 17.640 ;
        RECT 311.950 17.440 315.490 17.580 ;
        RECT 311.950 17.380 312.270 17.440 ;
        RECT 315.170 17.380 315.490 17.440 ;
      LAYER via ;
        RECT 315.200 1662.980 315.460 1663.240 ;
        RECT 393.400 1662.980 393.660 1663.240 ;
        RECT 311.980 17.380 312.240 17.640 ;
        RECT 315.200 17.380 315.460 17.640 ;
      LAYER met2 ;
        RECT 393.390 1663.435 393.670 1663.805 ;
        RECT 393.460 1663.270 393.600 1663.435 ;
        RECT 315.200 1662.950 315.460 1663.270 ;
        RECT 393.400 1662.950 393.660 1663.270 ;
        RECT 315.260 17.670 315.400 1662.950 ;
        RECT 311.980 17.350 312.240 17.670 ;
        RECT 315.200 17.350 315.460 17.670 ;
        RECT 312.040 2.400 312.180 17.350 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 393.390 1663.480 393.670 1663.760 ;
      LAYER met3 ;
        RECT 393.365 1663.770 393.695 1663.785 ;
        RECT 410.000 1663.770 414.000 1663.920 ;
        RECT 393.365 1663.470 414.000 1663.770 ;
        RECT 393.365 1663.455 393.695 1663.470 ;
        RECT 410.000 1663.320 414.000 1663.470 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 328.970 1918.520 329.290 1918.580 ;
        RECT 393.370 1918.520 393.690 1918.580 ;
        RECT 328.970 1918.380 393.690 1918.520 ;
        RECT 328.970 1918.320 329.290 1918.380 ;
        RECT 393.370 1918.320 393.690 1918.380 ;
      LAYER via ;
        RECT 329.000 1918.320 329.260 1918.580 ;
        RECT 393.400 1918.320 393.660 1918.580 ;
      LAYER met2 ;
        RECT 393.390 1919.115 393.670 1919.485 ;
        RECT 393.460 1918.610 393.600 1919.115 ;
        RECT 329.000 1918.290 329.260 1918.610 ;
        RECT 393.400 1918.290 393.660 1918.610 ;
        RECT 329.060 16.730 329.200 1918.290 ;
        RECT 329.060 16.590 330.120 16.730 ;
        RECT 329.980 2.400 330.120 16.590 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 393.390 1919.160 393.670 1919.440 ;
      LAYER met3 ;
        RECT 393.365 1919.450 393.695 1919.465 ;
        RECT 410.000 1919.450 414.000 1919.600 ;
        RECT 393.365 1919.150 414.000 1919.450 ;
        RECT 393.365 1919.135 393.695 1919.150 ;
        RECT 410.000 1919.000 414.000 1919.150 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 350.590 1476.860 350.910 1476.920 ;
        RECT 393.370 1476.860 393.690 1476.920 ;
        RECT 350.590 1476.720 393.690 1476.860 ;
        RECT 350.590 1476.660 350.910 1476.720 ;
        RECT 393.370 1476.660 393.690 1476.720 ;
        RECT 347.370 14.520 347.690 14.580 ;
        RECT 350.590 14.520 350.910 14.580 ;
        RECT 347.370 14.380 350.910 14.520 ;
        RECT 347.370 14.320 347.690 14.380 ;
        RECT 350.590 14.320 350.910 14.380 ;
      LAYER via ;
        RECT 350.620 1476.660 350.880 1476.920 ;
        RECT 393.400 1476.660 393.660 1476.920 ;
        RECT 347.400 14.320 347.660 14.580 ;
        RECT 350.620 14.320 350.880 14.580 ;
      LAYER met2 ;
        RECT 393.390 1481.195 393.670 1481.565 ;
        RECT 393.460 1476.950 393.600 1481.195 ;
        RECT 350.620 1476.630 350.880 1476.950 ;
        RECT 393.400 1476.630 393.660 1476.950 ;
        RECT 350.680 14.610 350.820 1476.630 ;
        RECT 347.400 14.290 347.660 14.610 ;
        RECT 350.620 14.290 350.880 14.610 ;
        RECT 347.460 2.400 347.600 14.290 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 393.390 1481.240 393.670 1481.520 ;
      LAYER met3 ;
        RECT 393.365 1481.530 393.695 1481.545 ;
        RECT 410.000 1481.530 414.000 1481.680 ;
        RECT 393.365 1481.230 414.000 1481.530 ;
        RECT 393.365 1481.215 393.695 1481.230 ;
        RECT 410.000 1481.080 414.000 1481.230 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1432.070 3010.515 1432.350 3010.885 ;
        RECT 1432.140 3010.000 1432.280 3010.515 ;
        RECT 1432.140 3009.340 1432.490 3010.000 ;
        RECT 1432.210 3006.000 1432.490 3009.340 ;
        RECT 365.330 17.155 365.610 17.525 ;
        RECT 365.400 2.400 365.540 17.155 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1432.070 3010.560 1432.350 3010.840 ;
        RECT 365.330 17.200 365.610 17.480 ;
      LAYER met3 ;
        RECT 362.750 3010.850 363.130 3010.860 ;
        RECT 1432.045 3010.850 1432.375 3010.865 ;
        RECT 362.750 3010.550 1432.375 3010.850 ;
        RECT 362.750 3010.540 363.130 3010.550 ;
        RECT 1432.045 3010.535 1432.375 3010.550 ;
        RECT 362.750 17.490 363.130 17.500 ;
        RECT 365.305 17.490 365.635 17.505 ;
        RECT 362.750 17.190 365.635 17.490 ;
        RECT 362.750 17.180 363.130 17.190 ;
        RECT 365.305 17.175 365.635 17.190 ;
      LAYER via3 ;
        RECT 362.780 3010.540 363.100 3010.860 ;
        RECT 362.780 17.180 363.100 17.500 ;
      LAYER met4 ;
        RECT 362.775 3010.535 363.105 3010.865 ;
        RECT 362.790 17.505 363.090 3010.535 ;
        RECT 362.775 17.175 363.105 17.505 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 16.900 383.570 16.960 ;
        RECT 386.010 16.900 386.330 16.960 ;
        RECT 383.250 16.760 386.330 16.900 ;
        RECT 383.250 16.700 383.570 16.760 ;
        RECT 386.010 16.700 386.330 16.760 ;
      LAYER via ;
        RECT 383.280 16.700 383.540 16.960 ;
        RECT 386.040 16.700 386.300 16.960 ;
      LAYER met2 ;
        RECT 2383.490 3006.690 2383.770 3010.000 ;
        RECT 2384.730 3006.690 2385.010 3006.805 ;
        RECT 2383.490 3006.550 2385.010 3006.690 ;
        RECT 2383.490 3006.000 2383.770 3006.550 ;
        RECT 2384.730 3006.435 2385.010 3006.550 ;
        RECT 386.030 451.675 386.310 452.045 ;
        RECT 386.100 16.990 386.240 451.675 ;
        RECT 383.280 16.670 383.540 16.990 ;
        RECT 386.040 16.670 386.300 16.990 ;
        RECT 383.340 2.400 383.480 16.670 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 2384.730 3006.480 2385.010 3006.760 ;
        RECT 386.030 451.720 386.310 452.000 ;
      LAYER met3 ;
        RECT 2384.705 3006.780 2385.035 3006.785 ;
        RECT 2384.705 3006.770 2385.290 3006.780 ;
        RECT 2384.705 3006.470 2385.490 3006.770 ;
        RECT 2384.705 3006.460 2385.290 3006.470 ;
        RECT 2384.705 3006.455 2385.035 3006.460 ;
        RECT 386.005 452.010 386.335 452.025 ;
        RECT 2545.910 452.010 2546.290 452.020 ;
        RECT 386.005 451.710 2546.290 452.010 ;
        RECT 386.005 451.695 386.335 451.710 ;
        RECT 2545.910 451.700 2546.290 451.710 ;
      LAYER via3 ;
        RECT 2384.940 3006.460 2385.260 3006.780 ;
        RECT 2545.940 451.700 2546.260 452.020 ;
      LAYER met4 ;
        RECT 2384.935 3006.455 2385.265 3006.785 ;
        RECT 2384.950 3004.490 2385.250 3006.455 ;
        RECT 2384.510 3003.310 2385.690 3004.490 ;
        RECT 2545.510 3003.310 2546.690 3004.490 ;
        RECT 2545.950 452.025 2546.250 3003.310 ;
        RECT 2545.935 451.695 2546.265 452.025 ;
      LAYER met5 ;
        RECT 2384.300 3003.100 2546.900 3004.700 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 321.610 2008.280 321.930 2008.340 ;
        RECT 393.370 2008.280 393.690 2008.340 ;
        RECT 321.610 2008.140 393.690 2008.280 ;
        RECT 321.610 2008.080 321.930 2008.140 ;
        RECT 393.370 2008.080 393.690 2008.140 ;
        RECT 321.610 20.300 321.930 20.360 ;
        RECT 401.190 20.300 401.510 20.360 ;
        RECT 321.610 20.160 401.510 20.300 ;
        RECT 321.610 20.100 321.930 20.160 ;
        RECT 401.190 20.100 401.510 20.160 ;
      LAYER via ;
        RECT 321.640 2008.080 321.900 2008.340 ;
        RECT 393.400 2008.080 393.660 2008.340 ;
        RECT 321.640 20.100 321.900 20.360 ;
        RECT 401.220 20.100 401.480 20.360 ;
      LAYER met2 ;
        RECT 393.390 2011.595 393.670 2011.965 ;
        RECT 393.460 2008.370 393.600 2011.595 ;
        RECT 321.640 2008.050 321.900 2008.370 ;
        RECT 393.400 2008.050 393.660 2008.370 ;
        RECT 321.700 20.390 321.840 2008.050 ;
        RECT 321.640 20.070 321.900 20.390 ;
        RECT 401.220 20.070 401.480 20.390 ;
        RECT 401.280 2.400 401.420 20.070 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 393.390 2011.640 393.670 2011.920 ;
      LAYER met3 ;
        RECT 393.365 2011.930 393.695 2011.945 ;
        RECT 410.000 2011.930 414.000 2012.080 ;
        RECT 393.365 2011.630 414.000 2011.930 ;
        RECT 393.365 2011.615 393.695 2011.630 ;
        RECT 410.000 2011.480 414.000 2011.630 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 731.580 86.410 731.640 ;
        RECT 393.370 731.580 393.690 731.640 ;
        RECT 86.090 731.440 393.690 731.580 ;
        RECT 86.090 731.380 86.410 731.440 ;
        RECT 393.370 731.380 393.690 731.440 ;
        RECT 62.170 22.000 62.490 22.060 ;
        RECT 86.090 22.000 86.410 22.060 ;
        RECT 62.170 21.860 86.410 22.000 ;
        RECT 62.170 21.800 62.490 21.860 ;
        RECT 86.090 21.800 86.410 21.860 ;
      LAYER via ;
        RECT 86.120 731.380 86.380 731.640 ;
        RECT 393.400 731.380 393.660 731.640 ;
        RECT 62.200 21.800 62.460 22.060 ;
        RECT 86.120 21.800 86.380 22.060 ;
      LAYER met2 ;
        RECT 393.390 733.195 393.670 733.565 ;
        RECT 393.460 731.670 393.600 733.195 ;
        RECT 86.120 731.350 86.380 731.670 ;
        RECT 393.400 731.350 393.660 731.670 ;
        RECT 86.180 22.090 86.320 731.350 ;
        RECT 62.200 21.770 62.460 22.090 ;
        RECT 86.120 21.770 86.380 22.090 ;
        RECT 62.260 2.400 62.400 21.770 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 393.390 733.240 393.670 733.520 ;
      LAYER met3 ;
        RECT 393.365 733.530 393.695 733.545 ;
        RECT 410.000 733.530 414.000 733.680 ;
        RECT 393.365 733.230 414.000 733.530 ;
        RECT 393.365 733.215 393.695 733.230 ;
        RECT 410.000 733.080 414.000 733.230 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.530 375.515 420.810 375.885 ;
        RECT 420.600 17.410 420.740 375.515 ;
        RECT 419.220 17.270 420.740 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 420.530 375.560 420.810 375.840 ;
      LAYER met3 ;
        RECT 2506.000 776.600 2510.000 777.200 ;
        RECT 2507.310 774.340 2507.610 776.600 ;
        RECT 2507.270 774.020 2507.650 774.340 ;
        RECT 2498.070 387.410 2498.450 387.420 ;
        RECT 2497.190 387.110 2498.450 387.410 ;
        RECT 2497.190 386.740 2497.490 387.110 ;
        RECT 2498.070 387.100 2498.450 387.110 ;
        RECT 2497.150 386.420 2497.530 386.740 ;
        RECT 420.505 375.850 420.835 375.865 ;
        RECT 2497.150 375.850 2497.530 375.860 ;
        RECT 420.505 375.550 2497.530 375.850 ;
        RECT 420.505 375.535 420.835 375.550 ;
        RECT 2497.150 375.540 2497.530 375.550 ;
      LAYER via3 ;
        RECT 2507.300 774.020 2507.620 774.340 ;
        RECT 2498.100 387.100 2498.420 387.420 ;
        RECT 2497.180 386.420 2497.500 386.740 ;
        RECT 2497.180 375.540 2497.500 375.860 ;
      LAYER met4 ;
        RECT 2507.295 774.015 2507.625 774.345 ;
        RECT 2507.310 760.490 2507.610 774.015 ;
        RECT 2496.750 759.310 2497.930 760.490 ;
        RECT 2506.870 759.310 2508.050 760.490 ;
        RECT 2497.190 736.690 2497.490 759.310 ;
        RECT 2490.310 735.510 2491.490 736.690 ;
        RECT 2496.750 735.510 2497.930 736.690 ;
        RECT 2490.750 716.290 2491.050 735.510 ;
        RECT 2490.310 715.110 2491.490 716.290 ;
        RECT 2494.910 715.110 2496.090 716.290 ;
        RECT 2495.350 712.450 2495.650 715.110 ;
        RECT 2495.350 712.150 2497.490 712.450 ;
        RECT 2497.190 647.850 2497.490 712.150 ;
        RECT 2496.270 647.550 2497.490 647.850 ;
        RECT 2496.270 641.050 2496.570 647.550 ;
        RECT 2496.270 640.750 2498.410 641.050 ;
        RECT 2498.110 624.050 2498.410 640.750 ;
        RECT 2497.190 623.750 2498.410 624.050 ;
        RECT 2497.190 433.650 2497.490 623.750 ;
        RECT 2497.190 433.350 2498.410 433.650 ;
        RECT 2498.110 387.425 2498.410 433.350 ;
        RECT 2498.095 387.095 2498.425 387.425 ;
        RECT 2497.175 386.415 2497.505 386.745 ;
        RECT 2497.190 375.865 2497.490 386.415 ;
        RECT 2497.175 375.535 2497.505 375.865 ;
      LAYER met5 ;
        RECT 2496.540 759.100 2508.260 760.700 ;
        RECT 2490.100 735.300 2498.140 736.900 ;
        RECT 2490.100 714.900 2496.300 716.500 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2215.000 2519.810 2215.060 ;
        RECT 2548.010 2215.000 2548.330 2215.060 ;
        RECT 2519.490 2214.860 2548.330 2215.000 ;
        RECT 2519.490 2214.800 2519.810 2214.860 ;
        RECT 2548.010 2214.800 2548.330 2214.860 ;
        RECT 441.210 320.860 441.530 320.920 ;
        RECT 2548.010 320.860 2548.330 320.920 ;
        RECT 441.210 320.720 2548.330 320.860 ;
        RECT 441.210 320.660 441.530 320.720 ;
        RECT 2548.010 320.660 2548.330 320.720 ;
        RECT 436.610 16.900 436.930 16.960 ;
        RECT 441.210 16.900 441.530 16.960 ;
        RECT 436.610 16.760 441.530 16.900 ;
        RECT 436.610 16.700 436.930 16.760 ;
        RECT 441.210 16.700 441.530 16.760 ;
      LAYER via ;
        RECT 2519.520 2214.800 2519.780 2215.060 ;
        RECT 2548.040 2214.800 2548.300 2215.060 ;
        RECT 441.240 320.660 441.500 320.920 ;
        RECT 2548.040 320.660 2548.300 320.920 ;
        RECT 436.640 16.700 436.900 16.960 ;
        RECT 441.240 16.700 441.500 16.960 ;
      LAYER met2 ;
        RECT 2519.510 2219.675 2519.790 2220.045 ;
        RECT 2519.580 2215.090 2519.720 2219.675 ;
        RECT 2519.520 2214.770 2519.780 2215.090 ;
        RECT 2548.040 2214.770 2548.300 2215.090 ;
        RECT 2548.100 320.950 2548.240 2214.770 ;
        RECT 441.240 320.630 441.500 320.950 ;
        RECT 2548.040 320.630 2548.300 320.950 ;
        RECT 441.300 16.990 441.440 320.630 ;
        RECT 436.640 16.670 436.900 16.990 ;
        RECT 441.240 16.670 441.500 16.990 ;
        RECT 436.700 2.400 436.840 16.670 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2219.720 2519.790 2220.000 ;
      LAYER met3 ;
        RECT 2506.000 2220.010 2510.000 2220.160 ;
        RECT 2519.485 2220.010 2519.815 2220.025 ;
        RECT 2506.000 2219.710 2519.815 2220.010 ;
        RECT 2506.000 2219.560 2510.000 2219.710 ;
        RECT 2519.485 2219.695 2519.815 2219.710 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 449.565 241.485 449.735 289.595 ;
        RECT 450.025 145.265 450.195 159.035 ;
        RECT 449.105 109.565 449.275 137.955 ;
      LAYER mcon ;
        RECT 449.565 289.425 449.735 289.595 ;
        RECT 450.025 158.865 450.195 159.035 ;
        RECT 449.105 137.785 449.275 137.955 ;
      LAYER met1 ;
        RECT 449.490 410.620 449.810 410.680 ;
        RECT 450.410 410.620 450.730 410.680 ;
        RECT 449.490 410.480 450.730 410.620 ;
        RECT 449.490 410.420 449.810 410.480 ;
        RECT 450.410 410.420 450.730 410.480 ;
        RECT 449.490 352.140 449.810 352.200 ;
        RECT 449.120 352.000 449.810 352.140 ;
        RECT 449.120 351.180 449.260 352.000 ;
        RECT 449.490 351.940 449.810 352.000 ;
        RECT 449.030 350.920 449.350 351.180 ;
        RECT 449.030 303.660 449.350 303.920 ;
        RECT 449.120 303.520 449.260 303.660 ;
        RECT 449.950 303.520 450.270 303.580 ;
        RECT 449.120 303.380 450.270 303.520 ;
        RECT 449.950 303.320 450.270 303.380 ;
        RECT 449.505 289.580 449.795 289.625 ;
        RECT 449.950 289.580 450.270 289.640 ;
        RECT 449.505 289.440 450.270 289.580 ;
        RECT 449.505 289.395 449.795 289.440 ;
        RECT 449.950 289.380 450.270 289.440 ;
        RECT 449.490 241.640 449.810 241.700 ;
        RECT 449.295 241.500 449.810 241.640 ;
        RECT 449.490 241.440 449.810 241.500 ;
        RECT 449.030 206.960 449.350 207.020 ;
        RECT 449.950 206.960 450.270 207.020 ;
        RECT 449.030 206.820 450.270 206.960 ;
        RECT 449.030 206.760 449.350 206.820 ;
        RECT 449.950 206.760 450.270 206.820 ;
        RECT 449.950 159.020 450.270 159.080 ;
        RECT 449.755 158.880 450.270 159.020 ;
        RECT 449.950 158.820 450.270 158.880 ;
        RECT 449.490 145.420 449.810 145.480 ;
        RECT 449.965 145.420 450.255 145.465 ;
        RECT 449.490 145.280 450.255 145.420 ;
        RECT 449.490 145.220 449.810 145.280 ;
        RECT 449.965 145.235 450.255 145.280 ;
        RECT 449.030 137.940 449.350 138.000 ;
        RECT 448.835 137.800 449.350 137.940 ;
        RECT 449.030 137.740 449.350 137.800 ;
        RECT 449.045 109.720 449.335 109.765 ;
        RECT 449.950 109.720 450.270 109.780 ;
        RECT 449.045 109.580 450.270 109.720 ;
        RECT 449.045 109.535 449.335 109.580 ;
        RECT 449.950 109.520 450.270 109.580 ;
        RECT 449.950 16.220 450.270 16.280 ;
        RECT 454.550 16.220 454.870 16.280 ;
        RECT 449.950 16.080 454.870 16.220 ;
        RECT 449.950 16.020 450.270 16.080 ;
        RECT 454.550 16.020 454.870 16.080 ;
      LAYER via ;
        RECT 449.520 410.420 449.780 410.680 ;
        RECT 450.440 410.420 450.700 410.680 ;
        RECT 449.520 351.940 449.780 352.200 ;
        RECT 449.060 350.920 449.320 351.180 ;
        RECT 449.060 303.660 449.320 303.920 ;
        RECT 449.980 303.320 450.240 303.580 ;
        RECT 449.980 289.380 450.240 289.640 ;
        RECT 449.520 241.440 449.780 241.700 ;
        RECT 449.060 206.760 449.320 207.020 ;
        RECT 449.980 206.760 450.240 207.020 ;
        RECT 449.980 158.820 450.240 159.080 ;
        RECT 449.520 145.220 449.780 145.480 ;
        RECT 449.060 137.740 449.320 138.000 ;
        RECT 449.980 109.520 450.240 109.780 ;
        RECT 449.980 16.020 450.240 16.280 ;
        RECT 454.580 16.020 454.840 16.280 ;
      LAYER met2 ;
        RECT 403.510 3006.435 403.790 3006.805 ;
        RECT 1393.890 3006.690 1394.170 3006.805 ;
        RECT 1395.410 3006.690 1395.690 3010.000 ;
        RECT 1393.890 3006.550 1395.690 3006.690 ;
        RECT 1393.890 3006.435 1394.170 3006.550 ;
        RECT 295.870 3005.075 296.150 3005.445 ;
        RECT 295.940 508.485 296.080 3005.075 ;
        RECT 403.580 3004.765 403.720 3006.435 ;
        RECT 1395.410 3006.000 1395.690 3006.550 ;
        RECT 403.510 3004.395 403.790 3004.765 ;
        RECT 295.870 508.115 296.150 508.485 ;
        RECT 449.970 508.115 450.250 508.485 ;
        RECT 450.040 448.530 450.180 508.115 ;
        RECT 449.580 448.390 450.180 448.530 ;
        RECT 449.580 410.710 449.720 448.390 ;
        RECT 449.520 410.390 449.780 410.710 ;
        RECT 450.440 410.390 450.700 410.710 ;
        RECT 450.500 386.765 450.640 410.390 ;
        RECT 449.510 386.650 449.790 386.765 ;
        RECT 449.120 386.510 449.790 386.650 ;
        RECT 449.120 385.970 449.260 386.510 ;
        RECT 449.510 386.395 449.790 386.510 ;
        RECT 450.430 386.395 450.710 386.765 ;
        RECT 449.120 385.830 449.720 385.970 ;
        RECT 449.580 352.230 449.720 385.830 ;
        RECT 449.520 351.910 449.780 352.230 ;
        RECT 449.060 350.890 449.320 351.210 ;
        RECT 449.120 303.950 449.260 350.890 ;
        RECT 449.060 303.630 449.320 303.950 ;
        RECT 449.980 303.290 450.240 303.610 ;
        RECT 450.040 289.670 450.180 303.290 ;
        RECT 449.980 289.350 450.240 289.670 ;
        RECT 449.520 241.410 449.780 241.730 ;
        RECT 449.580 207.130 449.720 241.410 ;
        RECT 449.120 207.050 449.720 207.130 ;
        RECT 449.060 206.990 449.720 207.050 ;
        RECT 449.060 206.730 449.320 206.990 ;
        RECT 449.980 206.730 450.240 207.050 ;
        RECT 450.040 159.110 450.180 206.730 ;
        RECT 449.980 158.790 450.240 159.110 ;
        RECT 449.520 145.250 449.780 145.510 ;
        RECT 449.120 145.190 449.780 145.250 ;
        RECT 449.120 145.110 449.720 145.190 ;
        RECT 449.120 138.030 449.260 145.110 ;
        RECT 449.060 137.710 449.320 138.030 ;
        RECT 449.980 109.490 450.240 109.810 ;
        RECT 450.040 16.310 450.180 109.490 ;
        RECT 449.980 15.990 450.240 16.310 ;
        RECT 454.580 15.990 454.840 16.310 ;
        RECT 454.640 2.400 454.780 15.990 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 403.510 3006.480 403.790 3006.760 ;
        RECT 1393.890 3006.480 1394.170 3006.760 ;
        RECT 295.870 3005.120 296.150 3005.400 ;
        RECT 403.510 3004.440 403.790 3004.720 ;
        RECT 295.870 508.160 296.150 508.440 ;
        RECT 449.970 508.160 450.250 508.440 ;
        RECT 449.510 386.440 449.790 386.720 ;
        RECT 450.430 386.440 450.710 386.720 ;
      LAYER met3 ;
        RECT 379.310 3006.770 379.690 3006.780 ;
        RECT 403.485 3006.770 403.815 3006.785 ;
        RECT 379.310 3006.470 403.815 3006.770 ;
        RECT 379.310 3006.460 379.690 3006.470 ;
        RECT 403.485 3006.455 403.815 3006.470 ;
        RECT 1303.910 3006.770 1304.290 3006.780 ;
        RECT 1351.750 3006.770 1352.130 3006.780 ;
        RECT 1303.910 3006.470 1352.130 3006.770 ;
        RECT 1303.910 3006.460 1304.290 3006.470 ;
        RECT 1351.750 3006.460 1352.130 3006.470 ;
        RECT 1352.670 3006.770 1353.050 3006.780 ;
        RECT 1393.865 3006.770 1394.195 3006.785 ;
        RECT 1352.670 3006.470 1394.195 3006.770 ;
        RECT 1352.670 3006.460 1353.050 3006.470 ;
        RECT 1393.865 3006.455 1394.195 3006.470 ;
        RECT 434.510 3006.090 434.890 3006.100 ;
        RECT 675.550 3006.090 675.930 3006.100 ;
        RECT 765.710 3006.090 766.090 3006.100 ;
        RECT 434.510 3005.790 435.770 3006.090 ;
        RECT 434.510 3005.780 434.890 3005.790 ;
        RECT 295.845 3005.410 296.175 3005.425 ;
        RECT 379.310 3005.410 379.690 3005.420 ;
        RECT 295.845 3005.110 379.690 3005.410 ;
        RECT 435.470 3005.410 435.770 3005.790 ;
        RECT 675.550 3005.790 676.810 3006.090 ;
        RECT 675.550 3005.780 675.930 3005.790 ;
        RECT 621.270 3005.410 621.650 3005.420 ;
        RECT 676.510 3005.410 676.810 3005.790 ;
        RECT 765.710 3005.790 790.890 3006.090 ;
        RECT 765.710 3005.780 766.090 3005.790 ;
        RECT 790.590 3005.410 790.890 3005.790 ;
        RECT 879.830 3005.790 883.810 3006.090 ;
        RECT 879.830 3005.410 880.130 3005.790 ;
        RECT 435.470 3005.110 565.490 3005.410 ;
        RECT 295.845 3005.095 296.175 3005.110 ;
        RECT 379.310 3005.100 379.690 3005.110 ;
        RECT 403.485 3004.730 403.815 3004.745 ;
        RECT 434.510 3004.730 434.890 3004.740 ;
        RECT 403.485 3004.430 434.890 3004.730 ;
        RECT 565.190 3004.730 565.490 3005.110 ;
        RECT 621.270 3005.110 662.090 3005.410 ;
        RECT 676.510 3005.110 748.570 3005.410 ;
        RECT 790.590 3005.110 880.130 3005.410 ;
        RECT 883.510 3005.410 883.810 3005.790 ;
        RECT 1076.670 3005.410 1077.050 3005.420 ;
        RECT 1173.270 3005.410 1173.650 3005.420 ;
        RECT 1269.870 3005.410 1270.250 3005.420 ;
        RECT 1303.910 3005.410 1304.290 3005.420 ;
        RECT 883.510 3005.110 940.850 3005.410 ;
        RECT 621.270 3005.100 621.650 3005.110 ;
        RECT 620.350 3004.730 620.730 3004.740 ;
        RECT 565.190 3004.430 620.730 3004.730 ;
        RECT 661.790 3004.730 662.090 3005.110 ;
        RECT 675.550 3004.730 675.930 3004.740 ;
        RECT 661.790 3004.430 675.930 3004.730 ;
        RECT 748.270 3004.730 748.570 3005.110 ;
        RECT 765.710 3004.730 766.090 3004.740 ;
        RECT 748.270 3004.430 766.090 3004.730 ;
        RECT 940.550 3004.730 940.850 3005.110 ;
        RECT 1027.950 3005.110 1029.170 3005.410 ;
        RECT 979.150 3004.730 979.530 3004.740 ;
        RECT 940.550 3004.430 979.530 3004.730 ;
        RECT 403.485 3004.415 403.815 3004.430 ;
        RECT 434.510 3004.420 434.890 3004.430 ;
        RECT 620.350 3004.420 620.730 3004.430 ;
        RECT 675.550 3004.420 675.930 3004.430 ;
        RECT 765.710 3004.420 766.090 3004.430 ;
        RECT 979.150 3004.420 979.530 3004.430 ;
        RECT 1014.110 3004.730 1014.490 3004.740 ;
        RECT 1027.950 3004.730 1028.250 3005.110 ;
        RECT 1014.110 3004.430 1028.250 3004.730 ;
        RECT 1028.870 3004.730 1029.170 3005.110 ;
        RECT 1076.670 3005.110 1134.970 3005.410 ;
        RECT 1076.670 3005.100 1077.050 3005.110 ;
        RECT 1075.750 3004.730 1076.130 3004.740 ;
        RECT 1028.870 3004.430 1076.130 3004.730 ;
        RECT 1134.670 3004.730 1134.970 3005.110 ;
        RECT 1173.270 3005.110 1231.570 3005.410 ;
        RECT 1173.270 3005.100 1173.650 3005.110 ;
        RECT 1172.350 3004.730 1172.730 3004.740 ;
        RECT 1134.670 3004.430 1172.730 3004.730 ;
        RECT 1231.270 3004.730 1231.570 3005.110 ;
        RECT 1269.870 3005.110 1304.290 3005.410 ;
        RECT 1269.870 3005.100 1270.250 3005.110 ;
        RECT 1303.910 3005.100 1304.290 3005.110 ;
        RECT 1351.750 3005.100 1352.130 3005.420 ;
        RECT 1268.950 3004.730 1269.330 3004.740 ;
        RECT 1231.270 3004.430 1269.330 3004.730 ;
        RECT 1351.790 3004.730 1352.090 3005.100 ;
        RECT 1352.670 3004.730 1353.050 3004.740 ;
        RECT 1351.790 3004.430 1353.050 3004.730 ;
        RECT 1014.110 3004.420 1014.490 3004.430 ;
        RECT 1075.750 3004.420 1076.130 3004.430 ;
        RECT 1172.350 3004.420 1172.730 3004.430 ;
        RECT 1268.950 3004.420 1269.330 3004.430 ;
        RECT 1352.670 3004.420 1353.050 3004.430 ;
        RECT 979.150 3001.330 979.530 3001.340 ;
        RECT 1013.190 3001.330 1013.570 3001.340 ;
        RECT 979.150 3001.030 1013.570 3001.330 ;
        RECT 979.150 3001.020 979.530 3001.030 ;
        RECT 1013.190 3001.020 1013.570 3001.030 ;
        RECT 295.845 508.450 296.175 508.465 ;
        RECT 449.945 508.450 450.275 508.465 ;
        RECT 295.845 508.150 450.275 508.450 ;
        RECT 295.845 508.135 296.175 508.150 ;
        RECT 449.945 508.135 450.275 508.150 ;
        RECT 449.485 386.730 449.815 386.745 ;
        RECT 450.405 386.730 450.735 386.745 ;
        RECT 449.485 386.430 450.735 386.730 ;
        RECT 449.485 386.415 449.815 386.430 ;
        RECT 450.405 386.415 450.735 386.430 ;
      LAYER via3 ;
        RECT 379.340 3006.460 379.660 3006.780 ;
        RECT 1303.940 3006.460 1304.260 3006.780 ;
        RECT 1351.780 3006.460 1352.100 3006.780 ;
        RECT 1352.700 3006.460 1353.020 3006.780 ;
        RECT 434.540 3005.780 434.860 3006.100 ;
        RECT 379.340 3005.100 379.660 3005.420 ;
        RECT 675.580 3005.780 675.900 3006.100 ;
        RECT 434.540 3004.420 434.860 3004.740 ;
        RECT 621.300 3005.100 621.620 3005.420 ;
        RECT 765.740 3005.780 766.060 3006.100 ;
        RECT 620.380 3004.420 620.700 3004.740 ;
        RECT 675.580 3004.420 675.900 3004.740 ;
        RECT 765.740 3004.420 766.060 3004.740 ;
        RECT 979.180 3004.420 979.500 3004.740 ;
        RECT 1014.140 3004.420 1014.460 3004.740 ;
        RECT 1076.700 3005.100 1077.020 3005.420 ;
        RECT 1075.780 3004.420 1076.100 3004.740 ;
        RECT 1173.300 3005.100 1173.620 3005.420 ;
        RECT 1172.380 3004.420 1172.700 3004.740 ;
        RECT 1269.900 3005.100 1270.220 3005.420 ;
        RECT 1303.940 3005.100 1304.260 3005.420 ;
        RECT 1351.780 3005.100 1352.100 3005.420 ;
        RECT 1268.980 3004.420 1269.300 3004.740 ;
        RECT 1352.700 3004.420 1353.020 3004.740 ;
        RECT 979.180 3001.020 979.500 3001.340 ;
        RECT 1013.220 3001.020 1013.540 3001.340 ;
      LAYER met4 ;
        RECT 379.335 3006.455 379.665 3006.785 ;
        RECT 1303.935 3006.455 1304.265 3006.785 ;
        RECT 1351.775 3006.455 1352.105 3006.785 ;
        RECT 1352.695 3006.455 1353.025 3006.785 ;
        RECT 379.350 3005.425 379.650 3006.455 ;
        RECT 434.535 3005.775 434.865 3006.105 ;
        RECT 675.575 3005.775 675.905 3006.105 ;
        RECT 765.735 3005.775 766.065 3006.105 ;
        RECT 379.335 3005.095 379.665 3005.425 ;
        RECT 434.550 3004.745 434.850 3005.775 ;
        RECT 621.295 3005.095 621.625 3005.425 ;
        RECT 434.535 3004.415 434.865 3004.745 ;
        RECT 620.375 3004.415 620.705 3004.745 ;
        RECT 620.390 3004.050 620.690 3004.415 ;
        RECT 621.310 3004.050 621.610 3005.095 ;
        RECT 675.590 3004.745 675.890 3005.775 ;
        RECT 765.750 3004.745 766.050 3005.775 ;
        RECT 1303.950 3005.425 1304.250 3006.455 ;
        RECT 1351.790 3005.425 1352.090 3006.455 ;
        RECT 1076.695 3005.095 1077.025 3005.425 ;
        RECT 1173.295 3005.095 1173.625 3005.425 ;
        RECT 1269.895 3005.095 1270.225 3005.425 ;
        RECT 1303.935 3005.095 1304.265 3005.425 ;
        RECT 1351.775 3005.095 1352.105 3005.425 ;
        RECT 675.575 3004.415 675.905 3004.745 ;
        RECT 765.735 3004.415 766.065 3004.745 ;
        RECT 979.175 3004.415 979.505 3004.745 ;
        RECT 1014.135 3004.415 1014.465 3004.745 ;
        RECT 1075.775 3004.415 1076.105 3004.745 ;
        RECT 620.390 3003.750 621.610 3004.050 ;
        RECT 979.190 3001.345 979.490 3004.415 ;
        RECT 1014.150 3004.050 1014.450 3004.415 ;
        RECT 1013.230 3003.750 1014.450 3004.050 ;
        RECT 1075.790 3004.050 1076.090 3004.415 ;
        RECT 1076.710 3004.050 1077.010 3005.095 ;
        RECT 1172.375 3004.415 1172.705 3004.745 ;
        RECT 1075.790 3003.750 1077.010 3004.050 ;
        RECT 1172.390 3004.050 1172.690 3004.415 ;
        RECT 1173.310 3004.050 1173.610 3005.095 ;
        RECT 1268.975 3004.415 1269.305 3004.745 ;
        RECT 1172.390 3003.750 1173.610 3004.050 ;
        RECT 1268.990 3004.050 1269.290 3004.415 ;
        RECT 1269.910 3004.050 1270.210 3005.095 ;
        RECT 1352.710 3004.745 1353.010 3006.455 ;
        RECT 1352.695 3004.415 1353.025 3004.745 ;
        RECT 1268.990 3003.750 1270.210 3004.050 ;
        RECT 1013.230 3001.345 1013.530 3003.750 ;
        RECT 979.175 3001.015 979.505 3001.345 ;
        RECT 1013.215 3001.015 1013.545 3001.345 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 3017.060 336.190 3017.120 ;
        RECT 1012.530 3017.060 1012.850 3017.120 ;
        RECT 335.870 3016.920 1012.850 3017.060 ;
        RECT 335.870 3016.860 336.190 3016.920 ;
        RECT 1012.530 3016.860 1012.850 3016.920 ;
        RECT 335.870 508.880 336.190 508.940 ;
        RECT 469.730 508.880 470.050 508.940 ;
        RECT 335.870 508.740 470.050 508.880 ;
        RECT 335.870 508.680 336.190 508.740 ;
        RECT 469.730 508.680 470.050 508.740 ;
        RECT 469.730 16.900 470.050 16.960 ;
        RECT 472.490 16.900 472.810 16.960 ;
        RECT 469.730 16.760 472.810 16.900 ;
        RECT 469.730 16.700 470.050 16.760 ;
        RECT 472.490 16.700 472.810 16.760 ;
      LAYER via ;
        RECT 335.900 3016.860 336.160 3017.120 ;
        RECT 1012.560 3016.860 1012.820 3017.120 ;
        RECT 335.900 508.680 336.160 508.940 ;
        RECT 469.760 508.680 470.020 508.940 ;
        RECT 469.760 16.700 470.020 16.960 ;
        RECT 472.520 16.700 472.780 16.960 ;
      LAYER met2 ;
        RECT 335.900 3016.830 336.160 3017.150 ;
        RECT 1012.560 3016.830 1012.820 3017.150 ;
        RECT 335.960 508.970 336.100 3016.830 ;
        RECT 1012.620 3010.000 1012.760 3016.830 ;
        RECT 1012.620 3009.340 1012.970 3010.000 ;
        RECT 1012.690 3006.000 1012.970 3009.340 ;
        RECT 335.900 508.650 336.160 508.970 ;
        RECT 469.760 508.650 470.020 508.970 ;
        RECT 469.820 16.990 469.960 508.650 ;
        RECT 469.760 16.670 470.020 16.990 ;
        RECT 472.520 16.670 472.780 16.990 ;
        RECT 472.580 2.400 472.720 16.670 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2201.400 2519.810 2201.460 ;
        RECT 2547.550 2201.400 2547.870 2201.460 ;
        RECT 2519.490 2201.260 2547.870 2201.400 ;
        RECT 2519.490 2201.200 2519.810 2201.260 ;
        RECT 2547.550 2201.200 2547.870 2201.260 ;
        RECT 496.410 306.920 496.730 306.980 ;
        RECT 2547.550 306.920 2547.870 306.980 ;
        RECT 496.410 306.780 2547.870 306.920 ;
        RECT 496.410 306.720 496.730 306.780 ;
        RECT 2547.550 306.720 2547.870 306.780 ;
        RECT 490.430 16.900 490.750 16.960 ;
        RECT 496.870 16.900 497.190 16.960 ;
        RECT 490.430 16.760 497.190 16.900 ;
        RECT 490.430 16.700 490.750 16.760 ;
        RECT 496.870 16.700 497.190 16.760 ;
      LAYER via ;
        RECT 2519.520 2201.200 2519.780 2201.460 ;
        RECT 2547.580 2201.200 2547.840 2201.460 ;
        RECT 496.440 306.720 496.700 306.980 ;
        RECT 2547.580 306.720 2547.840 306.980 ;
        RECT 490.460 16.700 490.720 16.960 ;
        RECT 496.900 16.700 497.160 16.960 ;
      LAYER met2 ;
        RECT 2519.510 2201.995 2519.790 2202.365 ;
        RECT 2519.580 2201.490 2519.720 2201.995 ;
        RECT 2519.520 2201.170 2519.780 2201.490 ;
        RECT 2547.580 2201.170 2547.840 2201.490 ;
        RECT 2547.640 307.010 2547.780 2201.170 ;
        RECT 496.440 306.690 496.700 307.010 ;
        RECT 2547.580 306.690 2547.840 307.010 ;
        RECT 496.500 18.090 496.640 306.690 ;
        RECT 496.500 17.950 497.100 18.090 ;
        RECT 496.960 16.990 497.100 17.950 ;
        RECT 490.460 16.670 490.720 16.990 ;
        RECT 496.900 16.670 497.160 16.990 ;
        RECT 490.520 2.400 490.660 16.670 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2202.040 2519.790 2202.320 ;
      LAYER met3 ;
        RECT 2506.000 2202.330 2510.000 2202.480 ;
        RECT 2519.485 2202.330 2519.815 2202.345 ;
        RECT 2506.000 2202.030 2519.815 2202.330 ;
        RECT 2506.000 2201.880 2510.000 2202.030 ;
        RECT 2519.485 2202.015 2519.815 2202.030 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1307.390 500.720 1307.710 500.780 ;
        RECT 1968.410 500.720 1968.730 500.780 ;
        RECT 1307.390 500.580 1968.730 500.720 ;
        RECT 1307.390 500.520 1307.710 500.580 ;
        RECT 1968.410 500.520 1968.730 500.580 ;
        RECT 510.210 424.220 510.530 424.280 ;
        RECT 1307.390 424.220 1307.710 424.280 ;
        RECT 510.210 424.080 1307.710 424.220 ;
        RECT 510.210 424.020 510.530 424.080 ;
        RECT 1307.390 424.020 1307.710 424.080 ;
        RECT 507.910 16.900 508.230 16.960 ;
        RECT 510.210 16.900 510.530 16.960 ;
        RECT 507.910 16.760 510.530 16.900 ;
        RECT 507.910 16.700 508.230 16.760 ;
        RECT 510.210 16.700 510.530 16.760 ;
      LAYER via ;
        RECT 1307.420 500.520 1307.680 500.780 ;
        RECT 1968.440 500.520 1968.700 500.780 ;
        RECT 510.240 424.020 510.500 424.280 ;
        RECT 1307.420 424.020 1307.680 424.280 ;
        RECT 507.940 16.700 508.200 16.960 ;
        RECT 510.240 16.700 510.500 16.960 ;
      LAYER met2 ;
        RECT 1968.570 510.340 1968.850 514.000 ;
        RECT 1968.500 510.000 1968.850 510.340 ;
        RECT 1968.500 500.810 1968.640 510.000 ;
        RECT 1307.420 500.490 1307.680 500.810 ;
        RECT 1968.440 500.490 1968.700 500.810 ;
        RECT 1307.480 424.310 1307.620 500.490 ;
        RECT 510.240 423.990 510.500 424.310 ;
        RECT 1307.420 423.990 1307.680 424.310 ;
        RECT 510.300 16.990 510.440 423.990 ;
        RECT 507.940 16.670 508.200 16.990 ;
        RECT 510.240 16.670 510.500 16.990 ;
        RECT 508.000 2.400 508.140 16.670 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 327.660 531.230 327.720 ;
        RECT 1041.970 327.660 1042.290 327.720 ;
        RECT 530.910 327.520 1042.290 327.660 ;
        RECT 530.910 327.460 531.230 327.520 ;
        RECT 1041.970 327.460 1042.290 327.520 ;
        RECT 525.850 16.900 526.170 16.960 ;
        RECT 530.910 16.900 531.230 16.960 ;
        RECT 525.850 16.760 531.230 16.900 ;
        RECT 525.850 16.700 526.170 16.760 ;
        RECT 530.910 16.700 531.230 16.760 ;
      LAYER via ;
        RECT 530.940 327.460 531.200 327.720 ;
        RECT 1042.000 327.460 1042.260 327.720 ;
        RECT 525.880 16.700 526.140 16.960 ;
        RECT 530.940 16.700 531.200 16.960 ;
      LAYER met2 ;
        RECT 1042.130 510.340 1042.410 514.000 ;
        RECT 1042.060 510.000 1042.410 510.340 ;
        RECT 1042.060 327.750 1042.200 510.000 ;
        RECT 530.940 327.430 531.200 327.750 ;
        RECT 1042.000 327.430 1042.260 327.750 ;
        RECT 531.000 16.990 531.140 327.430 ;
        RECT 525.880 16.670 526.140 16.990 ;
        RECT 530.940 16.670 531.200 16.990 ;
        RECT 525.940 2.400 526.080 16.670 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 414.145 554.965 414.315 621.095 ;
      LAYER mcon ;
        RECT 414.145 620.925 414.315 621.095 ;
      LAYER met1 ;
        RECT 414.530 663.240 414.850 663.300 ;
        RECT 414.530 663.100 415.220 663.240 ;
        RECT 414.530 663.040 414.850 663.100 ;
        RECT 412.690 662.560 413.010 662.620 ;
        RECT 415.080 662.560 415.220 663.100 ;
        RECT 412.690 662.420 415.220 662.560 ;
        RECT 412.690 662.360 413.010 662.420 ;
        RECT 414.085 621.080 414.375 621.125 ;
        RECT 414.530 621.080 414.850 621.140 ;
        RECT 414.085 620.940 414.850 621.080 ;
        RECT 414.085 620.895 414.375 620.940 ;
        RECT 414.530 620.880 414.850 620.940 ;
        RECT 414.085 555.120 414.375 555.165 ;
        RECT 414.530 555.120 414.850 555.180 ;
        RECT 414.085 554.980 414.850 555.120 ;
        RECT 414.085 554.935 414.375 554.980 ;
        RECT 414.530 554.920 414.850 554.980 ;
        RECT 415.450 512.280 415.770 512.340 ;
        RECT 418.210 512.280 418.530 512.340 ;
        RECT 415.450 512.140 418.530 512.280 ;
        RECT 415.450 512.080 415.770 512.140 ;
        RECT 418.210 512.080 418.530 512.140 ;
        RECT 418.210 509.220 418.530 509.280 ;
        RECT 538.270 509.220 538.590 509.280 ;
        RECT 418.210 509.080 538.590 509.220 ;
        RECT 418.210 509.020 418.530 509.080 ;
        RECT 538.270 509.020 538.590 509.080 ;
      LAYER via ;
        RECT 414.560 663.040 414.820 663.300 ;
        RECT 412.720 662.360 412.980 662.620 ;
        RECT 414.560 620.880 414.820 621.140 ;
        RECT 414.560 554.920 414.820 555.180 ;
        RECT 415.480 512.080 415.740 512.340 ;
        RECT 418.240 512.080 418.500 512.340 ;
        RECT 418.240 509.020 418.500 509.280 ;
        RECT 538.300 509.020 538.560 509.280 ;
      LAYER met2 ;
        RECT 412.710 693.755 412.990 694.125 ;
        RECT 412.780 662.650 412.920 693.755 ;
        RECT 414.620 663.950 416.600 664.090 ;
        RECT 414.620 663.330 414.760 663.950 ;
        RECT 414.560 663.010 414.820 663.330 ;
        RECT 412.720 662.330 412.980 662.650 ;
        RECT 416.460 643.010 416.600 663.950 ;
        RECT 416.460 642.870 417.060 643.010 ;
        RECT 416.920 621.930 417.060 642.870 ;
        RECT 416.000 621.790 417.060 621.930 ;
        RECT 416.000 621.250 416.140 621.790 ;
        RECT 414.620 621.170 416.140 621.250 ;
        RECT 414.560 621.110 416.140 621.170 ;
        RECT 414.560 620.850 414.820 621.110 ;
        RECT 414.560 554.890 414.820 555.210 ;
        RECT 414.620 554.610 414.760 554.890 ;
        RECT 414.620 554.470 415.680 554.610 ;
        RECT 415.540 512.370 415.680 554.470 ;
        RECT 415.480 512.050 415.740 512.370 ;
        RECT 418.240 512.050 418.500 512.370 ;
        RECT 418.300 509.310 418.440 512.050 ;
        RECT 418.240 508.990 418.500 509.310 ;
        RECT 538.300 508.990 538.560 509.310 ;
        RECT 538.360 18.770 538.500 508.990 ;
        RECT 538.360 18.630 544.020 18.770 ;
        RECT 543.880 2.400 544.020 18.630 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 412.710 693.800 412.990 694.080 ;
      LAYER met3 ;
        RECT 410.000 696.360 414.000 696.960 ;
        RECT 412.470 694.105 412.770 696.360 ;
        RECT 412.470 693.790 413.015 694.105 ;
        RECT 412.685 693.775 413.015 693.790 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 24.040 562.050 24.100 ;
        RECT 1186.870 24.040 1187.190 24.100 ;
        RECT 561.730 23.900 1187.190 24.040 ;
        RECT 561.730 23.840 562.050 23.900 ;
        RECT 1186.870 23.840 1187.190 23.900 ;
      LAYER via ;
        RECT 561.760 23.840 562.020 24.100 ;
        RECT 1186.900 23.840 1187.160 24.100 ;
      LAYER met2 ;
        RECT 1190.250 510.410 1190.530 514.000 ;
        RECT 1186.960 510.270 1190.530 510.410 ;
        RECT 1186.960 24.130 1187.100 510.270 ;
        RECT 1190.250 510.000 1190.530 510.270 ;
        RECT 561.760 23.810 562.020 24.130 ;
        RECT 1186.900 23.810 1187.160 24.130 ;
        RECT 561.820 2.400 561.960 23.810 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 368.990 539.480 369.310 539.540 ;
        RECT 370.830 539.480 371.150 539.540 ;
        RECT 368.990 539.340 371.150 539.480 ;
        RECT 368.990 539.280 369.310 539.340 ;
        RECT 370.830 539.280 371.150 539.340 ;
      LAYER via ;
        RECT 369.020 539.280 369.280 539.540 ;
        RECT 370.860 539.280 371.120 539.540 ;
      LAYER met2 ;
        RECT 1480.370 3006.690 1480.650 3006.805 ;
        RECT 1481.890 3006.690 1482.170 3010.000 ;
        RECT 1480.370 3006.550 1482.170 3006.690 ;
        RECT 1480.370 3006.435 1480.650 3006.550 ;
        RECT 1481.890 3006.000 1482.170 3006.550 ;
        RECT 370.850 3003.715 371.130 3004.085 ;
        RECT 370.920 539.570 371.060 3003.715 ;
        RECT 369.020 539.250 369.280 539.570 ;
        RECT 370.860 539.250 371.120 539.570 ;
        RECT 369.080 507.805 369.220 539.250 ;
        RECT 369.010 507.435 369.290 507.805 ;
        RECT 580.610 507.435 580.890 507.805 ;
        RECT 580.680 3.130 580.820 507.435 ;
        RECT 579.760 2.990 580.820 3.130 ;
        RECT 579.760 2.400 579.900 2.990 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 1480.370 3006.480 1480.650 3006.760 ;
        RECT 370.850 3003.760 371.130 3004.040 ;
        RECT 369.010 507.480 369.290 507.760 ;
        RECT 580.610 507.480 580.890 507.760 ;
      LAYER met3 ;
        RECT 1480.345 3006.770 1480.675 3006.785 ;
        RECT 1458.510 3006.470 1480.675 3006.770 ;
        RECT 838.390 3006.090 838.770 3006.100 ;
        RECT 861.390 3006.090 861.770 3006.100 ;
        RECT 838.390 3005.790 861.770 3006.090 ;
        RECT 838.390 3005.780 838.770 3005.790 ;
        RECT 861.390 3005.780 861.770 3005.790 ;
        RECT 861.390 3004.420 861.770 3004.740 ;
        RECT 370.825 3004.050 371.155 3004.065 ;
        RECT 838.390 3004.050 838.770 3004.060 ;
        RECT 370.825 3003.750 838.770 3004.050 ;
        RECT 861.430 3004.050 861.730 3004.420 ;
        RECT 1458.510 3004.050 1458.810 3006.470 ;
        RECT 1480.345 3006.455 1480.675 3006.470 ;
        RECT 861.430 3003.750 1458.810 3004.050 ;
        RECT 370.825 3003.735 371.155 3003.750 ;
        RECT 838.390 3003.740 838.770 3003.750 ;
        RECT 368.985 507.770 369.315 507.785 ;
        RECT 580.585 507.770 580.915 507.785 ;
        RECT 368.985 507.470 580.915 507.770 ;
        RECT 368.985 507.455 369.315 507.470 ;
        RECT 580.585 507.455 580.915 507.470 ;
      LAYER via3 ;
        RECT 838.420 3005.780 838.740 3006.100 ;
        RECT 861.420 3005.780 861.740 3006.100 ;
        RECT 861.420 3004.420 861.740 3004.740 ;
        RECT 838.420 3003.740 838.740 3004.060 ;
      LAYER met4 ;
        RECT 838.415 3005.775 838.745 3006.105 ;
        RECT 861.415 3005.775 861.745 3006.105 ;
        RECT 838.430 3004.065 838.730 3005.775 ;
        RECT 861.430 3004.745 861.730 3005.775 ;
        RECT 861.415 3004.415 861.745 3004.745 ;
        RECT 838.415 3003.735 838.745 3004.065 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 51.580 89.630 51.640 ;
        RECT 2187.370 51.580 2187.690 51.640 ;
        RECT 89.310 51.440 2187.690 51.580 ;
        RECT 89.310 51.380 89.630 51.440 ;
        RECT 2187.370 51.380 2187.690 51.440 ;
        RECT 86.090 17.580 86.410 17.640 ;
        RECT 89.310 17.580 89.630 17.640 ;
        RECT 86.090 17.440 89.630 17.580 ;
        RECT 86.090 17.380 86.410 17.440 ;
        RECT 89.310 17.380 89.630 17.440 ;
      LAYER via ;
        RECT 89.340 51.380 89.600 51.640 ;
        RECT 2187.400 51.380 2187.660 51.640 ;
        RECT 86.120 17.380 86.380 17.640 ;
        RECT 89.340 17.380 89.600 17.640 ;
      LAYER met2 ;
        RECT 2191.210 510.410 2191.490 514.000 ;
        RECT 2187.460 510.270 2191.490 510.410 ;
        RECT 2187.460 51.670 2187.600 510.270 ;
        RECT 2191.210 510.000 2191.490 510.270 ;
        RECT 89.340 51.350 89.600 51.670 ;
        RECT 2187.400 51.350 2187.660 51.670 ;
        RECT 89.400 17.670 89.540 51.350 ;
        RECT 86.120 17.350 86.380 17.670 ;
        RECT 89.340 17.350 89.600 17.670 ;
        RECT 86.180 2.400 86.320 17.350 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1449.320 2520.730 1449.380 ;
        RECT 2541.570 1449.320 2541.890 1449.380 ;
        RECT 2520.410 1449.180 2541.890 1449.320 ;
        RECT 2520.410 1449.120 2520.730 1449.180 ;
        RECT 2541.570 1449.120 2541.890 1449.180 ;
        RECT 599.910 334.460 600.230 334.520 ;
        RECT 2541.570 334.460 2541.890 334.520 ;
        RECT 599.910 334.320 2541.890 334.460 ;
        RECT 599.910 334.260 600.230 334.320 ;
        RECT 2541.570 334.260 2541.890 334.320 ;
        RECT 597.150 16.900 597.470 16.960 ;
        RECT 599.910 16.900 600.230 16.960 ;
        RECT 597.150 16.760 600.230 16.900 ;
        RECT 597.150 16.700 597.470 16.760 ;
        RECT 599.910 16.700 600.230 16.760 ;
      LAYER via ;
        RECT 2520.440 1449.120 2520.700 1449.380 ;
        RECT 2541.600 1449.120 2541.860 1449.380 ;
        RECT 599.940 334.260 600.200 334.520 ;
        RECT 2541.600 334.260 2541.860 334.520 ;
        RECT 597.180 16.700 597.440 16.960 ;
        RECT 599.940 16.700 600.200 16.960 ;
      LAYER met2 ;
        RECT 2520.430 1452.635 2520.710 1453.005 ;
        RECT 2520.500 1449.410 2520.640 1452.635 ;
        RECT 2520.440 1449.090 2520.700 1449.410 ;
        RECT 2541.600 1449.090 2541.860 1449.410 ;
        RECT 2541.660 334.550 2541.800 1449.090 ;
        RECT 599.940 334.230 600.200 334.550 ;
        RECT 2541.600 334.230 2541.860 334.550 ;
        RECT 600.000 16.990 600.140 334.230 ;
        RECT 597.180 16.670 597.440 16.990 ;
        RECT 599.940 16.670 600.200 16.990 ;
        RECT 597.240 2.400 597.380 16.670 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1452.680 2520.710 1452.960 ;
      LAYER met3 ;
        RECT 2506.000 1452.970 2510.000 1453.120 ;
        RECT 2520.405 1452.970 2520.735 1452.985 ;
        RECT 2506.000 1452.670 2520.735 1452.970 ;
        RECT 2506.000 1452.520 2510.000 1452.670 ;
        RECT 2520.405 1452.655 2520.735 1452.670 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 413.685 786.845 413.855 793.475 ;
        RECT 413.225 724.285 413.395 741.455 ;
        RECT 414.145 685.865 414.315 701.335 ;
        RECT 434.845 473.365 435.015 474.215 ;
        RECT 482.685 472.685 482.855 474.215 ;
        RECT 579.745 466.225 579.915 473.195 ;
      LAYER mcon ;
        RECT 413.685 793.305 413.855 793.475 ;
        RECT 413.225 741.285 413.395 741.455 ;
        RECT 414.145 701.165 414.315 701.335 ;
        RECT 434.845 474.045 435.015 474.215 ;
        RECT 482.685 474.045 482.855 474.215 ;
        RECT 579.745 473.025 579.915 473.195 ;
      LAYER met1 ;
        RECT 413.625 793.460 413.915 793.505 ;
        RECT 414.070 793.460 414.390 793.520 ;
        RECT 413.625 793.320 414.390 793.460 ;
        RECT 413.625 793.275 413.915 793.320 ;
        RECT 414.070 793.260 414.390 793.320 ;
        RECT 413.610 787.000 413.930 787.060 ;
        RECT 413.415 786.860 413.930 787.000 ;
        RECT 413.610 786.800 413.930 786.860 ;
        RECT 413.165 741.440 413.455 741.485 ;
        RECT 414.530 741.440 414.850 741.500 ;
        RECT 413.165 741.300 414.850 741.440 ;
        RECT 413.165 741.255 413.455 741.300 ;
        RECT 414.530 741.240 414.850 741.300 ;
        RECT 413.165 724.440 413.455 724.485 ;
        RECT 414.070 724.440 414.390 724.500 ;
        RECT 413.165 724.300 414.390 724.440 ;
        RECT 413.165 724.255 413.455 724.300 ;
        RECT 414.070 724.240 414.390 724.300 ;
        RECT 414.070 701.320 414.390 701.380 ;
        RECT 414.070 701.180 414.585 701.320 ;
        RECT 414.070 701.120 414.390 701.180 ;
        RECT 414.070 686.020 414.390 686.080 ;
        RECT 414.070 685.880 414.585 686.020 ;
        RECT 414.070 685.820 414.390 685.880 ;
        RECT 434.785 474.200 435.075 474.245 ;
        RECT 482.625 474.200 482.915 474.245 ;
        RECT 434.785 474.060 482.915 474.200 ;
        RECT 434.785 474.015 435.075 474.060 ;
        RECT 482.625 474.015 482.915 474.060 ;
        RECT 417.290 473.520 417.610 473.580 ;
        RECT 434.785 473.520 435.075 473.565 ;
        RECT 417.290 473.380 435.075 473.520 ;
        RECT 417.290 473.320 417.610 473.380 ;
        RECT 434.785 473.335 435.075 473.380 ;
        RECT 579.685 472.995 579.975 473.225 ;
        RECT 482.625 472.840 482.915 472.885 ;
        RECT 579.760 472.840 579.900 472.995 ;
        RECT 482.625 472.700 579.900 472.840 ;
        RECT 482.625 472.655 482.915 472.700 ;
        RECT 579.685 466.380 579.975 466.425 ;
        RECT 614.170 466.380 614.490 466.440 ;
        RECT 579.685 466.240 614.490 466.380 ;
        RECT 579.685 466.195 579.975 466.240 ;
        RECT 614.170 466.180 614.490 466.240 ;
      LAYER via ;
        RECT 414.100 793.260 414.360 793.520 ;
        RECT 413.640 786.800 413.900 787.060 ;
        RECT 414.560 741.240 414.820 741.500 ;
        RECT 414.100 724.240 414.360 724.500 ;
        RECT 414.100 701.120 414.360 701.380 ;
        RECT 414.100 685.820 414.360 686.080 ;
        RECT 417.320 473.320 417.580 473.580 ;
        RECT 614.200 466.180 614.460 466.440 ;
      LAYER met2 ;
        RECT 413.170 876.930 413.450 877.045 ;
        RECT 413.170 876.790 414.300 876.930 ;
        RECT 413.170 876.675 413.450 876.790 ;
        RECT 414.160 862.650 414.300 876.790 ;
        RECT 414.160 862.510 415.220 862.650 ;
        RECT 415.080 861.970 415.220 862.510 ;
        RECT 414.160 861.830 415.220 861.970 ;
        RECT 414.160 793.550 414.300 861.830 ;
        RECT 414.100 793.230 414.360 793.550 ;
        RECT 413.640 786.770 413.900 787.090 ;
        RECT 413.700 745.690 413.840 786.770 ;
        RECT 413.700 745.550 415.220 745.690 ;
        RECT 415.080 741.610 415.220 745.550 ;
        RECT 414.620 741.530 415.220 741.610 ;
        RECT 414.560 741.470 415.220 741.530 ;
        RECT 414.560 741.210 414.820 741.470 ;
        RECT 414.100 724.210 414.360 724.530 ;
        RECT 414.160 701.410 414.300 724.210 ;
        RECT 414.100 701.090 414.360 701.410 ;
        RECT 414.100 685.790 414.360 686.110 ;
        RECT 414.160 662.730 414.300 685.790 ;
        RECT 414.160 662.590 415.220 662.730 ;
        RECT 415.080 645.730 415.220 662.590 ;
        RECT 414.160 645.590 415.220 645.730 ;
        RECT 414.160 619.890 414.300 645.590 ;
        RECT 414.160 619.750 416.140 619.890 ;
        RECT 416.000 615.130 416.140 619.750 ;
        RECT 415.540 614.990 416.140 615.130 ;
        RECT 415.540 575.690 415.680 614.990 ;
        RECT 415.540 575.550 416.600 575.690 ;
        RECT 416.460 557.330 416.600 575.550 ;
        RECT 416.460 557.190 417.060 557.330 ;
        RECT 416.920 555.290 417.060 557.190 ;
        RECT 416.920 555.150 417.520 555.290 ;
        RECT 417.380 526.730 417.520 555.150 ;
        RECT 416.460 526.590 417.520 526.730 ;
        RECT 416.460 521.970 416.600 526.590 ;
        RECT 416.460 521.830 417.520 521.970 ;
        RECT 417.380 473.610 417.520 521.830 ;
        RECT 417.320 473.290 417.580 473.610 ;
        RECT 614.200 466.150 614.460 466.470 ;
        RECT 614.260 17.410 614.400 466.150 ;
        RECT 614.260 17.270 615.320 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 413.170 876.720 413.450 877.000 ;
      LAYER met3 ;
        RECT 410.000 878.600 414.000 879.200 ;
        RECT 413.390 877.025 413.690 878.600 ;
        RECT 413.145 876.710 413.690 877.025 ;
        RECT 413.145 876.695 413.475 876.710 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 501.060 1204.210 501.120 ;
        RECT 1783.490 501.060 1783.810 501.120 ;
        RECT 1203.890 500.920 1783.810 501.060 ;
        RECT 1203.890 500.860 1204.210 500.920 ;
        RECT 1783.490 500.860 1783.810 500.920 ;
        RECT 110.010 314.400 110.330 314.460 ;
        RECT 1203.890 314.400 1204.210 314.460 ;
        RECT 110.010 314.260 1204.210 314.400 ;
        RECT 110.010 314.200 110.330 314.260 ;
        RECT 1203.890 314.200 1204.210 314.260 ;
      LAYER via ;
        RECT 1203.920 500.860 1204.180 501.120 ;
        RECT 1783.520 500.860 1783.780 501.120 ;
        RECT 110.040 314.200 110.300 314.460 ;
        RECT 1203.920 314.200 1204.180 314.460 ;
      LAYER met2 ;
        RECT 1783.650 510.340 1783.930 514.000 ;
        RECT 1783.580 510.000 1783.930 510.340 ;
        RECT 1783.580 501.150 1783.720 510.000 ;
        RECT 1203.920 500.830 1204.180 501.150 ;
        RECT 1783.520 500.830 1783.780 501.150 ;
        RECT 1203.980 314.490 1204.120 500.830 ;
        RECT 110.040 314.170 110.300 314.490 ;
        RECT 1203.920 314.170 1204.180 314.490 ;
        RECT 110.100 17.410 110.240 314.170 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 3009.920 137.930 3009.980 ;
        RECT 1319.350 3009.920 1319.670 3009.980 ;
        RECT 137.610 3009.780 1319.670 3009.920 ;
        RECT 137.610 3009.720 137.930 3009.780 ;
        RECT 1319.350 3009.720 1319.670 3009.780 ;
        RECT 133.470 17.580 133.790 17.640 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 133.470 17.440 137.930 17.580 ;
        RECT 133.470 17.380 133.790 17.440 ;
        RECT 137.610 17.380 137.930 17.440 ;
      LAYER via ;
        RECT 137.640 3009.720 137.900 3009.980 ;
        RECT 1319.380 3009.720 1319.640 3009.980 ;
        RECT 133.500 17.380 133.760 17.640 ;
        RECT 137.640 17.380 137.900 17.640 ;
      LAYER met2 ;
        RECT 137.640 3009.690 137.900 3010.010 ;
        RECT 1319.380 3009.690 1319.640 3010.010 ;
        RECT 137.700 17.670 137.840 3009.690 ;
        RECT 1319.440 3009.410 1319.580 3009.690 ;
        RECT 1320.890 3009.410 1321.170 3010.000 ;
        RECT 1319.440 3009.270 1321.170 3009.410 ;
        RECT 1320.890 3006.000 1321.170 3009.270 ;
        RECT 133.500 17.350 133.760 17.670 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 133.560 2.400 133.700 17.350 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.590 501.400 1431.910 501.460 ;
        RECT 1573.730 501.400 1574.050 501.460 ;
        RECT 1431.590 501.260 1574.050 501.400 ;
        RECT 1431.590 501.200 1431.910 501.260 ;
        RECT 1573.730 501.200 1574.050 501.260 ;
        RECT 150.950 45.460 151.270 45.520 ;
        RECT 1431.590 45.460 1431.910 45.520 ;
        RECT 150.950 45.320 1431.910 45.460 ;
        RECT 150.950 45.260 151.270 45.320 ;
        RECT 1431.590 45.260 1431.910 45.320 ;
      LAYER via ;
        RECT 1431.620 501.200 1431.880 501.460 ;
        RECT 1573.760 501.200 1574.020 501.460 ;
        RECT 150.980 45.260 151.240 45.520 ;
        RECT 1431.620 45.260 1431.880 45.520 ;
      LAYER met2 ;
        RECT 1573.890 510.340 1574.170 514.000 ;
        RECT 1573.820 510.000 1574.170 510.340 ;
        RECT 1573.820 501.490 1573.960 510.000 ;
        RECT 1431.620 501.170 1431.880 501.490 ;
        RECT 1573.760 501.170 1574.020 501.490 ;
        RECT 1431.680 45.550 1431.820 501.170 ;
        RECT 150.980 45.230 151.240 45.550 ;
        RECT 1431.620 45.230 1431.880 45.550 ;
        RECT 151.040 17.410 151.180 45.230 ;
        RECT 151.040 17.270 151.640 17.410 ;
        RECT 151.500 2.400 151.640 17.270 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 51.920 172.430 51.980 ;
        RECT 1752.670 51.920 1752.990 51.980 ;
        RECT 172.110 51.780 1752.990 51.920 ;
        RECT 172.110 51.720 172.430 51.780 ;
        RECT 1752.670 51.720 1752.990 51.780 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 172.110 17.580 172.430 17.640 ;
        RECT 169.350 17.440 172.430 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 172.110 17.380 172.430 17.440 ;
      LAYER via ;
        RECT 172.140 51.720 172.400 51.980 ;
        RECT 1752.700 51.720 1752.960 51.980 ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 172.140 17.380 172.400 17.640 ;
      LAYER met2 ;
        RECT 1758.810 510.410 1759.090 514.000 ;
        RECT 1752.760 510.270 1759.090 510.410 ;
        RECT 1752.760 52.010 1752.900 510.270 ;
        RECT 1758.810 510.000 1759.090 510.270 ;
        RECT 172.140 51.690 172.400 52.010 ;
        RECT 1752.700 51.690 1752.960 52.010 ;
        RECT 172.200 17.670 172.340 51.690 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 172.140 17.350 172.400 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 134.880 193.130 134.940 ;
        RECT 765.970 134.880 766.290 134.940 ;
        RECT 192.810 134.740 766.290 134.880 ;
        RECT 192.810 134.680 193.130 134.740 ;
        RECT 765.970 134.680 766.290 134.740 ;
        RECT 186.830 17.580 187.150 17.640 ;
        RECT 192.810 17.580 193.130 17.640 ;
        RECT 186.830 17.440 193.130 17.580 ;
        RECT 186.830 17.380 187.150 17.440 ;
        RECT 192.810 17.380 193.130 17.440 ;
      LAYER via ;
        RECT 192.840 134.680 193.100 134.940 ;
        RECT 766.000 134.680 766.260 134.940 ;
        RECT 186.860 17.380 187.120 17.640 ;
        RECT 192.840 17.380 193.100 17.640 ;
      LAYER met2 ;
        RECT 770.730 510.410 771.010 514.000 ;
        RECT 766.060 510.270 771.010 510.410 ;
        RECT 766.060 134.970 766.200 510.270 ;
        RECT 770.730 510.000 771.010 510.270 ;
        RECT 192.840 134.650 193.100 134.970 ;
        RECT 766.000 134.650 766.260 134.970 ;
        RECT 192.900 17.670 193.040 134.650 ;
        RECT 186.860 17.350 187.120 17.670 ;
        RECT 192.840 17.350 193.100 17.670 ;
        RECT 186.920 2.400 187.060 17.350 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 279.290 1166.440 279.610 1166.500 ;
        RECT 393.370 1166.440 393.690 1166.500 ;
        RECT 279.290 1166.300 393.690 1166.440 ;
        RECT 279.290 1166.240 279.610 1166.300 ;
        RECT 393.370 1166.240 393.690 1166.300 ;
        RECT 204.770 24.040 205.090 24.100 ;
        RECT 279.290 24.040 279.610 24.100 ;
        RECT 204.770 23.900 279.610 24.040 ;
        RECT 204.770 23.840 205.090 23.900 ;
        RECT 279.290 23.840 279.610 23.900 ;
      LAYER via ;
        RECT 279.320 1166.240 279.580 1166.500 ;
        RECT 393.400 1166.240 393.660 1166.500 ;
        RECT 204.800 23.840 205.060 24.100 ;
        RECT 279.320 23.840 279.580 24.100 ;
      LAYER met2 ;
        RECT 393.390 1171.115 393.670 1171.485 ;
        RECT 393.460 1166.530 393.600 1171.115 ;
        RECT 279.320 1166.210 279.580 1166.530 ;
        RECT 393.400 1166.210 393.660 1166.530 ;
        RECT 279.380 24.130 279.520 1166.210 ;
        RECT 204.800 23.810 205.060 24.130 ;
        RECT 279.320 23.810 279.580 24.130 ;
        RECT 204.860 2.400 205.000 23.810 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 393.390 1171.160 393.670 1171.440 ;
      LAYER met3 ;
        RECT 393.365 1171.450 393.695 1171.465 ;
        RECT 410.000 1171.450 414.000 1171.600 ;
        RECT 393.365 1171.150 414.000 1171.450 ;
        RECT 393.365 1171.135 393.695 1171.150 ;
        RECT 410.000 1171.000 414.000 1171.150 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1852.950 501.060 1853.270 501.120 ;
        RECT 2042.930 501.060 2043.250 501.120 ;
        RECT 1852.950 500.920 2043.250 501.060 ;
        RECT 1852.950 500.860 1853.270 500.920 ;
        RECT 2042.930 500.860 2043.250 500.920 ;
        RECT 227.310 300.460 227.630 300.520 ;
        RECT 1852.950 300.460 1853.270 300.520 ;
        RECT 227.310 300.320 1853.270 300.460 ;
        RECT 227.310 300.260 227.630 300.320 ;
        RECT 1852.950 300.260 1853.270 300.320 ;
        RECT 222.710 17.580 223.030 17.640 ;
        RECT 227.310 17.580 227.630 17.640 ;
        RECT 222.710 17.440 227.630 17.580 ;
        RECT 222.710 17.380 223.030 17.440 ;
        RECT 227.310 17.380 227.630 17.440 ;
      LAYER via ;
        RECT 1852.980 500.860 1853.240 501.120 ;
        RECT 2042.960 500.860 2043.220 501.120 ;
        RECT 227.340 300.260 227.600 300.520 ;
        RECT 1852.980 300.260 1853.240 300.520 ;
        RECT 222.740 17.380 223.000 17.640 ;
        RECT 227.340 17.380 227.600 17.640 ;
      LAYER met2 ;
        RECT 2043.090 510.340 2043.370 514.000 ;
        RECT 2043.020 510.000 2043.370 510.340 ;
        RECT 2043.020 501.150 2043.160 510.000 ;
        RECT 1852.980 500.830 1853.240 501.150 ;
        RECT 2042.960 500.830 2043.220 501.150 ;
        RECT 1853.040 300.550 1853.180 500.830 ;
        RECT 227.340 300.230 227.600 300.550 ;
        RECT 1852.980 300.230 1853.240 300.550 ;
        RECT 227.400 17.670 227.540 300.230 ;
        RECT 222.740 17.350 223.000 17.670 ;
        RECT 227.340 17.350 227.600 17.670 ;
        RECT 222.800 2.400 222.940 17.350 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 3012.640 45.010 3012.700 ;
        RECT 666.610 3012.640 666.930 3012.700 ;
        RECT 44.690 3012.500 666.930 3012.640 ;
        RECT 44.690 3012.440 45.010 3012.500 ;
        RECT 666.610 3012.440 666.930 3012.500 ;
        RECT 20.310 14.520 20.630 14.580 ;
        RECT 44.690 14.520 45.010 14.580 ;
        RECT 20.310 14.380 45.010 14.520 ;
        RECT 20.310 14.320 20.630 14.380 ;
        RECT 44.690 14.320 45.010 14.380 ;
      LAYER via ;
        RECT 44.720 3012.440 44.980 3012.700 ;
        RECT 666.640 3012.440 666.900 3012.700 ;
        RECT 20.340 14.320 20.600 14.580 ;
        RECT 44.720 14.320 44.980 14.580 ;
      LAYER met2 ;
        RECT 44.720 3012.410 44.980 3012.730 ;
        RECT 666.640 3012.410 666.900 3012.730 ;
        RECT 44.780 14.610 44.920 3012.410 ;
        RECT 666.700 3010.000 666.840 3012.410 ;
        RECT 666.700 3009.340 667.050 3010.000 ;
        RECT 666.770 3006.000 667.050 3009.340 ;
        RECT 20.340 14.290 20.600 14.610 ;
        RECT 44.720 14.290 44.980 14.610 ;
        RECT 20.400 2.400 20.540 14.290 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1038.290 501.400 1038.610 501.460 ;
        RECT 1387.890 501.400 1388.210 501.460 ;
        RECT 1038.290 501.260 1388.210 501.400 ;
        RECT 1038.290 501.200 1038.610 501.260 ;
        RECT 1387.890 501.200 1388.210 501.260 ;
        RECT 47.910 148.820 48.230 148.880 ;
        RECT 1038.290 148.820 1038.610 148.880 ;
        RECT 47.910 148.680 1038.610 148.820 ;
        RECT 47.910 148.620 48.230 148.680 ;
        RECT 1038.290 148.620 1038.610 148.680 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 1038.320 501.200 1038.580 501.460 ;
        RECT 1387.920 501.200 1388.180 501.460 ;
        RECT 47.940 148.620 48.200 148.880 ;
        RECT 1038.320 148.620 1038.580 148.880 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 1388.050 510.340 1388.330 514.000 ;
        RECT 1387.980 510.000 1388.330 510.340 ;
        RECT 1387.980 501.490 1388.120 510.000 ;
        RECT 1038.320 501.170 1038.580 501.490 ;
        RECT 1387.920 501.170 1388.180 501.490 ;
        RECT 1038.380 148.910 1038.520 501.170 ;
        RECT 47.940 148.590 48.200 148.910 ;
        RECT 1038.320 148.590 1038.580 148.910 ;
        RECT 48.000 17.670 48.140 148.590 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1842.700 248.330 1842.760 ;
        RECT 393.370 1842.700 393.690 1842.760 ;
        RECT 248.010 1842.560 393.690 1842.700 ;
        RECT 248.010 1842.500 248.330 1842.560 ;
        RECT 393.370 1842.500 393.690 1842.560 ;
      LAYER via ;
        RECT 248.040 1842.500 248.300 1842.760 ;
        RECT 393.400 1842.500 393.660 1842.760 ;
      LAYER met2 ;
        RECT 393.390 1847.035 393.670 1847.405 ;
        RECT 393.460 1842.790 393.600 1847.035 ;
        RECT 248.040 1842.470 248.300 1842.790 ;
        RECT 393.400 1842.470 393.660 1842.790 ;
        RECT 248.100 17.410 248.240 1842.470 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 393.390 1847.080 393.670 1847.360 ;
      LAYER met3 ;
        RECT 393.365 1847.370 393.695 1847.385 ;
        RECT 410.000 1847.370 414.000 1847.520 ;
        RECT 393.365 1847.070 414.000 1847.370 ;
        RECT 393.365 1847.055 393.695 1847.070 ;
        RECT 410.000 1846.920 414.000 1847.070 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2036.105 3008.065 2036.275 3018.435 ;
      LAYER mcon ;
        RECT 2036.105 3018.265 2036.275 3018.435 ;
      LAYER met1 ;
        RECT 2036.045 3018.420 2036.335 3018.465 ;
        RECT 2346.530 3018.420 2346.850 3018.480 ;
        RECT 2036.045 3018.280 2346.850 3018.420 ;
        RECT 2036.045 3018.235 2036.335 3018.280 ;
        RECT 2346.530 3018.220 2346.850 3018.280 ;
        RECT 461.910 3008.220 462.230 3008.280 ;
        RECT 2036.045 3008.220 2036.335 3008.265 ;
        RECT 461.910 3008.080 2036.335 3008.220 ;
        RECT 461.910 3008.020 462.230 3008.080 ;
        RECT 2036.045 3008.035 2036.335 3008.080 ;
        RECT 264.110 17.580 264.430 17.640 ;
        RECT 268.710 17.580 269.030 17.640 ;
        RECT 264.110 17.440 269.030 17.580 ;
        RECT 264.110 17.380 264.430 17.440 ;
        RECT 268.710 17.380 269.030 17.440 ;
      LAYER via ;
        RECT 2346.560 3018.220 2346.820 3018.480 ;
        RECT 461.940 3008.020 462.200 3008.280 ;
        RECT 264.140 17.380 264.400 17.640 ;
        RECT 268.740 17.380 269.000 17.640 ;
      LAYER met2 ;
        RECT 2346.560 3018.190 2346.820 3018.510 ;
        RECT 2346.620 3010.000 2346.760 3018.190 ;
        RECT 2346.620 3009.340 2346.970 3010.000 ;
        RECT 461.940 3007.990 462.200 3008.310 ;
        RECT 462.000 3006.805 462.140 3007.990 ;
        RECT 416.850 3006.435 417.130 3006.805 ;
        RECT 461.930 3006.435 462.210 3006.805 ;
        RECT 416.920 3002.045 417.060 3006.435 ;
        RECT 2346.690 3006.000 2346.970 3009.340 ;
        RECT 268.730 3001.675 269.010 3002.045 ;
        RECT 416.850 3001.675 417.130 3002.045 ;
        RECT 268.800 17.670 268.940 3001.675 ;
        RECT 264.140 17.350 264.400 17.670 ;
        RECT 268.740 17.350 269.000 17.670 ;
        RECT 264.200 2.400 264.340 17.350 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 416.850 3006.480 417.130 3006.760 ;
        RECT 461.930 3006.480 462.210 3006.760 ;
        RECT 268.730 3001.720 269.010 3002.000 ;
        RECT 416.850 3001.720 417.130 3002.000 ;
      LAYER met3 ;
        RECT 416.825 3006.770 417.155 3006.785 ;
        RECT 461.905 3006.770 462.235 3006.785 ;
        RECT 416.825 3006.470 462.235 3006.770 ;
        RECT 416.825 3006.455 417.155 3006.470 ;
        RECT 461.905 3006.455 462.235 3006.470 ;
        RECT 268.705 3002.010 269.035 3002.025 ;
        RECT 416.825 3002.010 417.155 3002.025 ;
        RECT 268.705 3001.710 417.155 3002.010 ;
        RECT 268.705 3001.695 269.035 3001.710 ;
        RECT 416.825 3001.695 417.155 3001.710 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 655.760 286.510 655.820 ;
        RECT 393.370 655.760 393.690 655.820 ;
        RECT 286.190 655.620 393.690 655.760 ;
        RECT 286.190 655.560 286.510 655.620 ;
        RECT 393.370 655.560 393.690 655.620 ;
        RECT 282.510 76.060 282.830 76.120 ;
        RECT 286.190 76.060 286.510 76.120 ;
        RECT 282.510 75.920 286.510 76.060 ;
        RECT 282.510 75.860 282.830 75.920 ;
        RECT 286.190 75.860 286.510 75.920 ;
      LAYER via ;
        RECT 286.220 655.560 286.480 655.820 ;
        RECT 393.400 655.560 393.660 655.820 ;
        RECT 282.540 75.860 282.800 76.120 ;
        RECT 286.220 75.860 286.480 76.120 ;
      LAYER met2 ;
        RECT 393.390 659.755 393.670 660.125 ;
        RECT 393.460 655.850 393.600 659.755 ;
        RECT 286.220 655.530 286.480 655.850 ;
        RECT 393.400 655.530 393.660 655.850 ;
        RECT 286.280 76.150 286.420 655.530 ;
        RECT 282.540 75.830 282.800 76.150 ;
        RECT 286.220 75.830 286.480 76.150 ;
        RECT 282.600 3.130 282.740 75.830 ;
        RECT 282.140 2.990 282.740 3.130 ;
        RECT 282.140 2.400 282.280 2.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 393.390 659.800 393.670 660.080 ;
      LAYER met3 ;
        RECT 393.365 660.090 393.695 660.105 ;
        RECT 410.000 660.090 414.000 660.240 ;
        RECT 393.365 659.790 414.000 660.090 ;
        RECT 393.365 659.775 393.695 659.790 ;
        RECT 410.000 659.640 414.000 659.790 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 3017.400 1759.430 3017.460 ;
        RECT 2334.570 3017.400 2334.890 3017.460 ;
        RECT 1759.110 3017.260 2334.890 3017.400 ;
        RECT 1759.110 3017.200 1759.430 3017.260 ;
        RECT 2334.570 3017.200 2334.890 3017.260 ;
        RECT 441.670 3015.360 441.990 3015.420 ;
        RECT 1759.110 3015.360 1759.430 3015.420 ;
        RECT 441.670 3015.220 1759.430 3015.360 ;
        RECT 441.670 3015.160 441.990 3015.220 ;
        RECT 1759.110 3015.160 1759.430 3015.220 ;
        RECT 299.990 17.580 300.310 17.640 ;
        RECT 303.210 17.580 303.530 17.640 ;
        RECT 299.990 17.440 303.530 17.580 ;
        RECT 299.990 17.380 300.310 17.440 ;
        RECT 303.210 17.380 303.530 17.440 ;
      LAYER via ;
        RECT 1759.140 3017.200 1759.400 3017.460 ;
        RECT 2334.600 3017.200 2334.860 3017.460 ;
        RECT 441.700 3015.160 441.960 3015.420 ;
        RECT 1759.140 3015.160 1759.400 3015.420 ;
        RECT 300.020 17.380 300.280 17.640 ;
        RECT 303.240 17.380 303.500 17.640 ;
      LAYER met2 ;
        RECT 1759.140 3017.170 1759.400 3017.490 ;
        RECT 2334.600 3017.170 2334.860 3017.490 ;
        RECT 1759.200 3015.450 1759.340 3017.170 ;
        RECT 441.700 3015.130 441.960 3015.450 ;
        RECT 1759.140 3015.130 1759.400 3015.450 ;
        RECT 441.760 3011.565 441.900 3015.130 ;
        RECT 303.230 3011.195 303.510 3011.565 ;
        RECT 441.690 3011.195 441.970 3011.565 ;
        RECT 303.300 17.670 303.440 3011.195 ;
        RECT 2334.660 3010.000 2334.800 3017.170 ;
        RECT 2334.660 3009.340 2335.010 3010.000 ;
        RECT 2334.730 3006.000 2335.010 3009.340 ;
        RECT 300.020 17.350 300.280 17.670 ;
        RECT 303.240 17.350 303.500 17.670 ;
        RECT 300.080 2.400 300.220 17.350 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 303.230 3011.240 303.510 3011.520 ;
        RECT 441.690 3011.240 441.970 3011.520 ;
      LAYER met3 ;
        RECT 303.205 3011.530 303.535 3011.545 ;
        RECT 441.665 3011.530 441.995 3011.545 ;
        RECT 303.205 3011.230 441.995 3011.530 ;
        RECT 303.205 3011.215 303.535 3011.230 ;
        RECT 441.665 3011.215 441.995 3011.230 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2507.530 2780.560 2507.850 2780.820 ;
        RECT 2507.620 2780.140 2507.760 2780.560 ;
        RECT 2507.530 2779.880 2507.850 2780.140 ;
        RECT 317.930 17.580 318.250 17.640 ;
        RECT 321.150 17.580 321.470 17.640 ;
        RECT 317.930 17.440 321.470 17.580 ;
        RECT 317.930 17.380 318.250 17.440 ;
        RECT 321.150 17.380 321.470 17.440 ;
      LAYER via ;
        RECT 2507.560 2780.560 2507.820 2780.820 ;
        RECT 2507.560 2779.880 2507.820 2780.140 ;
        RECT 317.960 17.380 318.220 17.640 ;
        RECT 321.180 17.380 321.440 17.640 ;
      LAYER met2 ;
        RECT 2507.550 2947.275 2507.830 2947.645 ;
        RECT 2507.620 2780.850 2507.760 2947.275 ;
        RECT 2507.560 2780.530 2507.820 2780.850 ;
        RECT 2507.560 2779.850 2507.820 2780.170 ;
        RECT 2507.620 689.365 2507.760 2779.850 ;
        RECT 2507.550 688.995 2507.830 689.365 ;
        RECT 2500.190 227.275 2500.470 227.645 ;
        RECT 2500.260 196.365 2500.400 227.275 ;
        RECT 321.170 195.995 321.450 196.365 ;
        RECT 2500.190 195.995 2500.470 196.365 ;
        RECT 321.240 17.670 321.380 195.995 ;
        RECT 317.960 17.350 318.220 17.670 ;
        RECT 321.180 17.350 321.440 17.670 ;
        RECT 318.020 2.400 318.160 17.350 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 2507.550 2947.320 2507.830 2947.600 ;
        RECT 2507.550 689.040 2507.830 689.320 ;
        RECT 2500.190 227.320 2500.470 227.600 ;
        RECT 321.170 196.040 321.450 196.320 ;
        RECT 2500.190 196.040 2500.470 196.320 ;
      LAYER met3 ;
        RECT 2506.000 2949.880 2510.000 2950.480 ;
        RECT 2507.310 2947.625 2507.610 2949.880 ;
        RECT 2507.310 2947.310 2507.855 2947.625 ;
        RECT 2507.525 2947.295 2507.855 2947.310 ;
        RECT 2507.525 689.330 2507.855 689.345 ;
        RECT 2508.190 689.330 2508.570 689.340 ;
        RECT 2507.525 689.030 2508.570 689.330 ;
        RECT 2507.525 689.015 2507.855 689.030 ;
        RECT 2508.190 689.020 2508.570 689.030 ;
        RECT 2504.510 513.210 2504.890 513.220 ;
        RECT 2506.350 513.210 2506.730 513.220 ;
        RECT 2504.510 512.910 2506.730 513.210 ;
        RECT 2504.510 512.900 2504.890 512.910 ;
        RECT 2506.350 512.900 2506.730 512.910 ;
        RECT 2506.350 462.210 2506.730 462.220 ;
        RECT 2505.470 461.910 2506.730 462.210 ;
        RECT 2505.470 461.540 2505.770 461.910 ;
        RECT 2506.350 461.900 2506.730 461.910 ;
        RECT 2505.430 461.220 2505.810 461.540 ;
        RECT 2504.510 304.140 2504.890 304.460 ;
        RECT 2504.550 303.090 2504.850 304.140 ;
        RECT 2505.430 303.090 2505.810 303.100 ;
        RECT 2504.550 302.790 2505.810 303.090 ;
        RECT 2505.430 302.780 2505.810 302.790 ;
        RECT 2500.165 227.610 2500.495 227.625 ;
        RECT 2505.430 227.610 2505.810 227.620 ;
        RECT 2500.165 227.310 2505.810 227.610 ;
        RECT 2500.165 227.295 2500.495 227.310 ;
        RECT 2505.430 227.300 2505.810 227.310 ;
        RECT 321.145 196.330 321.475 196.345 ;
        RECT 2500.165 196.330 2500.495 196.345 ;
        RECT 321.145 196.030 2500.495 196.330 ;
        RECT 321.145 196.015 321.475 196.030 ;
        RECT 2500.165 196.015 2500.495 196.030 ;
      LAYER via3 ;
        RECT 2508.220 689.020 2508.540 689.340 ;
        RECT 2504.540 512.900 2504.860 513.220 ;
        RECT 2506.380 512.900 2506.700 513.220 ;
        RECT 2506.380 461.900 2506.700 462.220 ;
        RECT 2505.460 461.220 2505.780 461.540 ;
        RECT 2504.540 304.140 2504.860 304.460 ;
        RECT 2505.460 302.780 2505.780 303.100 ;
        RECT 2505.460 227.300 2505.780 227.620 ;
      LAYER met4 ;
        RECT 2508.215 689.015 2508.545 689.345 ;
        RECT 2508.230 607.050 2508.530 689.015 ;
        RECT 2505.470 606.750 2508.530 607.050 ;
        RECT 2505.470 603.650 2505.770 606.750 ;
        RECT 2504.550 603.350 2505.770 603.650 ;
        RECT 2504.550 513.225 2504.850 603.350 ;
        RECT 2504.535 512.895 2504.865 513.225 ;
        RECT 2506.375 512.895 2506.705 513.225 ;
        RECT 2506.390 462.225 2506.690 512.895 ;
        RECT 2506.375 461.895 2506.705 462.225 ;
        RECT 2505.455 461.215 2505.785 461.545 ;
        RECT 2505.470 335.050 2505.770 461.215 ;
        RECT 2504.550 334.750 2505.770 335.050 ;
        RECT 2504.550 304.465 2504.850 334.750 ;
        RECT 2504.535 304.135 2504.865 304.465 ;
        RECT 2505.455 302.775 2505.785 303.105 ;
        RECT 2505.470 227.625 2505.770 302.775 ;
        RECT 2505.455 227.295 2505.785 227.625 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 950.430 3018.760 950.750 3018.820 ;
        RECT 2087.090 3018.760 2087.410 3018.820 ;
        RECT 950.430 3018.620 2087.410 3018.760 ;
        RECT 950.430 3018.560 950.750 3018.620 ;
        RECT 2087.090 3018.560 2087.410 3018.620 ;
      LAYER via ;
        RECT 950.460 3018.560 950.720 3018.820 ;
        RECT 2087.120 3018.560 2087.380 3018.820 ;
      LAYER met2 ;
        RECT 950.450 3024.115 950.730 3024.485 ;
        RECT 950.520 3018.850 950.660 3024.115 ;
        RECT 950.460 3018.530 950.720 3018.850 ;
        RECT 2087.120 3018.530 2087.380 3018.850 ;
        RECT 2087.180 3010.000 2087.320 3018.530 ;
        RECT 2087.180 3009.340 2087.530 3010.000 ;
        RECT 2087.250 3006.000 2087.530 3009.340 ;
        RECT 334.970 2172.755 335.250 2173.125 ;
        RECT 335.040 2149.325 335.180 2172.755 ;
        RECT 334.970 2148.955 335.250 2149.325 ;
        RECT 334.510 1641.675 334.790 1642.045 ;
        RECT 334.580 1618.245 334.720 1641.675 ;
        RECT 334.510 1617.875 334.790 1618.245 ;
        RECT 335.430 1029.675 335.710 1030.045 ;
        RECT 335.500 1027.325 335.640 1029.675 ;
        RECT 335.430 1026.955 335.710 1027.325 ;
        RECT 335.890 17.155 336.170 17.525 ;
        RECT 335.960 2.400 336.100 17.155 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 950.450 3024.160 950.730 3024.440 ;
        RECT 334.970 2172.800 335.250 2173.080 ;
        RECT 334.970 2149.000 335.250 2149.280 ;
        RECT 334.510 1641.720 334.790 1642.000 ;
        RECT 334.510 1617.920 334.790 1618.200 ;
        RECT 335.430 1029.720 335.710 1030.000 ;
        RECT 335.430 1027.000 335.710 1027.280 ;
        RECT 335.890 17.200 336.170 17.480 ;
      LAYER met3 ;
        RECT 336.990 3024.450 337.370 3024.460 ;
        RECT 950.425 3024.450 950.755 3024.465 ;
        RECT 336.990 3024.150 950.755 3024.450 ;
        RECT 336.990 3024.140 337.370 3024.150 ;
        RECT 950.425 3024.135 950.755 3024.150 ;
        RECT 334.945 2173.090 335.275 2173.105 ;
        RECT 336.990 2173.090 337.370 2173.100 ;
        RECT 334.945 2172.790 337.370 2173.090 ;
        RECT 334.945 2172.775 335.275 2172.790 ;
        RECT 336.990 2172.780 337.370 2172.790 ;
        RECT 334.945 2149.290 335.275 2149.305 ;
        RECT 336.990 2149.290 337.370 2149.300 ;
        RECT 334.945 2148.990 337.370 2149.290 ;
        RECT 334.945 2148.975 335.275 2148.990 ;
        RECT 336.990 2148.980 337.370 2148.990 ;
        RECT 334.485 1642.010 334.815 1642.025 ;
        RECT 336.990 1642.010 337.370 1642.020 ;
        RECT 334.485 1641.710 337.370 1642.010 ;
        RECT 334.485 1641.695 334.815 1641.710 ;
        RECT 336.990 1641.700 337.370 1641.710 ;
        RECT 334.485 1618.210 334.815 1618.225 ;
        RECT 336.990 1618.210 337.370 1618.220 ;
        RECT 334.485 1617.910 337.370 1618.210 ;
        RECT 334.485 1617.895 334.815 1617.910 ;
        RECT 336.990 1617.900 337.370 1617.910 ;
        RECT 336.990 1210.210 337.370 1210.220 ;
        RECT 336.110 1209.910 337.370 1210.210 ;
        RECT 336.110 1208.170 336.410 1209.910 ;
        RECT 336.990 1209.900 337.370 1209.910 ;
        RECT 336.990 1208.170 337.370 1208.180 ;
        RECT 336.110 1207.870 337.370 1208.170 ;
        RECT 336.990 1207.860 337.370 1207.870 ;
        RECT 335.405 1030.010 335.735 1030.025 ;
        RECT 336.990 1030.010 337.370 1030.020 ;
        RECT 335.405 1029.710 337.370 1030.010 ;
        RECT 335.405 1029.695 335.735 1029.710 ;
        RECT 336.990 1029.700 337.370 1029.710 ;
        RECT 335.405 1027.290 335.735 1027.305 ;
        RECT 336.990 1027.290 337.370 1027.300 ;
        RECT 335.405 1026.990 337.370 1027.290 ;
        RECT 335.405 1026.975 335.735 1026.990 ;
        RECT 336.990 1026.980 337.370 1026.990 ;
        RECT 335.865 17.490 336.195 17.505 ;
        RECT 336.990 17.490 337.370 17.500 ;
        RECT 335.865 17.190 337.370 17.490 ;
        RECT 335.865 17.175 336.195 17.190 ;
        RECT 336.990 17.180 337.370 17.190 ;
      LAYER via3 ;
        RECT 337.020 3024.140 337.340 3024.460 ;
        RECT 337.020 2172.780 337.340 2173.100 ;
        RECT 337.020 2148.980 337.340 2149.300 ;
        RECT 337.020 1641.700 337.340 1642.020 ;
        RECT 337.020 1617.900 337.340 1618.220 ;
        RECT 337.020 1209.900 337.340 1210.220 ;
        RECT 337.020 1207.860 337.340 1208.180 ;
        RECT 337.020 1029.700 337.340 1030.020 ;
        RECT 337.020 1026.980 337.340 1027.300 ;
        RECT 337.020 17.180 337.340 17.500 ;
      LAYER met4 ;
        RECT 337.015 3024.135 337.345 3024.465 ;
        RECT 337.030 2173.105 337.330 3024.135 ;
        RECT 337.015 2172.775 337.345 2173.105 ;
        RECT 337.015 2148.975 337.345 2149.305 ;
        RECT 337.030 1642.025 337.330 2148.975 ;
        RECT 337.015 1641.695 337.345 1642.025 ;
        RECT 337.015 1617.895 337.345 1618.225 ;
        RECT 337.030 1210.225 337.330 1617.895 ;
        RECT 337.015 1209.895 337.345 1210.225 ;
        RECT 337.015 1207.855 337.345 1208.185 ;
        RECT 337.030 1030.025 337.330 1207.855 ;
        RECT 337.015 1029.695 337.345 1030.025 ;
        RECT 337.015 1026.975 337.345 1027.305 ;
        RECT 337.030 17.505 337.330 1026.975 ;
        RECT 337.015 17.175 337.345 17.505 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1127.990 500.380 1128.310 500.440 ;
        RECT 1202.970 500.380 1203.290 500.440 ;
        RECT 1127.990 500.240 1203.290 500.380 ;
        RECT 1127.990 500.180 1128.310 500.240 ;
        RECT 1202.970 500.180 1203.290 500.240 ;
        RECT 353.350 32.880 353.670 32.940 ;
        RECT 1127.990 32.880 1128.310 32.940 ;
        RECT 353.350 32.740 1128.310 32.880 ;
        RECT 353.350 32.680 353.670 32.740 ;
        RECT 1127.990 32.680 1128.310 32.740 ;
      LAYER via ;
        RECT 1128.020 500.180 1128.280 500.440 ;
        RECT 1203.000 500.180 1203.260 500.440 ;
        RECT 353.380 32.680 353.640 32.940 ;
        RECT 1128.020 32.680 1128.280 32.940 ;
      LAYER met2 ;
        RECT 1203.130 510.340 1203.410 514.000 ;
        RECT 1203.060 510.000 1203.410 510.340 ;
        RECT 1203.060 500.470 1203.200 510.000 ;
        RECT 1128.020 500.150 1128.280 500.470 ;
        RECT 1203.000 500.150 1203.260 500.470 ;
        RECT 1128.080 32.970 1128.220 500.150 ;
        RECT 353.380 32.650 353.640 32.970 ;
        RECT 1128.020 32.650 1128.280 32.970 ;
        RECT 353.440 2.400 353.580 32.650 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 615.625 3004.325 615.795 3006.535 ;
      LAYER mcon ;
        RECT 615.625 3006.365 615.795 3006.535 ;
      LAYER met1 ;
        RECT 615.550 3006.520 615.870 3006.580 ;
        RECT 615.355 3006.380 615.870 3006.520 ;
        RECT 615.550 3006.320 615.870 3006.380 ;
        RECT 371.750 3004.480 372.070 3004.540 ;
        RECT 615.565 3004.480 615.855 3004.525 ;
        RECT 371.750 3004.340 615.855 3004.480 ;
        RECT 371.750 3004.280 372.070 3004.340 ;
        RECT 615.565 3004.295 615.855 3004.340 ;
      LAYER via ;
        RECT 615.580 3006.320 615.840 3006.580 ;
        RECT 371.780 3004.280 372.040 3004.540 ;
      LAYER met2 ;
        RECT 617.090 3006.690 617.370 3010.000 ;
        RECT 615.640 3006.610 617.370 3006.690 ;
        RECT 615.580 3006.550 617.370 3006.610 ;
        RECT 615.580 3006.290 615.840 3006.550 ;
        RECT 617.090 3006.000 617.370 3006.550 ;
        RECT 371.780 3004.250 372.040 3004.570 ;
        RECT 371.840 3.130 371.980 3004.250 ;
        RECT 371.380 2.990 371.980 3.130 ;
        RECT 371.380 2.400 371.520 2.990 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 391.530 1227.980 391.850 1228.040 ;
        RECT 397.510 1227.980 397.830 1228.040 ;
        RECT 391.530 1227.840 397.830 1227.980 ;
        RECT 391.530 1227.780 391.850 1227.840 ;
        RECT 397.510 1227.780 397.830 1227.840 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 391.530 16.900 391.850 16.960 ;
        RECT 389.230 16.760 391.850 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 391.530 16.700 391.850 16.760 ;
      LAYER via ;
        RECT 391.560 1227.780 391.820 1228.040 ;
        RECT 397.540 1227.780 397.800 1228.040 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 391.560 16.700 391.820 16.960 ;
      LAYER met2 ;
        RECT 397.530 2467.195 397.810 2467.565 ;
        RECT 397.600 1228.070 397.740 2467.195 ;
        RECT 391.560 1227.750 391.820 1228.070 ;
        RECT 397.540 1227.750 397.800 1228.070 ;
        RECT 391.620 16.990 391.760 1227.750 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 391.560 16.670 391.820 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 397.530 2467.240 397.810 2467.520 ;
      LAYER met3 ;
        RECT 397.505 2467.530 397.835 2467.545 ;
        RECT 410.000 2467.530 414.000 2467.680 ;
        RECT 397.505 2467.230 414.000 2467.530 ;
        RECT 397.505 2467.215 397.835 2467.230 ;
        RECT 410.000 2467.080 414.000 2467.230 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 289.410 3043.240 289.730 3043.300 ;
        RECT 1568.210 3043.240 1568.530 3043.300 ;
        RECT 289.410 3043.100 1568.530 3043.240 ;
        RECT 289.410 3043.040 289.730 3043.100 ;
        RECT 1568.210 3043.040 1568.530 3043.100 ;
        RECT 289.410 486.780 289.730 486.840 ;
        RECT 407.170 486.780 407.490 486.840 ;
        RECT 289.410 486.640 407.490 486.780 ;
        RECT 289.410 486.580 289.730 486.640 ;
        RECT 407.170 486.580 407.490 486.640 ;
      LAYER via ;
        RECT 289.440 3043.040 289.700 3043.300 ;
        RECT 1568.240 3043.040 1568.500 3043.300 ;
        RECT 289.440 486.580 289.700 486.840 ;
        RECT 407.200 486.580 407.460 486.840 ;
      LAYER met2 ;
        RECT 289.440 3043.010 289.700 3043.330 ;
        RECT 1568.240 3043.010 1568.500 3043.330 ;
        RECT 289.500 486.870 289.640 3043.010 ;
        RECT 1568.300 3010.000 1568.440 3043.010 ;
        RECT 1568.300 3009.340 1568.650 3010.000 ;
        RECT 1568.370 3006.000 1568.650 3009.340 ;
        RECT 289.440 486.550 289.700 486.870 ;
        RECT 407.200 486.550 407.460 486.870 ;
        RECT 407.260 2.400 407.400 486.550 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 154.515 68.450 154.885 ;
        RECT 68.240 2.400 68.380 154.515 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 68.170 154.560 68.450 154.840 ;
      LAYER met3 ;
        RECT 2506.000 2092.170 2510.000 2092.320 ;
        RECT 2546.830 2092.170 2547.210 2092.180 ;
        RECT 2506.000 2091.870 2547.210 2092.170 ;
        RECT 2506.000 2091.720 2510.000 2091.870 ;
        RECT 2546.830 2091.860 2547.210 2091.870 ;
        RECT 68.145 154.850 68.475 154.865 ;
        RECT 2546.830 154.850 2547.210 154.860 ;
        RECT 68.145 154.550 2547.210 154.850 ;
        RECT 68.145 154.535 68.475 154.550 ;
        RECT 2546.830 154.540 2547.210 154.550 ;
      LAYER via3 ;
        RECT 2546.860 2091.860 2547.180 2092.180 ;
        RECT 2546.860 154.540 2547.180 154.860 ;
      LAYER met4 ;
        RECT 2546.855 2091.855 2547.185 2092.185 ;
        RECT 2546.870 154.865 2547.170 2091.855 ;
        RECT 2546.855 154.535 2547.185 154.865 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 2125.580 2519.810 2125.640 ;
        RECT 2547.090 2125.580 2547.410 2125.640 ;
        RECT 2519.490 2125.440 2547.410 2125.580 ;
        RECT 2519.490 2125.380 2519.810 2125.440 ;
        RECT 2547.090 2125.380 2547.410 2125.440 ;
        RECT 427.410 93.060 427.730 93.120 ;
        RECT 2547.090 93.060 2547.410 93.120 ;
        RECT 427.410 92.920 2547.410 93.060 ;
        RECT 427.410 92.860 427.730 92.920 ;
        RECT 2547.090 92.860 2547.410 92.920 ;
        RECT 424.650 15.200 424.970 15.260 ;
        RECT 427.410 15.200 427.730 15.260 ;
        RECT 424.650 15.060 427.730 15.200 ;
        RECT 424.650 15.000 424.970 15.060 ;
        RECT 427.410 15.000 427.730 15.060 ;
      LAYER via ;
        RECT 2519.520 2125.380 2519.780 2125.640 ;
        RECT 2547.120 2125.380 2547.380 2125.640 ;
        RECT 427.440 92.860 427.700 93.120 ;
        RECT 2547.120 92.860 2547.380 93.120 ;
        RECT 424.680 15.000 424.940 15.260 ;
        RECT 427.440 15.000 427.700 15.260 ;
      LAYER met2 ;
        RECT 2519.510 2128.555 2519.790 2128.925 ;
        RECT 2519.580 2125.670 2519.720 2128.555 ;
        RECT 2519.520 2125.350 2519.780 2125.670 ;
        RECT 2547.120 2125.350 2547.380 2125.670 ;
        RECT 2547.180 93.150 2547.320 2125.350 ;
        RECT 427.440 92.830 427.700 93.150 ;
        RECT 2547.120 92.830 2547.380 93.150 ;
        RECT 427.500 15.290 427.640 92.830 ;
        RECT 424.680 14.970 424.940 15.290 ;
        RECT 427.440 14.970 427.700 15.290 ;
        RECT 424.740 2.400 424.880 14.970 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 2519.510 2128.600 2519.790 2128.880 ;
      LAYER met3 ;
        RECT 2506.000 2128.890 2510.000 2129.040 ;
        RECT 2519.485 2128.890 2519.815 2128.905 ;
        RECT 2506.000 2128.590 2519.815 2128.890 ;
        RECT 2506.000 2128.440 2510.000 2128.590 ;
        RECT 2519.485 2128.575 2519.815 2128.590 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 3017.740 282.830 3017.800 ;
        RECT 555.290 3017.740 555.610 3017.800 ;
        RECT 282.510 3017.600 555.610 3017.740 ;
        RECT 282.510 3017.540 282.830 3017.600 ;
        RECT 555.290 3017.540 555.610 3017.600 ;
        RECT 282.510 508.540 282.830 508.600 ;
        RECT 442.590 508.540 442.910 508.600 ;
        RECT 282.510 508.400 442.910 508.540 ;
        RECT 282.510 508.340 282.830 508.400 ;
        RECT 442.590 508.340 442.910 508.400 ;
      LAYER via ;
        RECT 282.540 3017.540 282.800 3017.800 ;
        RECT 555.320 3017.540 555.580 3017.800 ;
        RECT 282.540 508.340 282.800 508.600 ;
        RECT 442.620 508.340 442.880 508.600 ;
      LAYER met2 ;
        RECT 282.540 3017.510 282.800 3017.830 ;
        RECT 555.320 3017.510 555.580 3017.830 ;
        RECT 282.600 508.630 282.740 3017.510 ;
        RECT 555.380 3010.000 555.520 3017.510 ;
        RECT 555.380 3009.340 555.730 3010.000 ;
        RECT 555.450 3006.000 555.730 3009.340 ;
        RECT 282.540 508.310 282.800 508.630 ;
        RECT 442.620 508.310 442.880 508.630 ;
        RECT 442.680 503.610 442.820 508.310 ;
        RECT 441.760 503.470 442.820 503.610 ;
        RECT 441.760 16.900 441.900 503.470 ;
        RECT 441.760 16.760 442.820 16.900 ;
        RECT 442.680 2.400 442.820 16.760 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 934.790 500.720 935.110 500.780 ;
        RECT 1066.810 500.720 1067.130 500.780 ;
        RECT 934.790 500.580 1067.130 500.720 ;
        RECT 934.790 500.520 935.110 500.580 ;
        RECT 1066.810 500.520 1067.130 500.580 ;
        RECT 461.910 74.700 462.230 74.760 ;
        RECT 934.790 74.700 935.110 74.760 ;
        RECT 461.910 74.560 935.110 74.700 ;
        RECT 461.910 74.500 462.230 74.560 ;
        RECT 934.790 74.500 935.110 74.560 ;
      LAYER via ;
        RECT 934.820 500.520 935.080 500.780 ;
        RECT 1066.840 500.520 1067.100 500.780 ;
        RECT 461.940 74.500 462.200 74.760 ;
        RECT 934.820 74.500 935.080 74.760 ;
      LAYER met2 ;
        RECT 1066.970 510.340 1067.250 514.000 ;
        RECT 1066.900 510.000 1067.250 510.340 ;
        RECT 1066.900 500.810 1067.040 510.000 ;
        RECT 934.820 500.490 935.080 500.810 ;
        RECT 1066.840 500.490 1067.100 500.810 ;
        RECT 934.880 74.790 935.020 500.490 ;
        RECT 461.940 74.470 462.200 74.790 ;
        RECT 934.820 74.470 935.080 74.790 ;
        RECT 462.000 16.900 462.140 74.470 ;
        RECT 460.620 16.760 462.140 16.900 ;
        RECT 460.620 2.400 460.760 16.760 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 341.600 482.930 341.660 ;
        RECT 2520.870 341.600 2521.190 341.660 ;
        RECT 482.610 341.460 2521.190 341.600 ;
        RECT 482.610 341.400 482.930 341.460 ;
        RECT 2520.870 341.400 2521.190 341.460 ;
        RECT 478.470 16.900 478.790 16.960 ;
        RECT 482.610 16.900 482.930 16.960 ;
        RECT 478.470 16.760 482.930 16.900 ;
        RECT 478.470 16.700 478.790 16.760 ;
        RECT 482.610 16.700 482.930 16.760 ;
      LAYER via ;
        RECT 482.640 341.400 482.900 341.660 ;
        RECT 2520.900 341.400 2521.160 341.660 ;
        RECT 478.500 16.700 478.760 16.960 ;
        RECT 482.640 16.700 482.900 16.960 ;
      LAYER met2 ;
        RECT 2520.890 867.835 2521.170 868.205 ;
        RECT 2520.960 341.690 2521.100 867.835 ;
        RECT 482.640 341.370 482.900 341.690 ;
        RECT 2520.900 341.370 2521.160 341.690 ;
        RECT 482.700 16.990 482.840 341.370 ;
        RECT 478.500 16.670 478.760 16.990 ;
        RECT 482.640 16.670 482.900 16.990 ;
        RECT 478.560 2.400 478.700 16.670 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 2520.890 867.880 2521.170 868.160 ;
      LAYER met3 ;
        RECT 2506.000 868.170 2510.000 868.320 ;
        RECT 2520.865 868.170 2521.195 868.185 ;
        RECT 2506.000 867.870 2521.195 868.170 ;
        RECT 2506.000 867.720 2510.000 867.870 ;
        RECT 2520.865 867.855 2521.195 867.870 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.970 134.115 496.250 134.485 ;
        RECT 496.040 17.410 496.180 134.115 ;
        RECT 496.040 17.270 496.640 17.410 ;
        RECT 496.500 2.400 496.640 17.270 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 495.970 134.160 496.250 134.440 ;
      LAYER met3 ;
        RECT 2506.000 960.650 2510.000 960.800 ;
        RECT 2520.150 960.650 2520.530 960.660 ;
        RECT 2506.000 960.350 2520.530 960.650 ;
        RECT 2506.000 960.200 2510.000 960.350 ;
        RECT 2520.150 960.340 2520.530 960.350 ;
        RECT 495.945 134.450 496.275 134.465 ;
        RECT 2520.150 134.450 2520.530 134.460 ;
        RECT 495.945 134.150 2520.530 134.450 ;
        RECT 495.945 134.135 496.275 134.150 ;
        RECT 2520.150 134.140 2520.530 134.150 ;
      LAYER via3 ;
        RECT 2520.180 960.340 2520.500 960.660 ;
        RECT 2520.180 134.140 2520.500 134.460 ;
      LAYER met4 ;
        RECT 2520.175 960.335 2520.505 960.665 ;
        RECT 2520.190 134.465 2520.490 960.335 ;
        RECT 2520.175 134.135 2520.505 134.465 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 142.020 517.430 142.080 ;
        RECT 2104.570 142.020 2104.890 142.080 ;
        RECT 517.110 141.880 2104.890 142.020 ;
        RECT 517.110 141.820 517.430 141.880 ;
        RECT 2104.570 141.820 2104.890 141.880 ;
        RECT 513.890 16.900 514.210 16.960 ;
        RECT 517.110 16.900 517.430 16.960 ;
        RECT 513.890 16.760 517.430 16.900 ;
        RECT 513.890 16.700 514.210 16.760 ;
        RECT 517.110 16.700 517.430 16.760 ;
      LAYER via ;
        RECT 517.140 141.820 517.400 142.080 ;
        RECT 2104.600 141.820 2104.860 142.080 ;
        RECT 513.920 16.700 514.180 16.960 ;
        RECT 517.140 16.700 517.400 16.960 ;
      LAYER met2 ;
        RECT 2104.730 510.340 2105.010 514.000 ;
        RECT 2104.660 510.000 2105.010 510.340 ;
        RECT 2104.660 142.110 2104.800 510.000 ;
        RECT 517.140 141.790 517.400 142.110 ;
        RECT 2104.600 141.790 2104.860 142.110 ;
        RECT 517.200 16.990 517.340 141.790 ;
        RECT 513.920 16.670 514.180 16.990 ;
        RECT 517.140 16.670 517.400 16.990 ;
        RECT 513.980 2.400 514.120 16.670 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 369.820 538.130 369.880 ;
        RECT 669.370 369.820 669.690 369.880 ;
        RECT 537.810 369.680 669.690 369.820 ;
        RECT 537.810 369.620 538.130 369.680 ;
        RECT 669.370 369.620 669.690 369.680 ;
        RECT 531.830 16.900 532.150 16.960 ;
        RECT 538.270 16.900 538.590 16.960 ;
        RECT 531.830 16.760 538.590 16.900 ;
        RECT 531.830 16.700 532.150 16.760 ;
        RECT 538.270 16.700 538.590 16.760 ;
      LAYER via ;
        RECT 537.840 369.620 538.100 369.880 ;
        RECT 669.400 369.620 669.660 369.880 ;
        RECT 531.860 16.700 532.120 16.960 ;
        RECT 538.300 16.700 538.560 16.960 ;
      LAYER met2 ;
        RECT 671.370 510.410 671.650 514.000 ;
        RECT 669.460 510.270 671.650 510.410 ;
        RECT 669.460 369.910 669.600 510.270 ;
        RECT 671.370 510.000 671.650 510.270 ;
        RECT 537.840 369.590 538.100 369.910 ;
        RECT 669.400 369.590 669.660 369.910 ;
        RECT 537.900 18.090 538.040 369.590 ;
        RECT 537.900 17.950 538.500 18.090 ;
        RECT 538.360 16.990 538.500 17.950 ;
        RECT 531.860 16.670 532.120 16.990 ;
        RECT 538.300 16.670 538.560 16.990 ;
        RECT 531.920 2.400 532.060 16.670 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2519.490 1890.980 2519.810 1891.040 ;
        RECT 2534.670 1890.980 2534.990 1891.040 ;
        RECT 2519.490 1890.840 2534.990 1890.980 ;
        RECT 2519.490 1890.780 2519.810 1890.840 ;
        RECT 2534.670 1890.780 2534.990 1890.840 ;
        RECT 551.150 217.500 551.470 217.560 ;
        RECT 2534.670 217.500 2534.990 217.560 ;
        RECT 551.150 217.360 2534.990 217.500 ;
        RECT 551.150 217.300 551.470 217.360 ;
        RECT 2534.670 217.300 2534.990 217.360 ;
      LAYER via ;
        RECT 2519.520 1890.780 2519.780 1891.040 ;
        RECT 2534.700 1890.780 2534.960 1891.040 ;
        RECT 551.180 217.300 551.440 217.560 ;
        RECT 2534.700 217.300 2534.960 217.560 ;
      LAYER met2 ;
        RECT 2519.520 1890.925 2519.780 1891.070 ;
        RECT 2519.510 1890.555 2519.790 1890.925 ;
        RECT 2534.700 1890.750 2534.960 1891.070 ;
        RECT 2534.760 217.590 2534.900 1890.750 ;
        RECT 551.180 217.270 551.440 217.590 ;
        RECT 2534.700 217.270 2534.960 217.590 ;
        RECT 551.240 17.410 551.380 217.270 ;
        RECT 549.860 17.270 551.380 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 2519.510 1890.600 2519.790 1890.880 ;
      LAYER met3 ;
        RECT 2506.000 1890.890 2510.000 1891.040 ;
        RECT 2519.485 1890.890 2519.815 1890.905 ;
        RECT 2506.000 1890.590 2519.815 1890.890 ;
        RECT 2506.000 1890.440 2510.000 1890.590 ;
        RECT 2519.485 1890.575 2519.815 1890.590 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 46.820 568.030 46.880 ;
        RECT 1683.670 46.820 1683.990 46.880 ;
        RECT 567.710 46.680 1683.990 46.820 ;
        RECT 567.710 46.620 568.030 46.680 ;
        RECT 1683.670 46.620 1683.990 46.680 ;
      LAYER via ;
        RECT 567.740 46.620 568.000 46.880 ;
        RECT 1683.700 46.620 1683.960 46.880 ;
      LAYER met2 ;
        RECT 1685.210 510.410 1685.490 514.000 ;
        RECT 1683.760 510.270 1685.490 510.410 ;
        RECT 1683.760 46.910 1683.900 510.270 ;
        RECT 1685.210 510.000 1685.490 510.270 ;
        RECT 567.740 46.590 568.000 46.910 ;
        RECT 1683.700 46.590 1683.960 46.910 ;
        RECT 567.800 2.400 567.940 46.590 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 748.490 500.040 748.810 500.100 ;
        RECT 1301.410 500.040 1301.730 500.100 ;
        RECT 748.490 499.900 1301.730 500.040 ;
        RECT 748.490 499.840 748.810 499.900 ;
        RECT 1301.410 499.840 1301.730 499.900 ;
        RECT 585.650 37.980 585.970 38.040 ;
        RECT 748.490 37.980 748.810 38.040 ;
        RECT 585.650 37.840 748.810 37.980 ;
        RECT 585.650 37.780 585.970 37.840 ;
        RECT 748.490 37.780 748.810 37.840 ;
      LAYER via ;
        RECT 748.520 499.840 748.780 500.100 ;
        RECT 1301.440 499.840 1301.700 500.100 ;
        RECT 585.680 37.780 585.940 38.040 ;
        RECT 748.520 37.780 748.780 38.040 ;
      LAYER met2 ;
        RECT 1301.570 510.340 1301.850 514.000 ;
        RECT 1301.500 510.000 1301.850 510.340 ;
        RECT 1301.500 500.130 1301.640 510.000 ;
        RECT 748.520 499.810 748.780 500.130 ;
        RECT 1301.440 499.810 1301.700 500.130 ;
        RECT 748.580 38.070 748.720 499.810 ;
        RECT 585.680 37.750 585.940 38.070 ;
        RECT 748.520 37.750 748.780 38.070 ;
        RECT 585.740 2.400 585.880 37.750 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 369.140 96.530 369.200 ;
        RECT 1690.570 369.140 1690.890 369.200 ;
        RECT 96.210 369.000 1690.890 369.140 ;
        RECT 96.210 368.940 96.530 369.000 ;
        RECT 1690.570 368.940 1690.890 369.000 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 96.210 17.580 96.530 17.640 ;
        RECT 91.610 17.440 96.530 17.580 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 96.210 17.380 96.530 17.440 ;
      LAYER via ;
        RECT 96.240 368.940 96.500 369.200 ;
        RECT 1690.600 368.940 1690.860 369.200 ;
        RECT 91.640 17.380 91.900 17.640 ;
        RECT 96.240 17.380 96.500 17.640 ;
      LAYER met2 ;
        RECT 1697.170 510.410 1697.450 514.000 ;
        RECT 1690.660 510.270 1697.450 510.410 ;
        RECT 1690.660 369.230 1690.800 510.270 ;
        RECT 1697.170 510.000 1697.450 510.270 ;
        RECT 96.240 368.910 96.500 369.230 ;
        RECT 1690.600 368.910 1690.860 369.230 ;
        RECT 96.300 17.670 96.440 368.910 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 96.240 17.350 96.500 17.670 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 600.370 2.960 600.690 3.020 ;
        RECT 603.130 2.960 603.450 3.020 ;
        RECT 600.370 2.820 603.450 2.960 ;
        RECT 600.370 2.760 600.690 2.820 ;
        RECT 603.130 2.760 603.450 2.820 ;
      LAYER via ;
        RECT 600.400 2.760 600.660 3.020 ;
        RECT 603.160 2.760 603.420 3.020 ;
      LAYER met2 ;
        RECT 600.390 494.515 600.670 494.885 ;
        RECT 600.460 3.050 600.600 494.515 ;
        RECT 600.400 2.730 600.660 3.050 ;
        RECT 603.160 2.730 603.420 3.050 ;
        RECT 603.220 2.400 603.360 2.730 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 600.390 494.560 600.670 494.840 ;
      LAYER met3 ;
        RECT 410.000 2339.240 414.000 2339.840 ;
        RECT 412.470 2338.340 412.770 2339.240 ;
        RECT 412.430 2338.020 412.810 2338.340 ;
        RECT 416.110 494.850 416.490 494.860 ;
        RECT 600.365 494.850 600.695 494.865 ;
        RECT 416.110 494.550 600.695 494.850 ;
        RECT 416.110 494.540 416.490 494.550 ;
        RECT 600.365 494.535 600.695 494.550 ;
      LAYER via3 ;
        RECT 412.460 2338.020 412.780 2338.340 ;
        RECT 416.140 494.540 416.460 494.860 ;
      LAYER met4 ;
        RECT 412.455 2338.015 412.785 2338.345 ;
        RECT 412.470 2337.650 412.770 2338.015 ;
        RECT 412.470 2337.350 416.450 2337.650 ;
        RECT 416.150 494.865 416.450 2337.350 ;
        RECT 416.135 494.535 416.465 494.865 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.510 86.600 627.830 86.660 ;
        RECT 2263.270 86.600 2263.590 86.660 ;
        RECT 627.510 86.460 2263.590 86.600 ;
        RECT 627.510 86.400 627.830 86.460 ;
        RECT 2263.270 86.400 2263.590 86.460 ;
        RECT 621.070 16.900 621.390 16.960 ;
        RECT 627.510 16.900 627.830 16.960 ;
        RECT 621.070 16.760 627.830 16.900 ;
        RECT 621.070 16.700 621.390 16.760 ;
        RECT 627.510 16.700 627.830 16.760 ;
      LAYER via ;
        RECT 627.540 86.400 627.800 86.660 ;
        RECT 2263.300 86.400 2263.560 86.660 ;
        RECT 621.100 16.700 621.360 16.960 ;
        RECT 627.540 16.700 627.800 16.960 ;
      LAYER met2 ;
        RECT 2265.730 510.410 2266.010 514.000 ;
        RECT 2263.360 510.270 2266.010 510.410 ;
        RECT 2263.360 86.690 2263.500 510.270 ;
        RECT 2265.730 510.000 2266.010 510.270 ;
        RECT 627.540 86.370 627.800 86.690 ;
        RECT 2263.300 86.370 2263.560 86.690 ;
        RECT 627.600 16.990 627.740 86.370 ;
        RECT 621.100 16.670 621.360 16.990 ;
        RECT 627.540 16.670 627.800 16.990 ;
        RECT 621.160 2.400 621.300 16.670 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1579.730 3009.835 1580.010 3010.205 ;
        RECT 1579.800 3009.410 1579.940 3009.835 ;
        RECT 1580.330 3009.410 1580.610 3010.000 ;
        RECT 1579.800 3009.270 1580.610 3009.410 ;
        RECT 1580.330 3006.000 1580.610 3009.270 ;
        RECT 115.550 18.515 115.830 18.885 ;
        RECT 115.620 2.400 115.760 18.515 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1579.730 3009.880 1580.010 3010.160 ;
        RECT 115.550 18.560 115.830 18.840 ;
      LAYER met3 ;
        RECT 375.630 3010.170 376.010 3010.180 ;
        RECT 1579.705 3010.170 1580.035 3010.185 ;
        RECT 375.630 3009.870 1580.035 3010.170 ;
        RECT 375.630 3009.860 376.010 3009.870 ;
        RECT 1579.705 3009.855 1580.035 3009.870 ;
        RECT 115.525 18.850 115.855 18.865 ;
        RECT 375.630 18.850 376.010 18.860 ;
        RECT 115.525 18.550 376.010 18.850 ;
        RECT 115.525 18.535 115.855 18.550 ;
        RECT 375.630 18.540 376.010 18.550 ;
      LAYER via3 ;
        RECT 375.660 3009.860 375.980 3010.180 ;
        RECT 375.660 18.540 375.980 18.860 ;
      LAYER met4 ;
        RECT 375.655 3009.855 375.985 3010.185 ;
        RECT 375.670 18.865 375.970 3009.855 ;
        RECT 375.655 18.535 375.985 18.865 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.990 500.380 714.310 500.440 ;
        RECT 993.210 500.380 993.530 500.440 ;
        RECT 713.990 500.240 993.530 500.380 ;
        RECT 713.990 500.180 714.310 500.240 ;
        RECT 993.210 500.180 993.530 500.240 ;
        RECT 144.510 114.140 144.830 114.200 ;
        RECT 713.990 114.140 714.310 114.200 ;
        RECT 144.510 114.000 714.310 114.140 ;
        RECT 144.510 113.940 144.830 114.000 ;
        RECT 713.990 113.940 714.310 114.000 ;
        RECT 139.450 17.580 139.770 17.640 ;
        RECT 144.510 17.580 144.830 17.640 ;
        RECT 139.450 17.440 144.830 17.580 ;
        RECT 139.450 17.380 139.770 17.440 ;
        RECT 144.510 17.380 144.830 17.440 ;
      LAYER via ;
        RECT 714.020 500.180 714.280 500.440 ;
        RECT 993.240 500.180 993.500 500.440 ;
        RECT 144.540 113.940 144.800 114.200 ;
        RECT 714.020 113.940 714.280 114.200 ;
        RECT 139.480 17.380 139.740 17.640 ;
        RECT 144.540 17.380 144.800 17.640 ;
      LAYER met2 ;
        RECT 993.370 510.340 993.650 514.000 ;
        RECT 993.300 510.000 993.650 510.340 ;
        RECT 993.300 500.470 993.440 510.000 ;
        RECT 714.020 500.150 714.280 500.470 ;
        RECT 993.240 500.150 993.500 500.470 ;
        RECT 714.080 114.230 714.220 500.150 ;
        RECT 144.540 113.910 144.800 114.230 ;
        RECT 714.020 113.910 714.280 114.230 ;
        RECT 144.600 17.670 144.740 113.910 ;
        RECT 139.480 17.350 139.740 17.670 ;
        RECT 144.540 17.350 144.800 17.670 ;
        RECT 139.540 2.400 139.680 17.350 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 3013.320 158.630 3013.380 ;
        RECT 1197.450 3013.320 1197.770 3013.380 ;
        RECT 158.310 3013.180 1197.770 3013.320 ;
        RECT 158.310 3013.120 158.630 3013.180 ;
        RECT 1197.450 3013.120 1197.770 3013.180 ;
      LAYER via ;
        RECT 158.340 3013.120 158.600 3013.380 ;
        RECT 1197.480 3013.120 1197.740 3013.380 ;
      LAYER met2 ;
        RECT 158.340 3013.090 158.600 3013.410 ;
        RECT 1197.480 3013.090 1197.740 3013.410 ;
        RECT 158.400 17.410 158.540 3013.090 ;
        RECT 1197.540 3010.000 1197.680 3013.090 ;
        RECT 1197.540 3009.340 1197.890 3010.000 ;
        RECT 1197.610 3006.000 1197.890 3009.340 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 17.580 175.190 17.640 ;
        RECT 179.010 17.580 179.330 17.640 ;
        RECT 174.870 17.440 179.330 17.580 ;
        RECT 174.870 17.380 175.190 17.440 ;
        RECT 179.010 17.380 179.330 17.440 ;
      LAYER via ;
        RECT 174.900 17.380 175.160 17.640 ;
        RECT 179.040 17.380 179.300 17.640 ;
      LAYER met2 ;
        RECT 2198.430 3020.715 2198.710 3021.085 ;
        RECT 2198.500 3010.000 2198.640 3020.715 ;
        RECT 2198.500 3009.340 2198.850 3010.000 ;
        RECT 2198.570 3006.000 2198.850 3009.340 ;
        RECT 179.030 2977.195 179.310 2977.565 ;
        RECT 179.100 17.670 179.240 2977.195 ;
        RECT 174.900 17.350 175.160 17.670 ;
        RECT 179.040 17.350 179.300 17.670 ;
        RECT 174.960 2.400 175.100 17.350 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 2198.430 3020.760 2198.710 3021.040 ;
        RECT 179.030 2977.240 179.310 2977.520 ;
      LAYER met3 ;
        RECT 542.150 3021.050 542.530 3021.060 ;
        RECT 548.590 3021.050 548.970 3021.060 ;
        RECT 542.150 3020.750 548.970 3021.050 ;
        RECT 542.150 3020.740 542.530 3020.750 ;
        RECT 548.590 3020.740 548.970 3020.750 ;
        RECT 737.190 3021.050 737.570 3021.060 ;
        RECT 789.630 3021.050 790.010 3021.060 ;
        RECT 737.190 3020.750 790.010 3021.050 ;
        RECT 737.190 3020.740 737.570 3020.750 ;
        RECT 789.630 3020.740 790.010 3020.750 ;
        RECT 1118.070 3021.050 1118.450 3021.060 ;
        RECT 1124.510 3021.050 1124.890 3021.060 ;
        RECT 1118.070 3020.750 1124.890 3021.050 ;
        RECT 1118.070 3020.740 1118.450 3020.750 ;
        RECT 1124.510 3020.740 1124.890 3020.750 ;
        RECT 1316.790 3021.050 1317.170 3021.060 ;
        RECT 1322.310 3021.050 1322.690 3021.060 ;
        RECT 1316.790 3020.750 1322.690 3021.050 ;
        RECT 1316.790 3020.740 1317.170 3020.750 ;
        RECT 1322.310 3020.740 1322.690 3020.750 ;
        RECT 1406.030 3021.050 1406.410 3021.060 ;
        RECT 1415.230 3021.050 1415.610 3021.060 ;
        RECT 1406.030 3020.750 1415.610 3021.050 ;
        RECT 1406.030 3020.740 1406.410 3020.750 ;
        RECT 1415.230 3020.740 1415.610 3020.750 ;
        RECT 1892.710 3021.050 1893.090 3021.060 ;
        RECT 1945.150 3021.050 1945.530 3021.060 ;
        RECT 1892.710 3020.750 1945.530 3021.050 ;
        RECT 1892.710 3020.740 1893.090 3020.750 ;
        RECT 1945.150 3020.740 1945.530 3020.750 ;
        RECT 2072.110 3021.050 2072.490 3021.060 ;
        RECT 2107.990 3021.050 2108.370 3021.060 ;
        RECT 2072.110 3020.750 2108.370 3021.050 ;
        RECT 2072.110 3020.740 2072.490 3020.750 ;
        RECT 2107.990 3020.740 2108.370 3020.750 ;
        RECT 2186.190 3021.050 2186.570 3021.060 ;
        RECT 2198.405 3021.050 2198.735 3021.065 ;
        RECT 2186.190 3020.750 2198.735 3021.050 ;
        RECT 2186.190 3020.740 2186.570 3020.750 ;
        RECT 2198.405 3020.735 2198.735 3020.750 ;
        RECT 179.005 2977.530 179.335 2977.545 ;
        RECT 412.430 2977.530 412.810 2977.540 ;
        RECT 179.005 2977.230 412.810 2977.530 ;
        RECT 179.005 2977.215 179.335 2977.230 ;
        RECT 412.430 2977.220 412.810 2977.230 ;
      LAYER via3 ;
        RECT 542.180 3020.740 542.500 3021.060 ;
        RECT 548.620 3020.740 548.940 3021.060 ;
        RECT 737.220 3020.740 737.540 3021.060 ;
        RECT 789.660 3020.740 789.980 3021.060 ;
        RECT 1118.100 3020.740 1118.420 3021.060 ;
        RECT 1124.540 3020.740 1124.860 3021.060 ;
        RECT 1316.820 3020.740 1317.140 3021.060 ;
        RECT 1322.340 3020.740 1322.660 3021.060 ;
        RECT 1406.060 3020.740 1406.380 3021.060 ;
        RECT 1415.260 3020.740 1415.580 3021.060 ;
        RECT 1892.740 3020.740 1893.060 3021.060 ;
        RECT 1945.180 3020.740 1945.500 3021.060 ;
        RECT 2072.140 3020.740 2072.460 3021.060 ;
        RECT 2108.020 3020.740 2108.340 3021.060 ;
        RECT 2186.220 3020.740 2186.540 3021.060 ;
        RECT 412.460 2977.220 412.780 2977.540 ;
      LAYER met4 ;
        RECT 789.230 3023.710 790.410 3024.890 ;
        RECT 415.710 3020.310 416.890 3021.490 ;
        RECT 541.750 3020.310 542.930 3021.490 ;
        RECT 548.190 3020.310 549.370 3021.490 ;
        RECT 736.790 3020.310 737.970 3021.490 ;
        RECT 789.670 3021.065 789.970 3023.710 ;
        RECT 789.655 3020.735 789.985 3021.065 ;
        RECT 1024.750 3021.050 1025.930 3021.490 ;
        RECT 1028.430 3021.050 1029.610 3021.490 ;
        RECT 1024.750 3020.750 1029.610 3021.050 ;
        RECT 1024.750 3020.310 1025.930 3020.750 ;
        RECT 1028.430 3020.310 1029.610 3020.750 ;
        RECT 1117.670 3020.310 1118.850 3021.490 ;
        RECT 1124.110 3020.310 1125.290 3021.490 ;
        RECT 1217.950 3021.050 1219.130 3021.490 ;
        RECT 1221.630 3021.050 1222.810 3021.490 ;
        RECT 1217.950 3020.750 1222.810 3021.050 ;
        RECT 1217.950 3020.310 1219.130 3020.750 ;
        RECT 1221.630 3020.310 1222.810 3020.750 ;
        RECT 1316.390 3020.310 1317.570 3021.490 ;
        RECT 1321.910 3020.310 1323.090 3021.490 ;
        RECT 1405.630 3020.310 1406.810 3021.490 ;
        RECT 1414.830 3020.310 1416.010 3021.490 ;
        RECT 1507.750 3021.050 1508.930 3021.490 ;
        RECT 1511.430 3021.050 1512.610 3021.490 ;
        RECT 1507.750 3020.750 1512.610 3021.050 ;
        RECT 1507.750 3020.310 1508.930 3020.750 ;
        RECT 1511.430 3020.310 1512.610 3020.750 ;
        RECT 1604.350 3021.050 1605.530 3021.490 ;
        RECT 1608.030 3021.050 1609.210 3021.490 ;
        RECT 1604.350 3020.750 1609.210 3021.050 ;
        RECT 1604.350 3020.310 1605.530 3020.750 ;
        RECT 1608.030 3020.310 1609.210 3020.750 ;
        RECT 1700.950 3021.050 1702.130 3021.490 ;
        RECT 1704.630 3021.050 1705.810 3021.490 ;
        RECT 1700.950 3020.750 1705.810 3021.050 ;
        RECT 1700.950 3020.310 1702.130 3020.750 ;
        RECT 1704.630 3020.310 1705.810 3020.750 ;
        RECT 1797.550 3021.050 1798.730 3021.490 ;
        RECT 1801.230 3021.050 1802.410 3021.490 ;
        RECT 1797.550 3020.750 1802.410 3021.050 ;
        RECT 1797.550 3020.310 1798.730 3020.750 ;
        RECT 1801.230 3020.310 1802.410 3020.750 ;
        RECT 1892.310 3020.310 1893.490 3021.490 ;
        RECT 1944.750 3020.310 1945.930 3021.490 ;
        RECT 2071.710 3020.310 2072.890 3021.490 ;
        RECT 2107.590 3020.310 2108.770 3021.490 ;
        RECT 2185.790 3020.310 2186.970 3021.490 ;
        RECT 416.150 2980.250 416.450 3020.310 ;
        RECT 414.310 2979.950 416.450 2980.250 ;
        RECT 412.455 2977.215 412.785 2977.545 ;
        RECT 412.470 2976.850 412.770 2977.215 ;
        RECT 414.310 2976.850 414.610 2979.950 ;
        RECT 412.470 2976.550 414.610 2976.850 ;
      LAYER met5 ;
        RECT 789.020 3023.500 884.460 3025.100 ;
        RECT 882.860 3021.700 884.460 3023.500 ;
        RECT 1992.380 3021.700 1994.900 3025.100 ;
        RECT 415.500 3020.100 543.140 3021.700 ;
        RECT 547.980 3020.100 738.180 3021.700 ;
        RECT 882.860 3020.100 1026.140 3021.700 ;
        RECT 1028.220 3020.100 1119.060 3021.700 ;
        RECT 1123.900 3020.100 1219.340 3021.700 ;
        RECT 1221.420 3020.100 1317.780 3021.700 ;
        RECT 1321.700 3020.100 1407.020 3021.700 ;
        RECT 1414.620 3020.100 1509.140 3021.700 ;
        RECT 1511.220 3020.100 1605.740 3021.700 ;
        RECT 1607.820 3020.100 1702.340 3021.700 ;
        RECT 1704.420 3020.100 1798.940 3021.700 ;
        RECT 1801.020 3020.100 1893.700 3021.700 ;
        RECT 1944.540 3020.100 2073.100 3021.700 ;
        RECT 2107.380 3020.100 2187.180 3021.700 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 2097.700 231.310 2097.760 ;
        RECT 393.370 2097.700 393.690 2097.760 ;
        RECT 230.990 2097.560 393.690 2097.700 ;
        RECT 230.990 2097.500 231.310 2097.560 ;
        RECT 393.370 2097.500 393.690 2097.560 ;
        RECT 192.350 30.840 192.670 30.900 ;
        RECT 230.990 30.840 231.310 30.900 ;
        RECT 192.350 30.700 231.310 30.840 ;
        RECT 192.350 30.640 192.670 30.700 ;
        RECT 230.990 30.640 231.310 30.700 ;
      LAYER via ;
        RECT 231.020 2097.500 231.280 2097.760 ;
        RECT 393.400 2097.500 393.660 2097.760 ;
        RECT 192.380 30.640 192.640 30.900 ;
        RECT 231.020 30.640 231.280 30.900 ;
      LAYER met2 ;
        RECT 393.390 2102.715 393.670 2103.085 ;
        RECT 393.460 2097.790 393.600 2102.715 ;
        RECT 231.020 2097.470 231.280 2097.790 ;
        RECT 393.400 2097.470 393.660 2097.790 ;
        RECT 231.080 30.930 231.220 2097.470 ;
        RECT 192.380 30.610 192.640 30.930 ;
        RECT 231.020 30.610 231.280 30.930 ;
        RECT 192.440 15.370 192.580 30.610 ;
        RECT 192.440 15.230 193.040 15.370 ;
        RECT 192.900 2.400 193.040 15.230 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 393.390 2102.760 393.670 2103.040 ;
      LAYER met3 ;
        RECT 393.365 2103.050 393.695 2103.065 ;
        RECT 410.000 2103.050 414.000 2103.200 ;
        RECT 393.365 2102.750 414.000 2103.050 ;
        RECT 393.365 2102.735 393.695 2102.750 ;
        RECT 410.000 2102.600 414.000 2102.750 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 415.910 3016.380 416.230 3016.440 ;
        RECT 1308.770 3016.380 1309.090 3016.440 ;
        RECT 415.910 3016.240 1309.090 3016.380 ;
        RECT 415.910 3016.180 416.230 3016.240 ;
        RECT 1308.770 3016.180 1309.090 3016.240 ;
        RECT 213.510 2963.340 213.830 2963.400 ;
        RECT 414.530 2963.340 414.850 2963.400 ;
        RECT 213.510 2963.200 414.850 2963.340 ;
        RECT 213.510 2963.140 213.830 2963.200 ;
        RECT 414.530 2963.140 414.850 2963.200 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 415.940 3016.180 416.200 3016.440 ;
        RECT 1308.800 3016.180 1309.060 3016.440 ;
        RECT 213.540 2963.140 213.800 2963.400 ;
        RECT 414.560 2963.140 414.820 2963.400 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 415.940 3016.150 416.200 3016.470 ;
        RECT 1308.800 3016.150 1309.060 3016.470 ;
        RECT 416.000 2963.850 416.140 3016.150 ;
        RECT 1308.860 3010.000 1309.000 3016.150 ;
        RECT 1308.860 3009.340 1309.210 3010.000 ;
        RECT 1308.930 3006.000 1309.210 3009.340 ;
        RECT 414.620 2963.710 416.140 2963.850 ;
        RECT 414.620 2963.430 414.760 2963.710 ;
        RECT 213.540 2963.110 213.800 2963.430 ;
        RECT 414.560 2963.110 414.820 2963.430 ;
        RECT 213.600 17.670 213.740 2963.110 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 233.750 59.740 234.070 59.800 ;
        RECT 2325.370 59.740 2325.690 59.800 ;
        RECT 233.750 59.600 2325.690 59.740 ;
        RECT 233.750 59.540 234.070 59.600 ;
        RECT 2325.370 59.540 2325.690 59.600 ;
        RECT 228.690 17.580 229.010 17.640 ;
        RECT 233.750 17.580 234.070 17.640 ;
        RECT 228.690 17.440 234.070 17.580 ;
        RECT 228.690 17.380 229.010 17.440 ;
        RECT 233.750 17.380 234.070 17.440 ;
      LAYER via ;
        RECT 233.780 59.540 234.040 59.800 ;
        RECT 2325.400 59.540 2325.660 59.800 ;
        RECT 228.720 17.380 228.980 17.640 ;
        RECT 233.780 17.380 234.040 17.640 ;
      LAYER met2 ;
        RECT 2327.370 510.410 2327.650 514.000 ;
        RECT 2325.460 510.270 2327.650 510.410 ;
        RECT 2325.460 59.830 2325.600 510.270 ;
        RECT 2327.370 510.000 2327.650 510.270 ;
        RECT 233.780 59.510 234.040 59.830 ;
        RECT 2325.400 59.510 2325.660 59.830 ;
        RECT 233.840 17.670 233.980 59.510 ;
        RECT 228.720 17.350 228.980 17.670 ;
        RECT 233.780 17.350 234.040 17.670 ;
        RECT 228.780 2.400 228.920 17.350 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 189.590 1808.020 189.910 1808.080 ;
        RECT 393.370 1808.020 393.690 1808.080 ;
        RECT 189.590 1807.880 393.690 1808.020 ;
        RECT 189.590 1807.820 189.910 1807.880 ;
        RECT 393.370 1807.820 393.690 1807.880 ;
        RECT 54.810 72.320 55.130 72.380 ;
        RECT 189.590 72.320 189.910 72.380 ;
        RECT 54.810 72.180 189.910 72.320 ;
        RECT 54.810 72.120 55.130 72.180 ;
        RECT 189.590 72.120 189.910 72.180 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 189.620 1807.820 189.880 1808.080 ;
        RECT 393.400 1807.820 393.660 1808.080 ;
        RECT 54.840 72.120 55.100 72.380 ;
        RECT 189.620 72.120 189.880 72.380 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 393.390 1810.315 393.670 1810.685 ;
        RECT 393.460 1808.110 393.600 1810.315 ;
        RECT 189.620 1807.790 189.880 1808.110 ;
        RECT 393.400 1807.790 393.660 1808.110 ;
        RECT 189.680 72.410 189.820 1807.790 ;
        RECT 54.840 72.090 55.100 72.410 ;
        RECT 189.620 72.090 189.880 72.410 ;
        RECT 54.900 17.670 55.040 72.090 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 393.390 1810.360 393.670 1810.640 ;
      LAYER met3 ;
        RECT 393.365 1810.650 393.695 1810.665 ;
        RECT 410.000 1810.650 414.000 1810.800 ;
        RECT 393.365 1810.350 414.000 1810.650 ;
        RECT 393.365 1810.335 393.695 1810.350 ;
        RECT 410.000 1810.200 414.000 1810.350 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2473.490 496.980 2473.810 497.040 ;
        RECT 2500.170 496.980 2500.490 497.040 ;
        RECT 2473.490 496.840 2500.490 496.980 ;
        RECT 2473.490 496.780 2473.810 496.840 ;
        RECT 2500.170 496.780 2500.490 496.840 ;
        RECT 254.910 59.400 255.230 59.460 ;
        RECT 2473.490 59.400 2473.810 59.460 ;
        RECT 254.910 59.260 2473.810 59.400 ;
        RECT 254.910 59.200 255.230 59.260 ;
        RECT 2473.490 59.200 2473.810 59.260 ;
        RECT 252.610 14.520 252.930 14.580 ;
        RECT 254.910 14.520 255.230 14.580 ;
        RECT 252.610 14.380 255.230 14.520 ;
        RECT 252.610 14.320 252.930 14.380 ;
        RECT 254.910 14.320 255.230 14.380 ;
      LAYER via ;
        RECT 2473.520 496.780 2473.780 497.040 ;
        RECT 2500.200 496.780 2500.460 497.040 ;
        RECT 254.940 59.200 255.200 59.460 ;
        RECT 2473.520 59.200 2473.780 59.460 ;
        RECT 252.640 14.320 252.900 14.580 ;
        RECT 254.940 14.320 255.200 14.580 ;
      LAYER met2 ;
        RECT 2500.330 510.340 2500.610 514.000 ;
        RECT 2500.260 510.000 2500.610 510.340 ;
        RECT 2500.260 497.070 2500.400 510.000 ;
        RECT 2473.520 496.750 2473.780 497.070 ;
        RECT 2500.200 496.750 2500.460 497.070 ;
        RECT 2473.580 59.490 2473.720 496.750 ;
        RECT 254.940 59.170 255.200 59.490 ;
        RECT 2473.520 59.170 2473.780 59.490 ;
        RECT 255.000 14.610 255.140 59.170 ;
        RECT 252.640 14.290 252.900 14.610 ;
        RECT 254.940 14.290 255.200 14.610 ;
        RECT 252.700 2.400 252.840 14.290 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 38.320 270.410 38.380 ;
        RECT 1497.370 38.320 1497.690 38.380 ;
        RECT 270.090 38.180 1497.690 38.320 ;
        RECT 270.090 38.120 270.410 38.180 ;
        RECT 1497.370 38.120 1497.690 38.180 ;
      LAYER via ;
        RECT 270.120 38.120 270.380 38.380 ;
        RECT 1497.400 38.120 1497.660 38.380 ;
      LAYER met2 ;
        RECT 1499.370 510.410 1499.650 514.000 ;
        RECT 1497.460 510.270 1499.650 510.410 ;
        RECT 1497.460 38.410 1497.600 510.270 ;
        RECT 1499.370 510.000 1499.650 510.270 ;
        RECT 270.120 38.090 270.380 38.410 ;
        RECT 1497.400 38.090 1497.660 38.410 ;
        RECT 270.180 2.400 270.320 38.090 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 1332.020 288.810 1332.080 ;
        RECT 393.370 1332.020 393.690 1332.080 ;
        RECT 288.490 1331.880 393.690 1332.020 ;
        RECT 288.490 1331.820 288.810 1331.880 ;
        RECT 393.370 1331.820 393.690 1331.880 ;
      LAYER via ;
        RECT 288.520 1331.820 288.780 1332.080 ;
        RECT 393.400 1331.820 393.660 1332.080 ;
      LAYER met2 ;
        RECT 393.390 1335.675 393.670 1336.045 ;
        RECT 393.460 1332.110 393.600 1335.675 ;
        RECT 288.520 1331.790 288.780 1332.110 ;
        RECT 393.400 1331.790 393.660 1332.110 ;
        RECT 288.580 3.130 288.720 1331.790 ;
        RECT 288.120 2.990 288.720 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 393.390 1335.720 393.670 1336.000 ;
      LAYER met3 ;
        RECT 393.365 1336.010 393.695 1336.025 ;
        RECT 410.000 1336.010 414.000 1336.160 ;
        RECT 393.365 1335.710 414.000 1336.010 ;
        RECT 393.365 1335.695 393.695 1335.710 ;
        RECT 410.000 1335.560 414.000 1335.710 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 565.945 3002.625 566.115 3006.535 ;
      LAYER mcon ;
        RECT 565.945 3006.365 566.115 3006.535 ;
      LAYER met1 ;
        RECT 565.870 3006.520 566.190 3006.580 ;
        RECT 565.675 3006.380 566.190 3006.520 ;
        RECT 565.870 3006.320 566.190 3006.380 ;
        RECT 310.110 3002.780 310.430 3002.840 ;
        RECT 565.885 3002.780 566.175 3002.825 ;
        RECT 310.110 3002.640 566.175 3002.780 ;
        RECT 310.110 3002.580 310.430 3002.640 ;
        RECT 565.885 3002.595 566.175 3002.640 ;
        RECT 305.970 17.580 306.290 17.640 ;
        RECT 310.110 17.580 310.430 17.640 ;
        RECT 305.970 17.440 310.430 17.580 ;
        RECT 305.970 17.380 306.290 17.440 ;
        RECT 310.110 17.380 310.430 17.440 ;
      LAYER via ;
        RECT 565.900 3006.320 566.160 3006.580 ;
        RECT 310.140 3002.580 310.400 3002.840 ;
        RECT 306.000 17.380 306.260 17.640 ;
        RECT 310.140 17.380 310.400 17.640 ;
      LAYER met2 ;
        RECT 567.410 3006.690 567.690 3010.000 ;
        RECT 565.960 3006.610 567.690 3006.690 ;
        RECT 565.900 3006.550 567.690 3006.610 ;
        RECT 565.900 3006.290 566.160 3006.550 ;
        RECT 567.410 3006.000 567.690 3006.550 ;
        RECT 310.140 3002.550 310.400 3002.870 ;
        RECT 310.200 17.670 310.340 3002.550 ;
        RECT 306.000 17.350 306.260 17.670 ;
        RECT 310.140 17.350 310.400 17.670 ;
        RECT 306.060 2.400 306.200 17.350 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.670 3015.275 2494.950 3015.645 ;
        RECT 2494.740 3010.000 2494.880 3015.275 ;
        RECT 2494.740 3009.340 2495.090 3010.000 ;
        RECT 2494.810 3006.000 2495.090 3009.340 ;
        RECT 323.010 57.955 323.290 58.325 ;
        RECT 323.080 17.410 323.220 57.955 ;
        RECT 323.080 17.270 324.140 17.410 ;
        RECT 324.000 2.400 324.140 17.270 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 2494.670 3015.320 2494.950 3015.600 ;
        RECT 323.010 58.000 323.290 58.280 ;
      LAYER met3 ;
        RECT 2479.670 3015.610 2480.050 3015.620 ;
        RECT 2494.645 3015.610 2494.975 3015.625 ;
        RECT 2479.670 3015.310 2494.975 3015.610 ;
        RECT 2479.670 3015.300 2480.050 3015.310 ;
        RECT 2494.645 3015.295 2494.975 3015.310 ;
        RECT 322.985 58.290 323.315 58.305 ;
        RECT 2479.670 58.290 2480.050 58.300 ;
        RECT 322.985 57.990 2480.050 58.290 ;
        RECT 322.985 57.975 323.315 57.990 ;
        RECT 2479.670 57.980 2480.050 57.990 ;
      LAYER via3 ;
        RECT 2479.700 3015.300 2480.020 3015.620 ;
        RECT 2479.700 57.980 2480.020 58.300 ;
      LAYER met4 ;
        RECT 2479.695 3015.295 2480.025 3015.625 ;
        RECT 2479.710 2963.250 2480.010 3015.295 ;
        RECT 2479.710 2962.950 2481.850 2963.250 ;
        RECT 2481.550 2946.930 2481.850 2962.950 ;
        RECT 2479.710 2946.630 2481.850 2946.930 ;
        RECT 2479.710 1675.090 2480.010 2946.630 ;
        RECT 2479.270 1673.910 2480.450 1675.090 ;
        RECT 2482.950 1673.910 2484.130 1675.090 ;
        RECT 2483.390 1667.850 2483.690 1673.910 ;
        RECT 2481.550 1667.550 2483.690 1667.850 ;
        RECT 2481.550 1623.650 2481.850 1667.550 ;
        RECT 2479.710 1623.350 2481.850 1623.650 ;
        RECT 2479.710 58.305 2480.010 1623.350 ;
        RECT 2479.695 57.975 2480.025 58.305 ;
      LAYER met5 ;
        RECT 2479.060 1673.700 2484.340 1675.300 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1617.890 496.980 1618.210 497.040 ;
        RECT 1622.490 496.980 1622.810 497.040 ;
        RECT 1617.890 496.840 1622.810 496.980 ;
        RECT 1617.890 496.780 1618.210 496.840 ;
        RECT 1622.490 496.780 1622.810 496.840 ;
        RECT 344.150 293.660 344.470 293.720 ;
        RECT 1617.890 293.660 1618.210 293.720 ;
        RECT 344.150 293.520 1618.210 293.660 ;
        RECT 344.150 293.460 344.470 293.520 ;
        RECT 1617.890 293.460 1618.210 293.520 ;
        RECT 341.390 17.580 341.710 17.640 ;
        RECT 344.150 17.580 344.470 17.640 ;
        RECT 341.390 17.440 344.470 17.580 ;
        RECT 341.390 17.380 341.710 17.440 ;
        RECT 344.150 17.380 344.470 17.440 ;
      LAYER via ;
        RECT 1617.920 496.780 1618.180 497.040 ;
        RECT 1622.520 496.780 1622.780 497.040 ;
        RECT 344.180 293.460 344.440 293.720 ;
        RECT 1617.920 293.460 1618.180 293.720 ;
        RECT 341.420 17.380 341.680 17.640 ;
        RECT 344.180 17.380 344.440 17.640 ;
      LAYER met2 ;
        RECT 1622.650 510.340 1622.930 514.000 ;
        RECT 1622.580 510.000 1622.930 510.340 ;
        RECT 1622.580 497.070 1622.720 510.000 ;
        RECT 1617.920 496.750 1618.180 497.070 ;
        RECT 1622.520 496.750 1622.780 497.070 ;
        RECT 1617.980 293.750 1618.120 496.750 ;
        RECT 344.180 293.430 344.440 293.750 ;
        RECT 1617.920 293.430 1618.180 293.750 ;
        RECT 344.240 17.670 344.380 293.430 ;
        RECT 341.420 17.350 341.680 17.670 ;
        RECT 344.180 17.350 344.440 17.670 ;
        RECT 341.480 2.400 341.620 17.350 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 624.290 501.060 624.610 501.120 ;
        RECT 634.410 501.060 634.730 501.120 ;
        RECT 624.290 500.920 634.730 501.060 ;
        RECT 624.290 500.860 624.610 500.920 ;
        RECT 634.410 500.860 634.730 500.920 ;
        RECT 364.390 65.520 364.710 65.580 ;
        RECT 624.290 65.520 624.610 65.580 ;
        RECT 364.390 65.380 624.610 65.520 ;
        RECT 364.390 65.320 364.710 65.380 ;
        RECT 624.290 65.320 624.610 65.380 ;
        RECT 359.330 17.580 359.650 17.640 ;
        RECT 364.390 17.580 364.710 17.640 ;
        RECT 359.330 17.440 364.710 17.580 ;
        RECT 359.330 17.380 359.650 17.440 ;
        RECT 364.390 17.380 364.710 17.440 ;
      LAYER via ;
        RECT 624.320 500.860 624.580 501.120 ;
        RECT 634.440 500.860 634.700 501.120 ;
        RECT 364.420 65.320 364.680 65.580 ;
        RECT 624.320 65.320 624.580 65.580 ;
        RECT 359.360 17.380 359.620 17.640 ;
        RECT 364.420 17.380 364.680 17.640 ;
      LAYER met2 ;
        RECT 634.570 510.340 634.850 514.000 ;
        RECT 634.500 510.000 634.850 510.340 ;
        RECT 634.500 501.150 634.640 510.000 ;
        RECT 624.320 500.830 624.580 501.150 ;
        RECT 634.440 500.830 634.700 501.150 ;
        RECT 624.380 65.610 624.520 500.830 ;
        RECT 364.420 65.290 364.680 65.610 ;
        RECT 624.320 65.290 624.580 65.610 ;
        RECT 364.480 17.670 364.620 65.290 ;
        RECT 359.360 17.350 359.620 17.670 ;
        RECT 364.420 17.350 364.680 17.670 ;
        RECT 359.420 2.400 359.560 17.350 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2235.230 3015.955 2235.510 3016.325 ;
        RECT 2235.300 3010.000 2235.440 3015.955 ;
        RECT 2235.300 3009.340 2235.650 3010.000 ;
        RECT 2235.370 3006.000 2235.650 3009.340 ;
        RECT 377.290 18.515 377.570 18.885 ;
        RECT 377.360 2.400 377.500 18.515 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 2235.230 3016.000 2235.510 3016.280 ;
        RECT 377.290 18.560 377.570 18.840 ;
      LAYER met3 ;
        RECT 414.270 3016.290 414.650 3016.300 ;
        RECT 2235.205 3016.290 2235.535 3016.305 ;
        RECT 414.270 3015.990 2235.535 3016.290 ;
        RECT 414.270 3015.980 414.650 3015.990 ;
        RECT 2235.205 3015.975 2235.535 3015.990 ;
        RECT 414.270 3001.330 414.650 3001.340 ;
        RECT 403.270 3001.030 414.650 3001.330 ;
        RECT 378.390 3000.650 378.770 3000.660 ;
        RECT 403.270 3000.650 403.570 3001.030 ;
        RECT 414.270 3001.020 414.650 3001.030 ;
        RECT 378.390 3000.350 403.570 3000.650 ;
        RECT 378.390 3000.340 378.770 3000.350 ;
        RECT 377.265 18.850 377.595 18.865 ;
        RECT 378.390 18.850 378.770 18.860 ;
        RECT 377.265 18.550 378.770 18.850 ;
        RECT 377.265 18.535 377.595 18.550 ;
        RECT 378.390 18.540 378.770 18.550 ;
      LAYER via3 ;
        RECT 414.300 3015.980 414.620 3016.300 ;
        RECT 378.420 3000.340 378.740 3000.660 ;
        RECT 414.300 3001.020 414.620 3001.340 ;
        RECT 378.420 18.540 378.740 18.860 ;
      LAYER met4 ;
        RECT 414.295 3015.975 414.625 3016.305 ;
        RECT 414.310 3001.345 414.610 3015.975 ;
        RECT 414.295 3001.015 414.625 3001.345 ;
        RECT 378.415 3000.335 378.745 3000.665 ;
        RECT 378.430 18.865 378.730 3000.335 ;
        RECT 378.415 18.535 378.745 18.865 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 379.185 3011.465 379.355 3029.995 ;
        RECT 489.125 3029.825 489.755 3029.995 ;
        RECT 516.725 3029.825 517.355 3029.995 ;
        RECT 614.245 3029.825 614.415 3033.395 ;
        RECT 703.485 3030.165 703.655 3033.395 ;
        RECT 752.245 3028.805 752.415 3030.335 ;
        RECT 776.165 3028.805 776.335 3030.335 ;
      LAYER mcon ;
        RECT 614.245 3033.225 614.415 3033.395 ;
        RECT 703.485 3033.225 703.655 3033.395 ;
        RECT 752.245 3030.165 752.415 3030.335 ;
        RECT 379.185 3029.825 379.355 3029.995 ;
        RECT 489.585 3029.825 489.755 3029.995 ;
        RECT 517.185 3029.825 517.355 3029.995 ;
        RECT 776.165 3030.165 776.335 3030.335 ;
      LAYER met1 ;
        RECT 614.185 3033.380 614.475 3033.425 ;
        RECT 703.425 3033.380 703.715 3033.425 ;
        RECT 614.185 3033.240 703.715 3033.380 ;
        RECT 614.185 3033.195 614.475 3033.240 ;
        RECT 703.425 3033.195 703.715 3033.240 ;
        RECT 703.425 3030.320 703.715 3030.365 ;
        RECT 752.185 3030.320 752.475 3030.365 ;
        RECT 703.425 3030.180 752.475 3030.320 ;
        RECT 703.425 3030.135 703.715 3030.180 ;
        RECT 752.185 3030.135 752.475 3030.180 ;
        RECT 776.105 3030.320 776.395 3030.365 ;
        RECT 839.570 3030.320 839.890 3030.380 ;
        RECT 776.105 3030.180 839.890 3030.320 ;
        RECT 776.105 3030.135 776.395 3030.180 ;
        RECT 839.570 3030.120 839.890 3030.180 ;
        RECT 379.125 3029.980 379.415 3030.025 ;
        RECT 489.065 3029.980 489.355 3030.025 ;
        RECT 379.125 3029.840 489.355 3029.980 ;
        RECT 379.125 3029.795 379.415 3029.840 ;
        RECT 489.065 3029.795 489.355 3029.840 ;
        RECT 489.525 3029.980 489.815 3030.025 ;
        RECT 516.665 3029.980 516.955 3030.025 ;
        RECT 489.525 3029.840 516.955 3029.980 ;
        RECT 489.525 3029.795 489.815 3029.840 ;
        RECT 516.665 3029.795 516.955 3029.840 ;
        RECT 517.125 3029.980 517.415 3030.025 ;
        RECT 614.185 3029.980 614.475 3030.025 ;
        RECT 517.125 3029.840 614.475 3029.980 ;
        RECT 517.125 3029.795 517.415 3029.840 ;
        RECT 614.185 3029.795 614.475 3029.840 ;
        RECT 752.185 3028.960 752.475 3029.005 ;
        RECT 776.105 3028.960 776.395 3029.005 ;
        RECT 752.185 3028.820 776.395 3028.960 ;
        RECT 752.185 3028.775 752.475 3028.820 ;
        RECT 776.105 3028.775 776.395 3028.820 ;
        RECT 296.310 3012.300 296.630 3012.360 ;
        RECT 296.310 3012.160 343.920 3012.300 ;
        RECT 296.310 3012.100 296.630 3012.160 ;
        RECT 343.780 3011.620 343.920 3012.160 ;
        RECT 379.125 3011.620 379.415 3011.665 ;
        RECT 343.780 3011.480 379.415 3011.620 ;
        RECT 379.125 3011.435 379.415 3011.480 ;
        RECT 296.310 465.700 296.630 465.760 ;
        RECT 393.370 465.700 393.690 465.760 ;
        RECT 296.310 465.560 393.690 465.700 ;
        RECT 296.310 465.500 296.630 465.560 ;
        RECT 393.370 465.500 393.690 465.560 ;
      LAYER via ;
        RECT 839.600 3030.120 839.860 3030.380 ;
        RECT 296.340 3012.100 296.600 3012.360 ;
        RECT 296.340 465.500 296.600 465.760 ;
        RECT 393.400 465.500 393.660 465.760 ;
      LAYER met2 ;
        RECT 839.600 3030.090 839.860 3030.410 ;
        RECT 296.340 3012.070 296.600 3012.390 ;
        RECT 296.400 465.790 296.540 3012.070 ;
        RECT 839.660 3010.000 839.800 3030.090 ;
        RECT 839.660 3009.340 840.010 3010.000 ;
        RECT 839.730 3006.000 840.010 3009.340 ;
        RECT 296.340 465.470 296.600 465.790 ;
        RECT 393.400 465.470 393.660 465.790 ;
        RECT 393.460 17.410 393.600 465.470 ;
        RECT 393.460 17.270 395.440 17.410 ;
        RECT 395.300 2.400 395.440 17.270 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 309.190 3032.360 309.510 3032.420 ;
        RECT 1123.850 3032.360 1124.170 3032.420 ;
        RECT 309.190 3032.220 1124.170 3032.360 ;
        RECT 309.190 3032.160 309.510 3032.220 ;
        RECT 1123.850 3032.160 1124.170 3032.220 ;
        RECT 309.190 487.120 309.510 487.180 ;
        RECT 409.470 487.120 409.790 487.180 ;
        RECT 309.190 486.980 409.790 487.120 ;
        RECT 309.190 486.920 309.510 486.980 ;
        RECT 409.470 486.920 409.790 486.980 ;
        RECT 409.470 16.900 409.790 16.960 ;
        RECT 413.150 16.900 413.470 16.960 ;
        RECT 409.470 16.760 413.470 16.900 ;
        RECT 409.470 16.700 409.790 16.760 ;
        RECT 413.150 16.700 413.470 16.760 ;
      LAYER via ;
        RECT 309.220 3032.160 309.480 3032.420 ;
        RECT 1123.880 3032.160 1124.140 3032.420 ;
        RECT 309.220 486.920 309.480 487.180 ;
        RECT 409.500 486.920 409.760 487.180 ;
        RECT 409.500 16.700 409.760 16.960 ;
        RECT 413.180 16.700 413.440 16.960 ;
      LAYER met2 ;
        RECT 309.220 3032.130 309.480 3032.450 ;
        RECT 1123.880 3032.130 1124.140 3032.450 ;
        RECT 309.280 487.210 309.420 3032.130 ;
        RECT 1123.940 3010.000 1124.080 3032.130 ;
        RECT 1123.940 3009.340 1124.290 3010.000 ;
        RECT 1124.010 3006.000 1124.290 3009.340 ;
        RECT 309.220 486.890 309.480 487.210 ;
        RECT 409.500 486.890 409.760 487.210 ;
        RECT 409.560 16.990 409.700 486.890 ;
        RECT 409.500 16.670 409.760 16.990 ;
        RECT 413.180 16.670 413.440 16.990 ;
        RECT 413.240 2.400 413.380 16.670 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 658.790 500.040 659.110 500.100 ;
        RECT 696.050 500.040 696.370 500.100 ;
        RECT 658.790 499.900 696.370 500.040 ;
        RECT 658.790 499.840 659.110 499.900 ;
        RECT 696.050 499.840 696.370 499.900 ;
        RECT 75.510 279.380 75.830 279.440 ;
        RECT 658.790 279.380 659.110 279.440 ;
        RECT 75.510 279.240 659.110 279.380 ;
        RECT 75.510 279.180 75.830 279.240 ;
        RECT 658.790 279.180 659.110 279.240 ;
      LAYER via ;
        RECT 658.820 499.840 659.080 500.100 ;
        RECT 696.080 499.840 696.340 500.100 ;
        RECT 75.540 279.180 75.800 279.440 ;
        RECT 658.820 279.180 659.080 279.440 ;
      LAYER met2 ;
        RECT 696.210 510.340 696.490 514.000 ;
        RECT 696.140 510.000 696.490 510.340 ;
        RECT 696.140 500.130 696.280 510.000 ;
        RECT 658.820 499.810 659.080 500.130 ;
        RECT 696.080 499.810 696.340 500.130 ;
        RECT 658.880 279.470 659.020 499.810 ;
        RECT 75.540 279.150 75.800 279.470 ;
        RECT 658.820 279.150 659.080 279.470 ;
        RECT 75.600 17.410 75.740 279.150 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 410.850 506.500 411.170 506.560 ;
        RECT 427.870 506.500 428.190 506.560 ;
        RECT 410.850 506.360 428.190 506.500 ;
        RECT 410.850 506.300 411.170 506.360 ;
        RECT 427.870 506.300 428.190 506.360 ;
      LAYER via ;
        RECT 410.880 506.300 411.140 506.560 ;
        RECT 427.900 506.300 428.160 506.560 ;
      LAYER met2 ;
        RECT 410.870 602.635 411.150 603.005 ;
        RECT 410.940 506.590 411.080 602.635 ;
        RECT 410.880 506.270 411.140 506.590 ;
        RECT 427.900 506.270 428.160 506.590 ;
        RECT 427.960 17.410 428.100 506.270 ;
        RECT 427.960 17.270 430.860 17.410 ;
        RECT 430.720 2.400 430.860 17.270 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 410.870 602.680 411.150 602.960 ;
      LAYER met3 ;
        RECT 410.000 605.240 414.000 605.840 ;
        RECT 410.630 602.985 410.930 605.240 ;
        RECT 410.630 602.670 411.175 602.985 ;
        RECT 410.845 602.655 411.175 602.670 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 454.550 237.900 454.870 237.960 ;
        RECT 1000.570 237.900 1000.890 237.960 ;
        RECT 454.550 237.760 1000.890 237.900 ;
        RECT 454.550 237.700 454.870 237.760 ;
        RECT 1000.570 237.700 1000.890 237.760 ;
        RECT 448.570 16.900 448.890 16.960 ;
        RECT 454.550 16.900 454.870 16.960 ;
        RECT 448.570 16.760 454.870 16.900 ;
        RECT 448.570 16.700 448.890 16.760 ;
        RECT 454.550 16.700 454.870 16.760 ;
      LAYER via ;
        RECT 454.580 237.700 454.840 237.960 ;
        RECT 1000.600 237.700 1000.860 237.960 ;
        RECT 448.600 16.700 448.860 16.960 ;
        RECT 454.580 16.700 454.840 16.960 ;
      LAYER met2 ;
        RECT 1005.330 510.410 1005.610 514.000 ;
        RECT 1000.660 510.270 1005.610 510.410 ;
        RECT 1000.660 237.990 1000.800 510.270 ;
        RECT 1005.330 510.000 1005.610 510.270 ;
        RECT 454.580 237.670 454.840 237.990 ;
        RECT 1000.600 237.670 1000.860 237.990 ;
        RECT 454.640 16.990 454.780 237.670 ;
        RECT 448.600 16.670 448.860 16.990 ;
        RECT 454.580 16.670 454.840 16.990 ;
        RECT 448.660 2.400 448.800 16.670 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 355.200 469.130 355.260 ;
        RECT 1828.570 355.200 1828.890 355.260 ;
        RECT 468.810 355.060 1828.890 355.200 ;
        RECT 468.810 355.000 469.130 355.060 ;
        RECT 1828.570 355.000 1828.890 355.060 ;
        RECT 466.510 16.900 466.830 16.960 ;
        RECT 468.810 16.900 469.130 16.960 ;
        RECT 466.510 16.760 469.130 16.900 ;
        RECT 466.510 16.700 466.830 16.760 ;
        RECT 468.810 16.700 469.130 16.760 ;
      LAYER via ;
        RECT 468.840 355.000 469.100 355.260 ;
        RECT 1828.600 355.000 1828.860 355.260 ;
        RECT 466.540 16.700 466.800 16.960 ;
        RECT 468.840 16.700 469.100 16.960 ;
      LAYER met2 ;
        RECT 1833.330 510.410 1833.610 514.000 ;
        RECT 1828.660 510.270 1833.610 510.410 ;
        RECT 1828.660 355.290 1828.800 510.270 ;
        RECT 1833.330 510.000 1833.610 510.270 ;
        RECT 468.840 354.970 469.100 355.290 ;
        RECT 1828.600 354.970 1828.860 355.290 ;
        RECT 468.900 16.990 469.040 354.970 ;
        RECT 466.540 16.670 466.800 16.990 ;
        RECT 468.840 16.670 469.100 16.990 ;
        RECT 466.600 2.400 466.740 16.670 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1259.090 500.380 1259.410 500.440 ;
        RECT 2030.970 500.380 2031.290 500.440 ;
        RECT 1259.090 500.240 2031.290 500.380 ;
        RECT 1259.090 500.180 1259.410 500.240 ;
        RECT 2030.970 500.180 2031.290 500.240 ;
        RECT 489.510 128.760 489.830 128.820 ;
        RECT 1259.090 128.760 1259.410 128.820 ;
        RECT 489.510 128.620 1259.410 128.760 ;
        RECT 489.510 128.560 489.830 128.620 ;
        RECT 1259.090 128.560 1259.410 128.620 ;
        RECT 484.450 16.900 484.770 16.960 ;
        RECT 489.510 16.900 489.830 16.960 ;
        RECT 484.450 16.760 489.830 16.900 ;
        RECT 484.450 16.700 484.770 16.760 ;
        RECT 489.510 16.700 489.830 16.760 ;
      LAYER via ;
        RECT 1259.120 500.180 1259.380 500.440 ;
        RECT 2031.000 500.180 2031.260 500.440 ;
        RECT 489.540 128.560 489.800 128.820 ;
        RECT 1259.120 128.560 1259.380 128.820 ;
        RECT 484.480 16.700 484.740 16.960 ;
        RECT 489.540 16.700 489.800 16.960 ;
      LAYER met2 ;
        RECT 2031.130 510.340 2031.410 514.000 ;
        RECT 2031.060 510.000 2031.410 510.340 ;
        RECT 2031.060 500.470 2031.200 510.000 ;
        RECT 1259.120 500.150 1259.380 500.470 ;
        RECT 2031.000 500.150 2031.260 500.470 ;
        RECT 1259.180 128.850 1259.320 500.150 ;
        RECT 489.540 128.530 489.800 128.850 ;
        RECT 1259.120 128.530 1259.380 128.850 ;
        RECT 489.600 16.990 489.740 128.530 ;
        RECT 484.480 16.670 484.740 16.990 ;
        RECT 489.540 16.670 489.800 16.990 ;
        RECT 484.540 2.400 484.680 16.670 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 413.685 1048.985 413.855 1053.575 ;
        RECT 413.685 861.305 413.855 867.595 ;
        RECT 414.605 723.945 414.775 789.395 ;
      LAYER mcon ;
        RECT 413.685 1053.405 413.855 1053.575 ;
        RECT 413.685 867.425 413.855 867.595 ;
        RECT 414.605 789.225 414.775 789.395 ;
      LAYER met1 ;
        RECT 413.625 1053.560 413.915 1053.605 ;
        RECT 414.530 1053.560 414.850 1053.620 ;
        RECT 413.625 1053.420 414.850 1053.560 ;
        RECT 413.625 1053.375 413.915 1053.420 ;
        RECT 414.530 1053.360 414.850 1053.420 ;
        RECT 413.625 1049.140 413.915 1049.185 ;
        RECT 414.530 1049.140 414.850 1049.200 ;
        RECT 413.625 1049.000 414.850 1049.140 ;
        RECT 413.625 1048.955 413.915 1049.000 ;
        RECT 414.530 1048.940 414.850 1049.000 ;
        RECT 414.530 914.640 414.850 914.900 ;
        RECT 414.620 913.880 414.760 914.640 ;
        RECT 414.530 913.620 414.850 913.880 ;
        RECT 413.625 867.580 413.915 867.625 ;
        RECT 414.530 867.580 414.850 867.640 ;
        RECT 413.625 867.440 414.850 867.580 ;
        RECT 413.625 867.395 413.915 867.440 ;
        RECT 414.530 867.380 414.850 867.440 ;
        RECT 413.625 861.460 413.915 861.505 ;
        RECT 414.530 861.460 414.850 861.520 ;
        RECT 413.625 861.320 414.850 861.460 ;
        RECT 413.625 861.275 413.915 861.320 ;
        RECT 414.530 861.260 414.850 861.320 ;
        RECT 414.070 789.380 414.390 789.440 ;
        RECT 414.545 789.380 414.835 789.425 ;
        RECT 414.070 789.240 414.835 789.380 ;
        RECT 414.070 789.180 414.390 789.240 ;
        RECT 414.545 789.195 414.835 789.240 ;
        RECT 414.530 724.100 414.850 724.160 ;
        RECT 414.530 723.960 415.045 724.100 ;
        RECT 414.530 723.900 414.850 723.960 ;
        RECT 417.750 500.380 418.070 500.440 ;
        RECT 497.330 500.380 497.650 500.440 ;
        RECT 417.750 500.240 497.650 500.380 ;
        RECT 417.750 500.180 418.070 500.240 ;
        RECT 497.330 500.180 497.650 500.240 ;
        RECT 497.330 2.960 497.650 3.020 ;
        RECT 502.390 2.960 502.710 3.020 ;
        RECT 497.330 2.820 502.710 2.960 ;
        RECT 497.330 2.760 497.650 2.820 ;
        RECT 502.390 2.760 502.710 2.820 ;
      LAYER via ;
        RECT 414.560 1053.360 414.820 1053.620 ;
        RECT 414.560 1048.940 414.820 1049.200 ;
        RECT 414.560 914.640 414.820 914.900 ;
        RECT 414.560 913.620 414.820 913.880 ;
        RECT 414.560 867.380 414.820 867.640 ;
        RECT 414.560 861.260 414.820 861.520 ;
        RECT 414.100 789.180 414.360 789.440 ;
        RECT 414.560 723.900 414.820 724.160 ;
        RECT 417.780 500.180 418.040 500.440 ;
        RECT 497.360 500.180 497.620 500.440 ;
        RECT 497.360 2.760 497.620 3.020 ;
        RECT 502.420 2.760 502.680 3.020 ;
      LAYER met2 ;
        RECT 413.170 2264.810 413.450 2264.925 ;
        RECT 413.170 2264.670 415.680 2264.810 ;
        RECT 413.170 2264.555 413.450 2264.670 ;
        RECT 415.540 2255.970 415.680 2264.670 ;
        RECT 414.160 2255.830 415.680 2255.970 ;
        RECT 414.160 2211.090 414.300 2255.830 ;
        RECT 414.160 2210.950 417.060 2211.090 ;
        RECT 416.920 2173.690 417.060 2210.950 ;
        RECT 416.920 2173.550 418.440 2173.690 ;
        RECT 418.300 2111.810 418.440 2173.550 ;
        RECT 417.380 2111.670 418.440 2111.810 ;
        RECT 417.380 2109.770 417.520 2111.670 ;
        RECT 417.380 2109.630 418.440 2109.770 ;
        RECT 418.300 1711.290 418.440 2109.630 ;
        RECT 415.540 1711.150 418.440 1711.290 ;
        RECT 415.540 1707.890 415.680 1711.150 ;
        RECT 415.540 1707.750 417.060 1707.890 ;
        RECT 416.920 1689.530 417.060 1707.750 ;
        RECT 416.000 1689.390 417.060 1689.530 ;
        RECT 416.000 1685.450 416.140 1689.390 ;
        RECT 416.000 1685.310 417.980 1685.450 ;
        RECT 417.840 1657.570 417.980 1685.310 ;
        RECT 417.380 1657.430 417.980 1657.570 ;
        RECT 417.380 1644.650 417.520 1657.430 ;
        RECT 417.380 1644.510 418.440 1644.650 ;
        RECT 418.300 1641.930 418.440 1644.510 ;
        RECT 417.840 1641.790 418.440 1641.930 ;
        RECT 417.840 1618.130 417.980 1641.790 ;
        RECT 417.840 1617.990 418.440 1618.130 ;
        RECT 418.300 1592.290 418.440 1617.990 ;
        RECT 417.840 1592.150 418.440 1592.290 ;
        RECT 417.840 1569.850 417.980 1592.150 ;
        RECT 417.840 1569.710 418.440 1569.850 ;
        RECT 418.300 1350.210 418.440 1569.710 ;
        RECT 416.920 1350.070 418.440 1350.210 ;
        RECT 416.920 1328.450 417.060 1350.070 ;
        RECT 416.920 1328.310 417.520 1328.450 ;
        RECT 417.380 1273.370 417.520 1328.310 ;
        RECT 417.380 1273.230 418.440 1273.370 ;
        RECT 418.300 1087.730 418.440 1273.230 ;
        RECT 414.620 1087.590 418.440 1087.730 ;
        RECT 414.620 1053.650 414.760 1087.590 ;
        RECT 414.560 1053.330 414.820 1053.650 ;
        RECT 414.560 1048.910 414.820 1049.230 ;
        RECT 414.620 1040.130 414.760 1048.910 ;
        RECT 414.620 1039.990 418.440 1040.130 ;
        RECT 418.300 934.730 418.440 1039.990 ;
        RECT 414.620 934.590 418.440 934.730 ;
        RECT 414.620 914.930 414.760 934.590 ;
        RECT 414.560 914.610 414.820 914.930 ;
        RECT 414.560 913.590 414.820 913.910 ;
        RECT 414.620 867.670 414.760 913.590 ;
        RECT 414.560 867.350 414.820 867.670 ;
        RECT 414.560 861.290 414.820 861.550 ;
        RECT 414.560 861.230 415.220 861.290 ;
        RECT 414.620 861.150 415.220 861.230 ;
        RECT 415.080 859.250 415.220 861.150 ;
        RECT 415.080 859.110 418.440 859.250 ;
        RECT 418.300 792.780 418.440 859.110 ;
        RECT 414.160 792.640 418.440 792.780 ;
        RECT 414.160 789.470 414.300 792.640 ;
        RECT 414.100 789.150 414.360 789.470 ;
        RECT 414.560 723.870 414.820 724.190 ;
        RECT 414.620 720.530 414.760 723.870 ;
        RECT 414.620 720.390 415.680 720.530 ;
        RECT 415.540 719.850 415.680 720.390 ;
        RECT 415.540 719.710 416.600 719.850 ;
        RECT 416.460 717.810 416.600 719.710 ;
        RECT 416.460 717.670 417.060 717.810 ;
        RECT 416.920 693.330 417.060 717.670 ;
        RECT 416.920 693.190 418.440 693.330 ;
        RECT 418.300 534.890 418.440 693.190 ;
        RECT 417.840 534.750 418.440 534.890 ;
        RECT 417.840 525.370 417.980 534.750 ;
        RECT 417.380 525.230 417.980 525.370 ;
        RECT 417.380 523.840 417.520 525.230 ;
        RECT 417.380 523.700 418.440 523.840 ;
        RECT 418.300 521.970 418.440 523.700 ;
        RECT 417.840 521.830 418.440 521.970 ;
        RECT 417.840 500.470 417.980 521.830 ;
        RECT 417.780 500.150 418.040 500.470 ;
        RECT 497.360 500.150 497.620 500.470 ;
        RECT 497.420 3.050 497.560 500.150 ;
        RECT 497.360 2.730 497.620 3.050 ;
        RECT 502.420 2.730 502.680 3.050 ;
        RECT 502.480 2.400 502.620 2.730 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 413.170 2264.600 413.450 2264.880 ;
      LAYER met3 ;
        RECT 410.000 2267.160 414.000 2267.760 ;
        RECT 413.390 2264.905 413.690 2267.160 ;
        RECT 413.145 2264.590 413.690 2264.905 ;
        RECT 413.145 2264.575 413.475 2264.590 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 357.950 3031.000 358.270 3031.060 ;
        RECT 999.650 3031.000 999.970 3031.060 ;
        RECT 357.950 3030.860 999.970 3031.000 ;
        RECT 357.950 3030.800 358.270 3030.860 ;
        RECT 999.650 3030.800 999.970 3030.860 ;
        RECT 357.950 508.200 358.270 508.260 ;
        RECT 518.030 508.200 518.350 508.260 ;
        RECT 357.950 508.060 518.350 508.200 ;
        RECT 357.950 508.000 358.270 508.060 ;
        RECT 518.030 508.000 518.350 508.060 ;
      LAYER via ;
        RECT 357.980 3030.800 358.240 3031.060 ;
        RECT 999.680 3030.800 999.940 3031.060 ;
        RECT 357.980 508.000 358.240 508.260 ;
        RECT 518.060 508.000 518.320 508.260 ;
      LAYER met2 ;
        RECT 357.980 3030.770 358.240 3031.090 ;
        RECT 999.680 3030.770 999.940 3031.090 ;
        RECT 358.040 508.290 358.180 3030.770 ;
        RECT 999.740 3010.000 999.880 3030.770 ;
        RECT 999.740 3009.340 1000.090 3010.000 ;
        RECT 999.810 3006.000 1000.090 3009.340 ;
        RECT 357.980 507.970 358.240 508.290 ;
        RECT 518.060 507.970 518.320 508.290 ;
        RECT 518.120 17.410 518.260 507.970 ;
        RECT 518.120 17.270 520.100 17.410 ;
        RECT 519.960 2.400 520.100 17.270 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 409.930 509.560 410.250 509.620 ;
        RECT 532.290 509.560 532.610 509.620 ;
        RECT 409.930 509.420 532.610 509.560 ;
        RECT 409.930 509.360 410.250 509.420 ;
        RECT 532.290 509.360 532.610 509.420 ;
      LAYER via ;
        RECT 409.960 509.360 410.220 509.620 ;
        RECT 532.320 509.360 532.580 509.620 ;
      LAYER met2 ;
        RECT 409.950 584.955 410.230 585.325 ;
        RECT 410.020 509.650 410.160 584.955 ;
        RECT 409.960 509.330 410.220 509.650 ;
        RECT 532.320 509.330 532.580 509.650 ;
        RECT 532.380 16.900 532.520 509.330 ;
        RECT 532.380 16.760 538.040 16.900 ;
        RECT 537.900 2.400 538.040 16.760 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 409.950 585.000 410.230 585.280 ;
      LAYER met3 ;
        RECT 410.000 586.200 414.000 586.800 ;
        RECT 409.925 585.290 410.255 585.305 ;
        RECT 410.630 585.290 410.930 586.200 ;
        RECT 409.925 584.990 410.930 585.290 ;
        RECT 409.925 584.975 410.255 584.990 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 407.170 500.040 407.490 500.100 ;
        RECT 552.070 500.040 552.390 500.100 ;
        RECT 407.170 499.900 552.390 500.040 ;
        RECT 407.170 499.840 407.490 499.900 ;
        RECT 552.070 499.840 552.390 499.900 ;
      LAYER via ;
        RECT 407.200 499.840 407.460 500.100 ;
        RECT 552.100 499.840 552.360 500.100 ;
      LAYER met2 ;
        RECT 407.190 2321.675 407.470 2322.045 ;
        RECT 407.260 500.130 407.400 2321.675 ;
        RECT 407.200 499.810 407.460 500.130 ;
        RECT 552.100 499.810 552.360 500.130 ;
        RECT 552.160 17.410 552.300 499.810 ;
        RECT 552.160 17.270 555.980 17.410 ;
        RECT 555.840 2.400 555.980 17.270 ;
        RECT 555.630 -4.800 556.190 2.400 ;
      LAYER via2 ;
        RECT 407.190 2321.720 407.470 2322.000 ;
      LAYER met3 ;
        RECT 407.165 2322.010 407.495 2322.025 ;
        RECT 410.000 2322.010 414.000 2322.160 ;
        RECT 407.165 2321.710 414.000 2322.010 ;
        RECT 407.165 2321.695 407.495 2321.710 ;
        RECT 410.000 2321.560 414.000 2321.710 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 16.900 574.010 16.960 ;
        RECT 578.750 16.900 579.070 16.960 ;
        RECT 573.690 16.760 579.070 16.900 ;
        RECT 573.690 16.700 574.010 16.760 ;
        RECT 578.750 16.700 579.070 16.760 ;
      LAYER via ;
        RECT 573.720 16.700 573.980 16.960 ;
        RECT 578.780 16.700 579.040 16.960 ;
      LAYER met2 ;
        RECT 578.770 251.075 579.050 251.445 ;
        RECT 578.840 16.990 578.980 251.075 ;
        RECT 573.720 16.670 573.980 16.990 ;
        RECT 578.780 16.670 579.040 16.990 ;
        RECT 573.780 2.400 573.920 16.670 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 578.770 251.120 579.050 251.400 ;
      LAYER met3 ;
        RECT 2506.000 2585.850 2510.000 2586.000 ;
        RECT 2512.790 2585.850 2513.170 2585.860 ;
        RECT 2506.000 2585.550 2513.170 2585.850 ;
        RECT 2506.000 2585.400 2510.000 2585.550 ;
        RECT 2512.790 2585.540 2513.170 2585.550 ;
        RECT 578.745 251.410 579.075 251.425 ;
        RECT 2512.790 251.410 2513.170 251.420 ;
        RECT 578.745 251.110 2513.170 251.410 ;
        RECT 578.745 251.095 579.075 251.110 ;
        RECT 2512.790 251.100 2513.170 251.110 ;
      LAYER via3 ;
        RECT 2512.820 2585.540 2513.140 2585.860 ;
        RECT 2512.820 251.100 2513.140 251.420 ;
      LAYER met4 ;
        RECT 2512.815 2585.535 2513.145 2585.865 ;
        RECT 2512.830 251.425 2513.130 2585.535 ;
        RECT 2512.815 251.095 2513.145 251.425 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1171.230 3006.320 1171.550 3006.580 ;
        RECT 377.730 3005.160 378.050 3005.220 ;
        RECT 1171.320 3005.160 1171.460 3006.320 ;
        RECT 377.730 3005.020 1171.460 3005.160 ;
        RECT 377.730 3004.960 378.050 3005.020 ;
        RECT 377.730 507.860 378.050 507.920 ;
        RECT 586.570 507.860 586.890 507.920 ;
        RECT 377.730 507.720 586.890 507.860 ;
        RECT 377.730 507.660 378.050 507.720 ;
        RECT 586.570 507.660 586.890 507.720 ;
        RECT 586.570 16.900 586.890 16.960 ;
        RECT 591.170 16.900 591.490 16.960 ;
        RECT 586.570 16.760 591.490 16.900 ;
        RECT 586.570 16.700 586.890 16.760 ;
        RECT 591.170 16.700 591.490 16.760 ;
      LAYER via ;
        RECT 1171.260 3006.320 1171.520 3006.580 ;
        RECT 377.760 3004.960 378.020 3005.220 ;
        RECT 377.760 507.660 378.020 507.920 ;
        RECT 586.600 507.660 586.860 507.920 ;
        RECT 586.600 16.700 586.860 16.960 ;
        RECT 591.200 16.700 591.460 16.960 ;
      LAYER met2 ;
        RECT 1172.770 3006.690 1173.050 3010.000 ;
        RECT 1171.320 3006.610 1173.050 3006.690 ;
        RECT 1171.260 3006.550 1173.050 3006.610 ;
        RECT 1171.260 3006.290 1171.520 3006.550 ;
        RECT 1172.770 3006.000 1173.050 3006.550 ;
        RECT 377.760 3004.930 378.020 3005.250 ;
        RECT 377.820 507.950 377.960 3004.930 ;
        RECT 377.760 507.630 378.020 507.950 ;
        RECT 586.600 507.630 586.860 507.950 ;
        RECT 586.660 16.990 586.800 507.630 ;
        RECT 586.600 16.670 586.860 16.990 ;
        RECT 591.200 16.670 591.460 16.990 ;
        RECT 591.260 2.400 591.400 16.670 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 127.740 103.430 127.800 ;
        RECT 455.470 127.740 455.790 127.800 ;
        RECT 103.110 127.600 455.790 127.740 ;
        RECT 103.110 127.540 103.430 127.600 ;
        RECT 455.470 127.540 455.790 127.600 ;
        RECT 97.590 17.580 97.910 17.640 ;
        RECT 103.110 17.580 103.430 17.640 ;
        RECT 97.590 17.440 103.430 17.580 ;
        RECT 97.590 17.380 97.910 17.440 ;
        RECT 103.110 17.380 103.430 17.440 ;
      LAYER via ;
        RECT 103.140 127.540 103.400 127.800 ;
        RECT 455.500 127.540 455.760 127.800 ;
        RECT 97.620 17.380 97.880 17.640 ;
        RECT 103.140 17.380 103.400 17.640 ;
      LAYER met2 ;
        RECT 461.610 510.410 461.890 514.000 ;
        RECT 455.560 510.270 461.890 510.410 ;
        RECT 455.560 127.830 455.700 510.270 ;
        RECT 461.610 510.000 461.890 510.270 ;
        RECT 103.140 127.510 103.400 127.830 ;
        RECT 455.500 127.510 455.760 127.830 ;
        RECT 103.200 17.670 103.340 127.510 ;
        RECT 97.620 17.350 97.880 17.670 ;
        RECT 103.140 17.350 103.400 17.670 ;
        RECT 97.680 2.400 97.820 17.350 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 307.350 1145.700 307.670 1145.760 ;
        RECT 393.370 1145.700 393.690 1145.760 ;
        RECT 307.350 1145.560 393.690 1145.700 ;
        RECT 307.350 1145.500 307.670 1145.560 ;
        RECT 393.370 1145.500 393.690 1145.560 ;
        RECT 307.350 48.180 307.670 48.240 ;
        RECT 609.110 48.180 609.430 48.240 ;
        RECT 307.350 48.040 609.430 48.180 ;
        RECT 307.350 47.980 307.670 48.040 ;
        RECT 609.110 47.980 609.430 48.040 ;
      LAYER via ;
        RECT 307.380 1145.500 307.640 1145.760 ;
        RECT 393.400 1145.500 393.660 1145.760 ;
        RECT 307.380 47.980 307.640 48.240 ;
        RECT 609.140 47.980 609.400 48.240 ;
      LAYER met2 ;
        RECT 393.390 1152.075 393.670 1152.445 ;
        RECT 393.460 1145.790 393.600 1152.075 ;
        RECT 307.380 1145.470 307.640 1145.790 ;
        RECT 393.400 1145.470 393.660 1145.790 ;
        RECT 307.440 48.270 307.580 1145.470 ;
        RECT 307.380 47.950 307.640 48.270 ;
        RECT 609.140 47.950 609.400 48.270 ;
        RECT 609.200 2.400 609.340 47.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 393.390 1152.120 393.670 1152.400 ;
      LAYER met3 ;
        RECT 393.365 1152.410 393.695 1152.425 ;
        RECT 410.000 1152.410 414.000 1152.560 ;
        RECT 393.365 1152.110 414.000 1152.410 ;
        RECT 393.365 1152.095 393.695 1152.110 ;
        RECT 410.000 1151.960 414.000 1152.110 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 344.610 3023.520 344.930 3023.580 ;
        RECT 505.610 3023.520 505.930 3023.580 ;
        RECT 344.610 3023.380 505.930 3023.520 ;
        RECT 344.610 3023.320 344.930 3023.380 ;
        RECT 505.610 3023.320 505.930 3023.380 ;
        RECT 344.610 33.220 344.930 33.280 ;
        RECT 627.050 33.220 627.370 33.280 ;
        RECT 344.610 33.080 627.370 33.220 ;
        RECT 344.610 33.020 344.930 33.080 ;
        RECT 627.050 33.020 627.370 33.080 ;
      LAYER via ;
        RECT 344.640 3023.320 344.900 3023.580 ;
        RECT 505.640 3023.320 505.900 3023.580 ;
        RECT 344.640 33.020 344.900 33.280 ;
        RECT 627.080 33.020 627.340 33.280 ;
      LAYER met2 ;
        RECT 344.640 3023.290 344.900 3023.610 ;
        RECT 505.640 3023.290 505.900 3023.610 ;
        RECT 344.700 33.310 344.840 3023.290 ;
        RECT 505.700 3010.000 505.840 3023.290 ;
        RECT 505.700 3009.340 506.050 3010.000 ;
        RECT 505.770 3006.000 506.050 3009.340 ;
        RECT 344.640 32.990 344.900 33.310 ;
        RECT 627.080 32.990 627.340 33.310 ;
        RECT 627.140 2.400 627.280 32.990 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.010 3006.690 1036.290 3006.805 ;
        RECT 1037.530 3006.690 1037.810 3010.000 ;
        RECT 1036.010 3006.550 1037.810 3006.690 ;
        RECT 1036.010 3006.435 1036.290 3006.550 ;
        RECT 1037.530 3006.000 1037.810 3006.550 ;
        RECT 123.370 3003.035 123.650 3003.405 ;
        RECT 123.440 17.410 123.580 3003.035 ;
        RECT 121.600 17.270 123.580 17.410 ;
        RECT 121.600 2.400 121.740 17.270 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 1036.010 3006.480 1036.290 3006.760 ;
        RECT 123.370 3003.080 123.650 3003.360 ;
      LAYER met3 ;
        RECT 1003.990 3006.770 1004.370 3006.780 ;
        RECT 1035.985 3006.770 1036.315 3006.785 ;
        RECT 1003.990 3006.470 1036.315 3006.770 ;
        RECT 1003.990 3006.460 1004.370 3006.470 ;
        RECT 1035.985 3006.455 1036.315 3006.470 ;
        RECT 123.345 3003.370 123.675 3003.385 ;
        RECT 838.390 3003.370 838.770 3003.380 ;
        RECT 123.345 3003.070 838.770 3003.370 ;
        RECT 123.345 3003.055 123.675 3003.070 ;
        RECT 838.390 3003.060 838.770 3003.070 ;
        RECT 861.390 3003.370 861.770 3003.380 ;
        RECT 1003.990 3003.370 1004.370 3003.380 ;
        RECT 861.390 3003.070 1004.370 3003.370 ;
        RECT 861.390 3003.060 861.770 3003.070 ;
        RECT 1003.990 3003.060 1004.370 3003.070 ;
        RECT 838.390 3001.330 838.770 3001.340 ;
        RECT 861.390 3001.330 861.770 3001.340 ;
        RECT 838.390 3001.030 861.770 3001.330 ;
        RECT 838.390 3001.020 838.770 3001.030 ;
        RECT 861.390 3001.020 861.770 3001.030 ;
      LAYER via3 ;
        RECT 1004.020 3006.460 1004.340 3006.780 ;
        RECT 838.420 3003.060 838.740 3003.380 ;
        RECT 861.420 3003.060 861.740 3003.380 ;
        RECT 1004.020 3003.060 1004.340 3003.380 ;
        RECT 838.420 3001.020 838.740 3001.340 ;
        RECT 861.420 3001.020 861.740 3001.340 ;
      LAYER met4 ;
        RECT 1004.015 3006.455 1004.345 3006.785 ;
        RECT 1004.030 3003.385 1004.330 3006.455 ;
        RECT 838.415 3003.055 838.745 3003.385 ;
        RECT 861.415 3003.055 861.745 3003.385 ;
        RECT 1004.015 3003.055 1004.345 3003.385 ;
        RECT 838.430 3001.345 838.730 3003.055 ;
        RECT 861.430 3001.345 861.730 3003.055 ;
        RECT 838.415 3001.015 838.745 3001.345 ;
        RECT 861.415 3001.015 861.745 3001.345 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 407.170 3019.100 407.490 3019.160 ;
        RECT 2050.290 3019.100 2050.610 3019.160 ;
        RECT 407.170 3018.960 2050.610 3019.100 ;
        RECT 407.170 3018.900 407.490 3018.960 ;
        RECT 2050.290 3018.900 2050.610 3018.960 ;
        RECT 151.410 2984.080 151.730 2984.140 ;
        RECT 407.170 2984.080 407.490 2984.140 ;
        RECT 151.410 2983.940 407.490 2984.080 ;
        RECT 151.410 2983.880 151.730 2983.940 ;
        RECT 407.170 2983.880 407.490 2983.940 ;
        RECT 145.430 17.920 145.750 17.980 ;
        RECT 151.410 17.920 151.730 17.980 ;
        RECT 145.430 17.780 151.730 17.920 ;
        RECT 145.430 17.720 145.750 17.780 ;
        RECT 151.410 17.720 151.730 17.780 ;
      LAYER via ;
        RECT 407.200 3018.900 407.460 3019.160 ;
        RECT 2050.320 3018.900 2050.580 3019.160 ;
        RECT 151.440 2983.880 151.700 2984.140 ;
        RECT 407.200 2983.880 407.460 2984.140 ;
        RECT 145.460 17.720 145.720 17.980 ;
        RECT 151.440 17.720 151.700 17.980 ;
      LAYER met2 ;
        RECT 407.200 3018.870 407.460 3019.190 ;
        RECT 2050.320 3018.870 2050.580 3019.190 ;
        RECT 407.260 2984.170 407.400 3018.870 ;
        RECT 2050.380 3010.000 2050.520 3018.870 ;
        RECT 2050.380 3009.340 2050.730 3010.000 ;
        RECT 2050.450 3006.000 2050.730 3009.340 ;
        RECT 151.440 2983.850 151.700 2984.170 ;
        RECT 407.200 2983.850 407.460 2984.170 ;
        RECT 151.500 18.010 151.640 2983.850 ;
        RECT 145.460 17.690 145.720 18.010 ;
        RECT 151.440 17.690 151.700 18.010 ;
        RECT 145.520 2.400 145.660 17.690 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1753.150 3017.995 1753.430 3018.365 ;
        RECT 1753.220 3010.000 1753.360 3017.995 ;
        RECT 1753.220 3009.340 1753.570 3010.000 ;
        RECT 1753.290 3006.000 1753.570 3009.340 ;
        RECT 165.230 120.515 165.510 120.885 ;
        RECT 165.300 17.410 165.440 120.515 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 1753.150 3018.040 1753.430 3018.320 ;
        RECT 165.230 120.560 165.510 120.840 ;
      LAYER met3 ;
        RECT 354.470 3018.330 354.850 3018.340 ;
        RECT 1753.125 3018.330 1753.455 3018.345 ;
        RECT 354.470 3018.030 1753.455 3018.330 ;
        RECT 354.470 3018.020 354.850 3018.030 ;
        RECT 1753.125 3018.015 1753.455 3018.030 ;
        RECT 165.205 120.850 165.535 120.865 ;
        RECT 354.470 120.850 354.850 120.860 ;
        RECT 165.205 120.550 354.850 120.850 ;
        RECT 165.205 120.535 165.535 120.550 ;
        RECT 354.470 120.540 354.850 120.550 ;
      LAYER via3 ;
        RECT 354.500 3018.020 354.820 3018.340 ;
        RECT 354.500 120.540 354.820 120.860 ;
      LAYER met4 ;
        RECT 354.495 3018.015 354.825 3018.345 ;
        RECT 354.510 120.865 354.810 3018.015 ;
        RECT 354.495 120.535 354.825 120.865 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 320.690 3016.720 321.010 3016.780 ;
        RECT 753.090 3016.720 753.410 3016.780 ;
        RECT 320.690 3016.580 753.410 3016.720 ;
        RECT 320.690 3016.520 321.010 3016.580 ;
        RECT 753.090 3016.520 753.410 3016.580 ;
        RECT 185.910 93.060 186.230 93.120 ;
        RECT 320.690 93.060 321.010 93.120 ;
        RECT 185.910 92.920 321.010 93.060 ;
        RECT 185.910 92.860 186.230 92.920 ;
        RECT 320.690 92.860 321.010 92.920 ;
        RECT 180.850 17.580 181.170 17.640 ;
        RECT 185.910 17.580 186.230 17.640 ;
        RECT 180.850 17.440 186.230 17.580 ;
        RECT 180.850 17.380 181.170 17.440 ;
        RECT 185.910 17.380 186.230 17.440 ;
      LAYER via ;
        RECT 320.720 3016.520 320.980 3016.780 ;
        RECT 753.120 3016.520 753.380 3016.780 ;
        RECT 185.940 92.860 186.200 93.120 ;
        RECT 320.720 92.860 320.980 93.120 ;
        RECT 180.880 17.380 181.140 17.640 ;
        RECT 185.940 17.380 186.200 17.640 ;
      LAYER met2 ;
        RECT 320.720 3016.490 320.980 3016.810 ;
        RECT 753.120 3016.490 753.380 3016.810 ;
        RECT 320.780 93.150 320.920 3016.490 ;
        RECT 753.180 3010.000 753.320 3016.490 ;
        RECT 753.180 3009.340 753.530 3010.000 ;
        RECT 753.250 3006.000 753.530 3009.340 ;
        RECT 185.940 92.830 186.200 93.150 ;
        RECT 320.720 92.830 320.980 93.150 ;
        RECT 186.000 17.670 186.140 92.830 ;
        RECT 180.880 17.350 181.140 17.670 ;
        RECT 185.940 17.350 186.200 17.670 ;
        RECT 180.940 2.400 181.080 17.350 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1638.590 501.400 1638.910 501.460 ;
        RECT 1708.970 501.400 1709.290 501.460 ;
        RECT 1638.590 501.260 1709.290 501.400 ;
        RECT 1638.590 501.200 1638.910 501.260 ;
        RECT 1708.970 501.200 1709.290 501.260 ;
        RECT 199.710 79.460 200.030 79.520 ;
        RECT 1638.590 79.460 1638.910 79.520 ;
        RECT 199.710 79.320 1638.910 79.460 ;
        RECT 199.710 79.260 200.030 79.320 ;
        RECT 1638.590 79.260 1638.910 79.320 ;
      LAYER via ;
        RECT 1638.620 501.200 1638.880 501.460 ;
        RECT 1709.000 501.200 1709.260 501.460 ;
        RECT 199.740 79.260 200.000 79.520 ;
        RECT 1638.620 79.260 1638.880 79.520 ;
      LAYER met2 ;
        RECT 1709.130 510.340 1709.410 514.000 ;
        RECT 1709.060 510.000 1709.410 510.340 ;
        RECT 1709.060 501.490 1709.200 510.000 ;
        RECT 1638.620 501.170 1638.880 501.490 ;
        RECT 1709.000 501.170 1709.260 501.490 ;
        RECT 1638.680 79.550 1638.820 501.170 ;
        RECT 199.740 79.230 200.000 79.550 ;
        RECT 1638.620 79.230 1638.880 79.550 ;
        RECT 199.800 17.410 199.940 79.230 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.490 496.980 1576.810 497.040 ;
        RECT 1585.690 496.980 1586.010 497.040 ;
        RECT 1576.490 496.840 1586.010 496.980 ;
        RECT 1576.490 496.780 1576.810 496.840 ;
        RECT 1585.690 496.780 1586.010 496.840 ;
        RECT 216.730 17.920 217.050 17.980 ;
        RECT 1576.490 17.920 1576.810 17.980 ;
        RECT 216.730 17.780 1576.810 17.920 ;
        RECT 216.730 17.720 217.050 17.780 ;
        RECT 1576.490 17.720 1576.810 17.780 ;
      LAYER via ;
        RECT 1576.520 496.780 1576.780 497.040 ;
        RECT 1585.720 496.780 1585.980 497.040 ;
        RECT 216.760 17.720 217.020 17.980 ;
        RECT 1576.520 17.720 1576.780 17.980 ;
      LAYER met2 ;
        RECT 1585.850 510.340 1586.130 514.000 ;
        RECT 1585.780 510.000 1586.130 510.340 ;
        RECT 1585.780 497.070 1585.920 510.000 ;
        RECT 1576.520 496.750 1576.780 497.070 ;
        RECT 1585.720 496.750 1585.980 497.070 ;
        RECT 1576.580 18.010 1576.720 496.750 ;
        RECT 216.760 17.690 217.020 18.010 ;
        RECT 1576.520 17.690 1576.780 18.010 ;
        RECT 216.820 2.400 216.960 17.690 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 251.690 2849.780 252.010 2849.840 ;
        RECT 393.370 2849.780 393.690 2849.840 ;
        RECT 251.690 2849.640 393.690 2849.780 ;
        RECT 251.690 2849.580 252.010 2849.640 ;
        RECT 393.370 2849.580 393.690 2849.640 ;
        RECT 234.670 27.780 234.990 27.840 ;
        RECT 251.690 27.780 252.010 27.840 ;
        RECT 234.670 27.640 252.010 27.780 ;
        RECT 234.670 27.580 234.990 27.640 ;
        RECT 251.690 27.580 252.010 27.640 ;
      LAYER via ;
        RECT 251.720 2849.580 251.980 2849.840 ;
        RECT 393.400 2849.580 393.660 2849.840 ;
        RECT 234.700 27.580 234.960 27.840 ;
        RECT 251.720 27.580 251.980 27.840 ;
      LAYER met2 ;
        RECT 393.390 2850.715 393.670 2851.085 ;
        RECT 393.460 2849.870 393.600 2850.715 ;
        RECT 251.720 2849.550 251.980 2849.870 ;
        RECT 393.400 2849.550 393.660 2849.870 ;
        RECT 251.780 27.870 251.920 2849.550 ;
        RECT 234.700 27.550 234.960 27.870 ;
        RECT 251.720 27.550 251.980 27.870 ;
        RECT 234.760 2.400 234.900 27.550 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 393.390 2850.760 393.670 2851.040 ;
      LAYER met3 ;
        RECT 393.365 2851.050 393.695 2851.065 ;
        RECT 410.000 2851.050 414.000 2851.200 ;
        RECT 393.365 2850.750 414.000 2851.050 ;
        RECT 393.365 2850.735 393.695 2850.750 ;
        RECT 410.000 2850.600 414.000 2850.750 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 99.890 2139.180 100.210 2139.240 ;
        RECT 393.370 2139.180 393.690 2139.240 ;
        RECT 99.890 2139.040 393.690 2139.180 ;
        RECT 99.890 2138.980 100.210 2139.040 ;
        RECT 393.370 2138.980 393.690 2139.040 ;
        RECT 56.190 30.840 56.510 30.900 ;
        RECT 99.890 30.840 100.210 30.900 ;
        RECT 56.190 30.700 100.210 30.840 ;
        RECT 56.190 30.640 56.510 30.700 ;
        RECT 99.890 30.640 100.210 30.700 ;
      LAYER via ;
        RECT 99.920 2138.980 100.180 2139.240 ;
        RECT 393.400 2138.980 393.660 2139.240 ;
        RECT 56.220 30.640 56.480 30.900 ;
        RECT 99.920 30.640 100.180 30.900 ;
      LAYER met2 ;
        RECT 393.390 2139.435 393.670 2139.805 ;
        RECT 393.460 2139.270 393.600 2139.435 ;
        RECT 99.920 2138.950 100.180 2139.270 ;
        RECT 393.400 2138.950 393.660 2139.270 ;
        RECT 99.980 30.930 100.120 2138.950 ;
        RECT 56.220 30.610 56.480 30.930 ;
        RECT 99.920 30.610 100.180 30.930 ;
        RECT 56.280 2.400 56.420 30.610 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 393.390 2139.480 393.670 2139.760 ;
      LAYER met3 ;
        RECT 393.365 2139.770 393.695 2139.785 ;
        RECT 410.000 2139.770 414.000 2139.920 ;
        RECT 393.365 2139.470 414.000 2139.770 ;
        RECT 393.365 2139.455 393.695 2139.470 ;
        RECT 410.000 2139.320 414.000 2139.470 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2491.910 143.635 2492.190 144.005 ;
        RECT 2491.980 105.925 2492.120 143.635 ;
        RECT 2491.910 105.555 2492.190 105.925 ;
        RECT 80.130 44.355 80.410 44.725 ;
        RECT 80.200 2.400 80.340 44.355 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 2491.910 143.680 2492.190 143.960 ;
        RECT 2491.910 105.600 2492.190 105.880 ;
        RECT 80.130 44.400 80.410 44.680 ;
      LAYER met3 ;
        RECT 2506.000 1744.920 2510.000 1745.520 ;
        RECT 2508.230 1742.660 2508.530 1744.920 ;
        RECT 2508.190 1742.340 2508.570 1742.660 ;
        RECT 2491.630 144.340 2492.010 144.660 ;
        RECT 2491.670 143.985 2491.970 144.340 ;
        RECT 2491.670 143.670 2492.215 143.985 ;
        RECT 2491.885 143.655 2492.215 143.670 ;
        RECT 2491.885 105.890 2492.215 105.905 ;
        RECT 2492.550 105.890 2492.930 105.900 ;
        RECT 2491.885 105.590 2492.930 105.890 ;
        RECT 2491.885 105.575 2492.215 105.590 ;
        RECT 2492.550 105.580 2492.930 105.590 ;
        RECT 80.105 44.690 80.435 44.705 ;
        RECT 2492.550 44.690 2492.930 44.700 ;
        RECT 80.105 44.390 2492.930 44.690 ;
        RECT 80.105 44.375 80.435 44.390 ;
        RECT 2492.550 44.380 2492.930 44.390 ;
      LAYER via3 ;
        RECT 2508.220 1742.340 2508.540 1742.660 ;
        RECT 2491.660 144.340 2491.980 144.660 ;
        RECT 2492.580 105.580 2492.900 105.900 ;
        RECT 2492.580 44.380 2492.900 44.700 ;
      LAYER met4 ;
        RECT 2508.215 1742.335 2508.545 1742.665 ;
        RECT 2508.230 1715.890 2508.530 1742.335 ;
        RECT 2493.070 1714.710 2494.250 1715.890 ;
        RECT 2507.790 1714.710 2508.970 1715.890 ;
        RECT 2493.510 1589.650 2493.810 1714.710 ;
        RECT 2492.590 1589.350 2493.810 1589.650 ;
        RECT 2492.590 1511.450 2492.890 1589.350 ;
        RECT 2492.590 1511.150 2493.810 1511.450 ;
        RECT 2493.510 1208.850 2493.810 1511.150 ;
        RECT 2493.510 1208.550 2494.730 1208.850 ;
        RECT 2494.430 1202.050 2494.730 1208.550 ;
        RECT 2493.510 1201.750 2494.730 1202.050 ;
        RECT 2493.510 1103.450 2493.810 1201.750 ;
        RECT 2493.510 1103.150 2494.730 1103.450 ;
        RECT 2494.430 1098.010 2494.730 1103.150 ;
        RECT 2493.510 1097.710 2494.730 1098.010 ;
        RECT 2493.510 831.450 2493.810 1097.710 ;
        RECT 2492.590 831.150 2493.810 831.450 ;
        RECT 2492.590 736.250 2492.890 831.150 ;
        RECT 2492.590 735.950 2493.810 736.250 ;
        RECT 2493.510 335.050 2493.810 735.950 ;
        RECT 2492.590 334.750 2493.810 335.050 ;
        RECT 2492.590 307.850 2492.890 334.750 ;
        RECT 2492.590 307.550 2493.810 307.850 ;
        RECT 2493.510 158.250 2493.810 307.550 ;
        RECT 2491.670 157.950 2493.810 158.250 ;
        RECT 2491.670 144.665 2491.970 157.950 ;
        RECT 2491.655 144.335 2491.985 144.665 ;
        RECT 2492.575 105.575 2492.905 105.905 ;
        RECT 2492.590 97.050 2492.890 105.575 ;
        RECT 2492.590 96.750 2493.810 97.050 ;
        RECT 2493.510 73.250 2493.810 96.750 ;
        RECT 2491.670 72.950 2493.810 73.250 ;
        RECT 2491.670 59.650 2491.970 72.950 ;
        RECT 2491.670 59.350 2492.890 59.650 ;
        RECT 2492.590 44.705 2492.890 59.350 ;
        RECT 2492.575 44.375 2492.905 44.705 ;
      LAYER met5 ;
        RECT 2492.860 1714.500 2509.180 1716.100 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 589.790 500.720 590.110 500.780 ;
        RECT 795.410 500.720 795.730 500.780 ;
        RECT 589.790 500.580 795.730 500.720 ;
        RECT 589.790 500.520 590.110 500.580 ;
        RECT 795.410 500.520 795.730 500.580 ;
        RECT 109.550 99.860 109.870 99.920 ;
        RECT 589.790 99.860 590.110 99.920 ;
        RECT 109.550 99.720 590.110 99.860 ;
        RECT 109.550 99.660 109.870 99.720 ;
        RECT 589.790 99.660 590.110 99.720 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 109.550 17.920 109.870 17.980 ;
        RECT 103.570 17.780 109.870 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 109.550 17.720 109.870 17.780 ;
      LAYER via ;
        RECT 589.820 500.520 590.080 500.780 ;
        RECT 795.440 500.520 795.700 500.780 ;
        RECT 109.580 99.660 109.840 99.920 ;
        RECT 589.820 99.660 590.080 99.920 ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 109.580 17.720 109.840 17.980 ;
      LAYER met2 ;
        RECT 795.570 510.340 795.850 514.000 ;
        RECT 795.500 510.000 795.850 510.340 ;
        RECT 795.500 500.810 795.640 510.000 ;
        RECT 589.820 500.490 590.080 500.810 ;
        RECT 795.440 500.490 795.700 500.810 ;
        RECT 589.880 99.950 590.020 500.490 ;
        RECT 109.580 99.630 109.840 99.950 ;
        RECT 589.820 99.630 590.080 99.950 ;
        RECT 109.640 18.010 109.780 99.630 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 109.580 17.690 109.840 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 3016.040 141.610 3016.100 ;
        RECT 1518.530 3016.040 1518.850 3016.100 ;
        RECT 141.290 3015.900 1518.850 3016.040 ;
        RECT 141.290 3015.840 141.610 3015.900 ;
        RECT 1518.530 3015.840 1518.850 3015.900 ;
        RECT 130.710 115.840 131.030 115.900 ;
        RECT 141.290 115.840 141.610 115.900 ;
        RECT 130.710 115.700 141.610 115.840 ;
        RECT 130.710 115.640 131.030 115.700 ;
        RECT 141.290 115.640 141.610 115.700 ;
        RECT 127.490 17.580 127.810 17.640 ;
        RECT 130.710 17.580 131.030 17.640 ;
        RECT 127.490 17.440 131.030 17.580 ;
        RECT 127.490 17.380 127.810 17.440 ;
        RECT 130.710 17.380 131.030 17.440 ;
      LAYER via ;
        RECT 141.320 3015.840 141.580 3016.100 ;
        RECT 1518.560 3015.840 1518.820 3016.100 ;
        RECT 130.740 115.640 131.000 115.900 ;
        RECT 141.320 115.640 141.580 115.900 ;
        RECT 127.520 17.380 127.780 17.640 ;
        RECT 130.740 17.380 131.000 17.640 ;
      LAYER met2 ;
        RECT 141.320 3015.810 141.580 3016.130 ;
        RECT 1518.560 3015.810 1518.820 3016.130 ;
        RECT 141.380 115.930 141.520 3015.810 ;
        RECT 1518.620 3010.000 1518.760 3015.810 ;
        RECT 1518.620 3009.340 1518.970 3010.000 ;
        RECT 1518.690 3006.000 1518.970 3009.340 ;
        RECT 130.740 115.610 131.000 115.930 ;
        RECT 141.320 115.610 141.580 115.930 ;
        RECT 130.800 17.670 130.940 115.610 ;
        RECT 127.520 17.350 127.780 17.670 ;
        RECT 130.740 17.350 131.000 17.670 ;
        RECT 127.580 2.400 127.720 17.350 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2520.410 1614.900 2520.730 1614.960 ;
        RECT 2560.890 1614.900 2561.210 1614.960 ;
        RECT 2520.410 1614.760 2561.210 1614.900 ;
        RECT 2520.410 1614.700 2520.730 1614.760 ;
        RECT 2560.890 1614.700 2561.210 1614.760 ;
        RECT 668.450 20.980 668.770 21.040 ;
        RECT 668.450 20.840 669.600 20.980 ;
        RECT 668.450 20.780 668.770 20.840 ;
        RECT 669.460 20.640 669.600 20.840 ;
        RECT 669.460 20.500 2543.180 20.640 ;
        RECT 2543.040 20.300 2543.180 20.500 ;
        RECT 2560.890 20.300 2561.210 20.360 ;
        RECT 2543.040 20.160 2561.210 20.300 ;
        RECT 2560.890 20.100 2561.210 20.160 ;
      LAYER via ;
        RECT 2520.440 1614.700 2520.700 1614.960 ;
        RECT 2560.920 1614.700 2561.180 1614.960 ;
        RECT 668.480 20.780 668.740 21.040 ;
        RECT 2560.920 20.100 2561.180 20.360 ;
      LAYER met2 ;
        RECT 2520.430 1617.195 2520.710 1617.565 ;
        RECT 2520.500 1614.990 2520.640 1617.195 ;
        RECT 2520.440 1614.670 2520.700 1614.990 ;
        RECT 2560.920 1614.670 2561.180 1614.990 ;
        RECT 668.480 20.750 668.740 21.070 ;
        RECT 668.540 14.125 668.680 20.750 ;
        RECT 2560.980 20.390 2561.120 1614.670 ;
        RECT 2560.920 20.070 2561.180 20.390 ;
        RECT 26.310 13.755 26.590 14.125 ;
        RECT 668.470 13.755 668.750 14.125 ;
        RECT 26.380 2.400 26.520 13.755 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 2520.430 1617.240 2520.710 1617.520 ;
        RECT 26.310 13.800 26.590 14.080 ;
        RECT 668.470 13.800 668.750 14.080 ;
      LAYER met3 ;
        RECT 2506.000 1617.530 2510.000 1617.680 ;
        RECT 2520.405 1617.530 2520.735 1617.545 ;
        RECT 2506.000 1617.230 2520.735 1617.530 ;
        RECT 2506.000 1617.080 2510.000 1617.230 ;
        RECT 2520.405 1617.215 2520.735 1617.230 ;
        RECT 26.285 14.090 26.615 14.105 ;
        RECT 668.445 14.090 668.775 14.105 ;
        RECT 26.285 13.790 668.775 14.090 ;
        RECT 26.285 13.775 26.615 13.790 ;
        RECT 668.445 13.775 668.775 13.790 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 72.290 745.520 72.610 745.580 ;
        RECT 393.370 745.520 393.690 745.580 ;
        RECT 72.290 745.380 393.690 745.520 ;
        RECT 72.290 745.320 72.610 745.380 ;
        RECT 393.370 745.320 393.690 745.380 ;
        RECT 32.270 24.040 32.590 24.100 ;
        RECT 72.290 24.040 72.610 24.100 ;
        RECT 32.270 23.900 72.610 24.040 ;
        RECT 32.270 23.840 32.590 23.900 ;
        RECT 72.290 23.840 72.610 23.900 ;
      LAYER via ;
        RECT 72.320 745.320 72.580 745.580 ;
        RECT 393.400 745.320 393.660 745.580 ;
        RECT 32.300 23.840 32.560 24.100 ;
        RECT 72.320 23.840 72.580 24.100 ;
      LAYER met2 ;
        RECT 393.390 750.875 393.670 751.245 ;
        RECT 393.460 745.610 393.600 750.875 ;
        RECT 72.320 745.290 72.580 745.610 ;
        RECT 393.400 745.290 393.660 745.610 ;
        RECT 72.380 24.130 72.520 745.290 ;
        RECT 32.300 23.810 32.560 24.130 ;
        RECT 72.320 23.810 72.580 24.130 ;
        RECT 32.360 2.400 32.500 23.810 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 393.390 750.920 393.670 751.200 ;
      LAYER met3 ;
        RECT 393.365 751.210 393.695 751.225 ;
        RECT 410.000 751.210 414.000 751.360 ;
        RECT 393.365 750.910 414.000 751.210 ;
        RECT 393.365 750.895 393.695 750.910 ;
        RECT 410.000 750.760 414.000 750.910 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 3010.000 547.020 3528.900 ;
        RECT 724.020 3010.000 727.020 3528.900 ;
        RECT 904.020 3010.000 907.020 3528.900 ;
        RECT 1084.020 3010.000 1087.020 3528.900 ;
        RECT 1264.020 3010.000 1267.020 3528.900 ;
        RECT 1444.020 3010.000 1447.020 3528.900 ;
        RECT 1624.020 3010.000 1627.020 3528.900 ;
        RECT 1804.020 3010.000 1807.020 3528.900 ;
        RECT 1984.020 3010.000 1987.020 3528.900 ;
        RECT 2164.020 3010.000 2167.020 3528.900 ;
        RECT 2344.020 3010.000 2347.020 3528.900 ;
        RECT 544.020 -9.220 547.020 510.000 ;
        RECT 724.020 -9.220 727.020 510.000 ;
        RECT 904.020 -9.220 907.020 510.000 ;
        RECT 1084.020 -9.220 1087.020 510.000 ;
        RECT 1264.020 -9.220 1267.020 510.000 ;
        RECT 1444.020 -9.220 1447.020 510.000 ;
        RECT 1624.020 -9.220 1627.020 510.000 ;
        RECT 1804.020 -9.220 1807.020 510.000 ;
        RECT 1984.020 -9.220 1987.020 510.000 ;
        RECT 2164.020 -9.220 2167.020 510.000 ;
        RECT 2344.020 -9.220 2347.020 510.000 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 3010.000 457.020 3528.900 ;
        RECT 634.020 3010.000 637.020 3528.900 ;
        RECT 814.020 3010.000 817.020 3528.900 ;
        RECT 994.020 3010.000 997.020 3528.900 ;
        RECT 1174.020 3010.000 1177.020 3528.900 ;
        RECT 1354.020 3010.000 1357.020 3528.900 ;
        RECT 1534.020 3010.000 1537.020 3528.900 ;
        RECT 1714.020 3010.000 1717.020 3528.900 ;
        RECT 1894.020 3010.000 1897.020 3528.900 ;
        RECT 2074.020 3010.000 2077.020 3528.900 ;
        RECT 2254.020 3010.000 2257.020 3528.900 ;
        RECT 2434.020 3010.000 2437.020 3528.900 ;
        RECT 454.020 -9.220 457.020 510.000 ;
        RECT 634.020 -9.220 637.020 510.000 ;
        RECT 814.020 -9.220 817.020 510.000 ;
        RECT 994.020 -9.220 997.020 510.000 ;
        RECT 1174.020 -9.220 1177.020 510.000 ;
        RECT 1354.020 -9.220 1357.020 510.000 ;
        RECT 1534.020 -9.220 1537.020 510.000 ;
        RECT 1714.020 -9.220 1717.020 510.000 ;
        RECT 1894.020 -9.220 1897.020 510.000 ;
        RECT 2074.020 -9.220 2077.020 510.000 ;
        RECT 2254.020 -9.220 2257.020 510.000 ;
        RECT 2434.020 -9.220 2437.020 510.000 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 3010.000 565.020 3538.100 ;
        RECT 742.020 3010.000 745.020 3538.100 ;
        RECT 922.020 3010.000 925.020 3538.100 ;
        RECT 1102.020 3010.000 1105.020 3538.100 ;
        RECT 1282.020 3010.000 1285.020 3538.100 ;
        RECT 1462.020 3010.000 1465.020 3538.100 ;
        RECT 1642.020 3010.000 1645.020 3538.100 ;
        RECT 1822.020 3010.000 1825.020 3538.100 ;
        RECT 2002.020 3010.000 2005.020 3538.100 ;
        RECT 2182.020 3010.000 2185.020 3538.100 ;
        RECT 2362.020 3010.000 2365.020 3538.100 ;
        RECT 562.020 -18.420 565.020 510.000 ;
        RECT 742.020 -18.420 745.020 510.000 ;
        RECT 922.020 -18.420 925.020 510.000 ;
        RECT 1102.020 -18.420 1105.020 510.000 ;
        RECT 1282.020 -18.420 1285.020 510.000 ;
        RECT 1462.020 -18.420 1465.020 510.000 ;
        RECT 1642.020 -18.420 1645.020 510.000 ;
        RECT 1822.020 -18.420 1825.020 510.000 ;
        RECT 2002.020 -18.420 2005.020 510.000 ;
        RECT 2182.020 -18.420 2185.020 510.000 ;
        RECT 2362.020 -18.420 2365.020 510.000 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 3010.000 583.020 3547.300 ;
        RECT 760.020 3010.000 763.020 3547.300 ;
        RECT 940.020 3010.000 943.020 3547.300 ;
        RECT 1120.020 3010.000 1123.020 3547.300 ;
        RECT 1300.020 3010.000 1303.020 3547.300 ;
        RECT 1480.020 3010.000 1483.020 3547.300 ;
        RECT 1660.020 3010.000 1663.020 3547.300 ;
        RECT 1840.020 3010.000 1843.020 3547.300 ;
        RECT 2020.020 3010.000 2023.020 3547.300 ;
        RECT 2200.020 3010.000 2203.020 3547.300 ;
        RECT 2380.020 3010.000 2383.020 3547.300 ;
        RECT 580.020 -27.620 583.020 510.000 ;
        RECT 760.020 -27.620 763.020 510.000 ;
        RECT 940.020 -27.620 943.020 510.000 ;
        RECT 1120.020 -27.620 1123.020 510.000 ;
        RECT 1300.020 -27.620 1303.020 510.000 ;
        RECT 1480.020 -27.620 1483.020 510.000 ;
        RECT 1660.020 -27.620 1663.020 510.000 ;
        RECT 1840.020 -27.620 1843.020 510.000 ;
        RECT 2020.020 -27.620 2023.020 510.000 ;
        RECT 2200.020 -27.620 2203.020 510.000 ;
        RECT 2380.020 -27.620 2383.020 510.000 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 3010.000 493.020 3547.300 ;
        RECT 670.020 3010.000 673.020 3547.300 ;
        RECT 850.020 3010.000 853.020 3547.300 ;
        RECT 1030.020 3010.000 1033.020 3547.300 ;
        RECT 1210.020 3010.000 1213.020 3547.300 ;
        RECT 1390.020 3010.000 1393.020 3547.300 ;
        RECT 1570.020 3010.000 1573.020 3547.300 ;
        RECT 1750.020 3010.000 1753.020 3547.300 ;
        RECT 1930.020 3010.000 1933.020 3547.300 ;
        RECT 2110.020 3010.000 2113.020 3547.300 ;
        RECT 2290.020 3010.000 2293.020 3547.300 ;
        RECT 2470.020 3010.000 2473.020 3547.300 ;
        RECT 490.020 -27.620 493.020 510.000 ;
        RECT 670.020 -27.620 673.020 510.000 ;
        RECT 850.020 -27.620 853.020 510.000 ;
        RECT 1030.020 -27.620 1033.020 510.000 ;
        RECT 1210.020 -27.620 1213.020 510.000 ;
        RECT 1390.020 -27.620 1393.020 510.000 ;
        RECT 1570.020 -27.620 1573.020 510.000 ;
        RECT 1750.020 -27.620 1753.020 510.000 ;
        RECT 1930.020 -27.620 1933.020 510.000 ;
        RECT 2110.020 -27.620 2113.020 510.000 ;
        RECT 2290.020 -27.620 2293.020 510.000 ;
        RECT 2470.020 -27.620 2473.020 510.000 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 3010.000 421.020 3556.500 ;
        RECT 598.020 3010.000 601.020 3556.500 ;
        RECT 778.020 3010.000 781.020 3556.500 ;
        RECT 958.020 3010.000 961.020 3556.500 ;
        RECT 1138.020 3010.000 1141.020 3556.500 ;
        RECT 1318.020 3010.000 1321.020 3556.500 ;
        RECT 1498.020 3010.000 1501.020 3556.500 ;
        RECT 1678.020 3010.000 1681.020 3556.500 ;
        RECT 1858.020 3010.000 1861.020 3556.500 ;
        RECT 2038.020 3010.000 2041.020 3556.500 ;
        RECT 2218.020 3010.000 2221.020 3556.500 ;
        RECT 2398.020 3010.000 2401.020 3556.500 ;
        RECT 418.020 -36.820 421.020 510.000 ;
        RECT 598.020 -36.820 601.020 510.000 ;
        RECT 778.020 -36.820 781.020 510.000 ;
        RECT 958.020 -36.820 961.020 510.000 ;
        RECT 1138.020 -36.820 1141.020 510.000 ;
        RECT 1318.020 -36.820 1321.020 510.000 ;
        RECT 1498.020 -36.820 1501.020 510.000 ;
        RECT 1678.020 -36.820 1681.020 510.000 ;
        RECT 1858.020 -36.820 1861.020 510.000 ;
        RECT 2038.020 -36.820 2041.020 510.000 ;
        RECT 2218.020 -36.820 2221.020 510.000 ;
        RECT 2398.020 -36.820 2401.020 510.000 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 3010.000 511.020 3556.500 ;
        RECT 688.020 3010.000 691.020 3556.500 ;
        RECT 868.020 3010.000 871.020 3556.500 ;
        RECT 1048.020 3010.000 1051.020 3556.500 ;
        RECT 1228.020 3010.000 1231.020 3556.500 ;
        RECT 1408.020 3010.000 1411.020 3556.500 ;
        RECT 1588.020 3010.000 1591.020 3556.500 ;
        RECT 1768.020 3010.000 1771.020 3556.500 ;
        RECT 1948.020 3010.000 1951.020 3556.500 ;
        RECT 2128.020 3010.000 2131.020 3556.500 ;
        RECT 2308.020 3010.000 2311.020 3556.500 ;
        RECT 2488.020 3010.000 2491.020 3556.500 ;
        RECT 508.020 -36.820 511.020 510.000 ;
        RECT 688.020 -36.820 691.020 510.000 ;
        RECT 868.020 -36.820 871.020 510.000 ;
        RECT 1048.020 -36.820 1051.020 510.000 ;
        RECT 1228.020 -36.820 1231.020 510.000 ;
        RECT 1408.020 -36.820 1411.020 510.000 ;
        RECT 1588.020 -36.820 1591.020 510.000 ;
        RECT 1768.020 -36.820 1771.020 510.000 ;
        RECT 1948.020 -36.820 1951.020 510.000 ;
        RECT 2128.020 -36.820 2131.020 510.000 ;
        RECT 2308.020 -36.820 2311.020 510.000 ;
        RECT 2488.020 -36.820 2491.020 510.000 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 415.520 520.795 2504.380 2998.885 ;
      LAYER met1 ;
        RECT 415.520 514.460 2507.070 2999.040 ;
      LAYER met2 ;
        RECT 418.840 3005.720 419.010 3006.010 ;
        RECT 419.850 3005.720 431.890 3006.010 ;
        RECT 432.730 3005.720 443.850 3006.010 ;
        RECT 444.690 3005.720 455.810 3006.010 ;
        RECT 456.650 3005.720 468.690 3006.010 ;
        RECT 469.530 3005.720 480.650 3006.010 ;
        RECT 481.490 3005.720 493.530 3006.010 ;
        RECT 494.370 3005.720 505.490 3006.010 ;
        RECT 506.330 3005.720 518.370 3006.010 ;
        RECT 519.210 3005.720 530.330 3006.010 ;
        RECT 531.170 3005.720 542.290 3006.010 ;
        RECT 543.130 3005.720 555.170 3006.010 ;
        RECT 556.010 3005.720 567.130 3006.010 ;
        RECT 567.970 3005.720 580.010 3006.010 ;
        RECT 580.850 3005.720 591.970 3006.010 ;
        RECT 592.810 3005.720 604.850 3006.010 ;
        RECT 605.690 3005.720 616.810 3006.010 ;
        RECT 617.650 3005.720 628.770 3006.010 ;
        RECT 629.610 3005.720 641.650 3006.010 ;
        RECT 642.490 3005.720 653.610 3006.010 ;
        RECT 654.450 3005.720 666.490 3006.010 ;
        RECT 667.330 3005.720 678.450 3006.010 ;
        RECT 679.290 3005.720 691.330 3006.010 ;
        RECT 692.170 3005.720 703.290 3006.010 ;
        RECT 704.130 3005.720 715.250 3006.010 ;
        RECT 716.090 3005.720 728.130 3006.010 ;
        RECT 728.970 3005.720 740.090 3006.010 ;
        RECT 740.930 3005.720 752.970 3006.010 ;
        RECT 753.810 3005.720 764.930 3006.010 ;
        RECT 765.770 3005.720 777.810 3006.010 ;
        RECT 778.650 3005.720 789.770 3006.010 ;
        RECT 790.610 3005.720 801.730 3006.010 ;
        RECT 802.570 3005.720 814.610 3006.010 ;
        RECT 815.450 3005.720 826.570 3006.010 ;
        RECT 827.410 3005.720 839.450 3006.010 ;
        RECT 840.290 3005.720 851.410 3006.010 ;
        RECT 852.250 3005.720 864.290 3006.010 ;
        RECT 865.130 3005.720 876.250 3006.010 ;
        RECT 877.090 3005.720 888.210 3006.010 ;
        RECT 889.050 3005.720 901.090 3006.010 ;
        RECT 901.930 3005.720 913.050 3006.010 ;
        RECT 913.890 3005.720 925.930 3006.010 ;
        RECT 926.770 3005.720 937.890 3006.010 ;
        RECT 938.730 3005.720 950.770 3006.010 ;
        RECT 951.610 3005.720 962.730 3006.010 ;
        RECT 963.570 3005.720 974.690 3006.010 ;
        RECT 975.530 3005.720 987.570 3006.010 ;
        RECT 988.410 3005.720 999.530 3006.010 ;
        RECT 1000.370 3005.720 1012.410 3006.010 ;
        RECT 1013.250 3005.720 1024.370 3006.010 ;
        RECT 1025.210 3005.720 1037.250 3006.010 ;
        RECT 1038.090 3005.720 1049.210 3006.010 ;
        RECT 1050.050 3005.720 1061.170 3006.010 ;
        RECT 1062.010 3005.720 1074.050 3006.010 ;
        RECT 1074.890 3005.720 1086.010 3006.010 ;
        RECT 1086.850 3005.720 1098.890 3006.010 ;
        RECT 1099.730 3005.720 1110.850 3006.010 ;
        RECT 1111.690 3005.720 1123.730 3006.010 ;
        RECT 1124.570 3005.720 1135.690 3006.010 ;
        RECT 1136.530 3005.720 1147.650 3006.010 ;
        RECT 1148.490 3005.720 1160.530 3006.010 ;
        RECT 1161.370 3005.720 1172.490 3006.010 ;
        RECT 1173.330 3005.720 1185.370 3006.010 ;
        RECT 1186.210 3005.720 1197.330 3006.010 ;
        RECT 1198.170 3005.720 1210.210 3006.010 ;
        RECT 1211.050 3005.720 1222.170 3006.010 ;
        RECT 1223.010 3005.720 1234.130 3006.010 ;
        RECT 1234.970 3005.720 1247.010 3006.010 ;
        RECT 1247.850 3005.720 1258.970 3006.010 ;
      LAYER met2 ;
        RECT 1259.250 3006.000 1259.530 3010.000 ;
        RECT 2012.730 3006.690 2013.010 3010.000 ;
        RECT 2014.430 3006.690 2014.710 3006.805 ;
        RECT 2012.730 3006.550 2014.710 3006.690 ;
      LAYER met2 ;
        RECT 1259.810 3005.720 1271.850 3006.010 ;
        RECT 1272.690 3005.720 1283.810 3006.010 ;
        RECT 1284.650 3005.720 1296.690 3006.010 ;
        RECT 1297.530 3005.720 1308.650 3006.010 ;
        RECT 1309.490 3005.720 1320.610 3006.010 ;
        RECT 1321.450 3005.720 1333.490 3006.010 ;
        RECT 1334.330 3005.720 1345.450 3006.010 ;
        RECT 1346.290 3005.720 1358.330 3006.010 ;
        RECT 1359.170 3005.720 1370.290 3006.010 ;
        RECT 1371.130 3005.720 1383.170 3006.010 ;
        RECT 1384.010 3005.720 1395.130 3006.010 ;
        RECT 1395.970 3005.720 1407.090 3006.010 ;
        RECT 1407.930 3005.720 1419.970 3006.010 ;
        RECT 1420.810 3005.720 1431.930 3006.010 ;
        RECT 1432.770 3005.720 1444.810 3006.010 ;
        RECT 1445.650 3005.720 1456.770 3006.010 ;
        RECT 1457.610 3005.720 1469.650 3006.010 ;
        RECT 1470.490 3005.720 1481.610 3006.010 ;
        RECT 1482.450 3005.720 1493.570 3006.010 ;
        RECT 1494.410 3005.720 1506.450 3006.010 ;
        RECT 1507.290 3005.720 1518.410 3006.010 ;
        RECT 1519.250 3005.720 1531.290 3006.010 ;
        RECT 1532.130 3005.720 1543.250 3006.010 ;
        RECT 1544.090 3005.720 1556.130 3006.010 ;
        RECT 1556.970 3005.720 1568.090 3006.010 ;
        RECT 1568.930 3005.720 1580.050 3006.010 ;
        RECT 1580.890 3005.720 1592.930 3006.010 ;
        RECT 1593.770 3005.720 1604.890 3006.010 ;
        RECT 1605.730 3005.720 1617.770 3006.010 ;
        RECT 1618.610 3005.720 1629.730 3006.010 ;
        RECT 1630.570 3005.720 1642.610 3006.010 ;
        RECT 1643.450 3005.720 1654.570 3006.010 ;
        RECT 1655.410 3005.720 1666.530 3006.010 ;
        RECT 1667.370 3005.720 1679.410 3006.010 ;
        RECT 1680.250 3005.720 1691.370 3006.010 ;
        RECT 1692.210 3005.720 1704.250 3006.010 ;
        RECT 1705.090 3005.720 1716.210 3006.010 ;
        RECT 1717.050 3005.720 1729.090 3006.010 ;
        RECT 1729.930 3005.720 1741.050 3006.010 ;
        RECT 1741.890 3005.720 1753.010 3006.010 ;
        RECT 1753.850 3005.720 1765.890 3006.010 ;
        RECT 1766.730 3005.720 1777.850 3006.010 ;
        RECT 1778.690 3005.720 1790.730 3006.010 ;
        RECT 1791.570 3005.720 1802.690 3006.010 ;
        RECT 1803.530 3005.720 1815.570 3006.010 ;
        RECT 1816.410 3005.720 1827.530 3006.010 ;
        RECT 1828.370 3005.720 1839.490 3006.010 ;
        RECT 1840.330 3005.720 1852.370 3006.010 ;
        RECT 1853.210 3005.720 1864.330 3006.010 ;
        RECT 1865.170 3005.720 1877.210 3006.010 ;
        RECT 1878.050 3005.720 1889.170 3006.010 ;
        RECT 1890.010 3005.720 1902.050 3006.010 ;
        RECT 1902.890 3005.720 1914.010 3006.010 ;
        RECT 1914.850 3005.720 1925.970 3006.010 ;
        RECT 1926.810 3005.720 1938.850 3006.010 ;
        RECT 1939.690 3005.720 1950.810 3006.010 ;
        RECT 1951.650 3005.720 1963.690 3006.010 ;
        RECT 1964.530 3005.720 1975.650 3006.010 ;
        RECT 1976.490 3005.720 1988.530 3006.010 ;
        RECT 1989.370 3005.720 2000.490 3006.010 ;
        RECT 2001.330 3005.720 2012.450 3006.010 ;
      LAYER met2 ;
        RECT 2012.730 3006.000 2013.010 3006.550 ;
        RECT 2014.430 3006.435 2014.710 3006.550 ;
      LAYER met2 ;
        RECT 2013.290 3005.720 2025.330 3006.010 ;
        RECT 2026.170 3005.720 2037.290 3006.010 ;
        RECT 2038.130 3005.720 2050.170 3006.010 ;
        RECT 2051.010 3005.720 2062.130 3006.010 ;
        RECT 2062.970 3005.720 2075.010 3006.010 ;
        RECT 2075.850 3005.720 2086.970 3006.010 ;
        RECT 2087.810 3005.720 2098.930 3006.010 ;
        RECT 2099.770 3005.720 2111.810 3006.010 ;
        RECT 2112.650 3005.720 2123.770 3006.010 ;
        RECT 2124.610 3005.720 2136.650 3006.010 ;
        RECT 2137.490 3005.720 2148.610 3006.010 ;
        RECT 2149.450 3005.720 2161.490 3006.010 ;
        RECT 2162.330 3005.720 2173.450 3006.010 ;
        RECT 2174.290 3005.720 2185.410 3006.010 ;
        RECT 2186.250 3005.720 2198.290 3006.010 ;
        RECT 2199.130 3005.720 2210.250 3006.010 ;
        RECT 2211.090 3005.720 2223.130 3006.010 ;
        RECT 2223.970 3005.720 2235.090 3006.010 ;
        RECT 2235.930 3005.720 2247.970 3006.010 ;
        RECT 2248.810 3005.720 2259.930 3006.010 ;
        RECT 2260.770 3005.720 2271.890 3006.010 ;
        RECT 2272.730 3005.720 2284.770 3006.010 ;
        RECT 2285.610 3005.720 2296.730 3006.010 ;
        RECT 2297.570 3005.720 2309.610 3006.010 ;
        RECT 2310.450 3005.720 2321.570 3006.010 ;
        RECT 2322.410 3005.720 2334.450 3006.010 ;
        RECT 2335.290 3005.720 2346.410 3006.010 ;
        RECT 2347.250 3005.720 2358.370 3006.010 ;
        RECT 2359.210 3005.720 2371.250 3006.010 ;
        RECT 2372.090 3005.720 2383.210 3006.010 ;
        RECT 2384.050 3005.720 2396.090 3006.010 ;
        RECT 2396.930 3005.720 2408.050 3006.010 ;
        RECT 2408.890 3005.720 2420.930 3006.010 ;
        RECT 2421.770 3005.720 2432.890 3006.010 ;
        RECT 2433.730 3005.720 2444.850 3006.010 ;
        RECT 2445.690 3005.720 2457.730 3006.010 ;
        RECT 2458.570 3005.720 2469.690 3006.010 ;
        RECT 2470.530 3005.720 2482.570 3006.010 ;
        RECT 2483.410 3005.720 2494.530 3006.010 ;
        RECT 2495.370 3005.720 2506.490 3006.010 ;
        RECT 418.840 514.280 2507.040 3005.720 ;
        RECT 418.840 514.000 424.530 514.280 ;
        RECT 425.370 514.000 436.490 514.280 ;
        RECT 437.330 514.000 449.370 514.280 ;
        RECT 450.210 514.000 461.330 514.280 ;
        RECT 462.170 514.000 474.210 514.280 ;
        RECT 475.050 514.000 486.170 514.280 ;
        RECT 487.010 514.000 498.130 514.280 ;
        RECT 498.970 514.000 511.010 514.280 ;
        RECT 511.850 514.000 522.970 514.280 ;
        RECT 523.810 514.000 535.850 514.280 ;
        RECT 536.690 514.000 547.810 514.280 ;
        RECT 548.650 514.000 560.690 514.280 ;
        RECT 561.530 514.000 572.650 514.280 ;
        RECT 573.490 514.000 584.610 514.280 ;
        RECT 585.450 514.000 597.490 514.280 ;
        RECT 598.330 514.000 609.450 514.280 ;
        RECT 610.290 514.000 622.330 514.280 ;
        RECT 623.170 514.000 634.290 514.280 ;
        RECT 635.130 514.000 647.170 514.280 ;
        RECT 648.010 514.000 659.130 514.280 ;
        RECT 659.970 514.000 671.090 514.280 ;
        RECT 671.930 514.000 683.970 514.280 ;
        RECT 684.810 514.000 695.930 514.280 ;
        RECT 696.770 514.000 708.810 514.280 ;
        RECT 709.650 514.000 720.770 514.280 ;
        RECT 721.610 514.000 733.650 514.280 ;
        RECT 734.490 514.000 745.610 514.280 ;
        RECT 746.450 514.000 757.570 514.280 ;
        RECT 758.410 514.000 770.450 514.280 ;
        RECT 771.290 514.000 782.410 514.280 ;
        RECT 783.250 514.000 795.290 514.280 ;
        RECT 796.130 514.000 807.250 514.280 ;
        RECT 808.090 514.000 820.130 514.280 ;
        RECT 820.970 514.000 832.090 514.280 ;
        RECT 832.930 514.000 844.050 514.280 ;
        RECT 844.890 514.000 856.930 514.280 ;
        RECT 857.770 514.000 868.890 514.280 ;
        RECT 869.730 514.000 881.770 514.280 ;
        RECT 882.610 514.000 893.730 514.280 ;
        RECT 894.570 514.000 906.610 514.280 ;
        RECT 907.450 514.000 918.570 514.280 ;
        RECT 919.410 514.000 930.530 514.280 ;
        RECT 931.370 514.000 943.410 514.280 ;
        RECT 944.250 514.000 955.370 514.280 ;
        RECT 956.210 514.000 968.250 514.280 ;
        RECT 969.090 514.000 980.210 514.280 ;
        RECT 981.050 514.000 993.090 514.280 ;
        RECT 993.930 514.000 1005.050 514.280 ;
        RECT 1005.890 514.000 1017.010 514.280 ;
        RECT 1017.850 514.000 1029.890 514.280 ;
        RECT 1030.730 514.000 1041.850 514.280 ;
        RECT 1042.690 514.000 1054.730 514.280 ;
        RECT 1055.570 514.000 1066.690 514.280 ;
        RECT 1067.530 514.000 1079.570 514.280 ;
        RECT 1080.410 514.000 1091.530 514.280 ;
        RECT 1092.370 514.000 1103.490 514.280 ;
        RECT 1104.330 514.000 1116.370 514.280 ;
        RECT 1117.210 514.000 1128.330 514.280 ;
        RECT 1129.170 514.000 1141.210 514.280 ;
        RECT 1142.050 514.000 1153.170 514.280 ;
        RECT 1154.010 514.000 1166.050 514.280 ;
        RECT 1166.890 514.000 1178.010 514.280 ;
        RECT 1178.850 514.000 1189.970 514.280 ;
        RECT 1190.810 514.000 1202.850 514.280 ;
        RECT 1203.690 514.000 1214.810 514.280 ;
        RECT 1215.650 514.000 1227.690 514.280 ;
        RECT 1228.530 514.000 1239.650 514.280 ;
        RECT 1240.490 514.000 1252.530 514.280 ;
        RECT 1253.370 514.000 1264.490 514.280 ;
        RECT 1265.330 514.000 1276.450 514.280 ;
        RECT 1277.290 514.000 1289.330 514.280 ;
        RECT 1290.170 514.000 1301.290 514.280 ;
        RECT 1302.130 514.000 1314.170 514.280 ;
        RECT 1315.010 514.000 1326.130 514.280 ;
        RECT 1326.970 514.000 1339.010 514.280 ;
        RECT 1339.850 514.000 1350.970 514.280 ;
        RECT 1351.810 514.000 1362.930 514.280 ;
        RECT 1363.770 514.000 1375.810 514.280 ;
        RECT 1376.650 514.000 1387.770 514.280 ;
        RECT 1388.610 514.000 1400.650 514.280 ;
        RECT 1401.490 514.000 1412.610 514.280 ;
        RECT 1413.450 514.000 1425.490 514.280 ;
        RECT 1426.330 514.000 1437.450 514.280 ;
        RECT 1438.290 514.000 1449.410 514.280 ;
        RECT 1450.250 514.000 1462.290 514.280 ;
        RECT 1463.130 514.000 1474.250 514.280 ;
        RECT 1475.090 514.000 1487.130 514.280 ;
        RECT 1487.970 514.000 1499.090 514.280 ;
        RECT 1499.930 514.000 1511.970 514.280 ;
        RECT 1512.810 514.000 1523.930 514.280 ;
        RECT 1524.770 514.000 1535.890 514.280 ;
        RECT 1536.730 514.000 1548.770 514.280 ;
        RECT 1549.610 514.000 1560.730 514.280 ;
        RECT 1561.570 514.000 1573.610 514.280 ;
        RECT 1574.450 514.000 1585.570 514.280 ;
        RECT 1586.410 514.000 1598.450 514.280 ;
        RECT 1599.290 514.000 1610.410 514.280 ;
        RECT 1611.250 514.000 1622.370 514.280 ;
        RECT 1623.210 514.000 1635.250 514.280 ;
        RECT 1636.090 514.000 1647.210 514.280 ;
        RECT 1648.050 514.000 1660.090 514.280 ;
        RECT 1660.930 514.000 1672.050 514.280 ;
        RECT 1672.890 514.000 1684.930 514.280 ;
        RECT 1685.770 514.000 1696.890 514.280 ;
        RECT 1697.730 514.000 1708.850 514.280 ;
        RECT 1709.690 514.000 1721.730 514.280 ;
        RECT 1722.570 514.000 1733.690 514.280 ;
        RECT 1734.530 514.000 1746.570 514.280 ;
        RECT 1747.410 514.000 1758.530 514.280 ;
        RECT 1759.370 514.000 1771.410 514.280 ;
        RECT 1772.250 514.000 1783.370 514.280 ;
        RECT 1784.210 514.000 1795.330 514.280 ;
        RECT 1796.170 514.000 1808.210 514.280 ;
        RECT 1809.050 514.000 1820.170 514.280 ;
        RECT 1821.010 514.000 1833.050 514.280 ;
        RECT 1833.890 514.000 1845.010 514.280 ;
        RECT 1845.850 514.000 1857.890 514.280 ;
        RECT 1858.730 514.000 1869.850 514.280 ;
        RECT 1870.690 514.000 1881.810 514.280 ;
        RECT 1882.650 514.000 1894.690 514.280 ;
        RECT 1895.530 514.000 1906.650 514.280 ;
        RECT 1907.490 514.000 1919.530 514.280 ;
        RECT 1920.370 514.000 1931.490 514.280 ;
        RECT 1932.330 514.000 1944.370 514.280 ;
        RECT 1945.210 514.000 1956.330 514.280 ;
        RECT 1957.170 514.000 1968.290 514.280 ;
        RECT 1969.130 514.000 1981.170 514.280 ;
        RECT 1982.010 514.000 1993.130 514.280 ;
        RECT 1993.970 514.000 2006.010 514.280 ;
        RECT 2006.850 514.000 2017.970 514.280 ;
        RECT 2018.810 514.000 2030.850 514.280 ;
        RECT 2031.690 514.000 2042.810 514.280 ;
        RECT 2043.650 514.000 2054.770 514.280 ;
        RECT 2055.610 514.000 2067.650 514.280 ;
        RECT 2068.490 514.000 2079.610 514.280 ;
        RECT 2080.450 514.000 2092.490 514.280 ;
        RECT 2093.330 514.000 2104.450 514.280 ;
        RECT 2105.290 514.000 2117.330 514.280 ;
        RECT 2118.170 514.000 2129.290 514.280 ;
        RECT 2130.130 514.000 2141.250 514.280 ;
        RECT 2142.090 514.000 2154.130 514.280 ;
        RECT 2154.970 514.000 2166.090 514.280 ;
        RECT 2166.930 514.000 2178.970 514.280 ;
        RECT 2179.810 514.000 2190.930 514.280 ;
        RECT 2191.770 514.000 2203.810 514.280 ;
        RECT 2204.650 514.000 2215.770 514.280 ;
        RECT 2216.610 514.000 2227.730 514.280 ;
        RECT 2228.570 514.000 2240.610 514.280 ;
        RECT 2241.450 514.000 2252.570 514.280 ;
        RECT 2253.410 514.000 2265.450 514.280 ;
        RECT 2266.290 514.000 2277.410 514.280 ;
        RECT 2278.250 514.000 2290.290 514.280 ;
        RECT 2291.130 514.000 2302.250 514.280 ;
        RECT 2303.090 514.000 2314.210 514.280 ;
        RECT 2315.050 514.000 2327.090 514.280 ;
        RECT 2327.930 514.000 2339.050 514.280 ;
        RECT 2339.890 514.000 2351.930 514.280 ;
        RECT 2352.770 514.000 2363.890 514.280 ;
        RECT 2364.730 514.000 2376.770 514.280 ;
        RECT 2377.610 514.000 2388.730 514.280 ;
        RECT 2389.570 514.000 2400.690 514.280 ;
        RECT 2401.530 514.000 2413.570 514.280 ;
        RECT 2414.410 514.000 2425.530 514.280 ;
        RECT 2426.370 514.000 2438.410 514.280 ;
        RECT 2439.250 514.000 2450.370 514.280 ;
        RECT 2451.210 514.000 2463.250 514.280 ;
        RECT 2464.090 514.000 2475.210 514.280 ;
        RECT 2476.050 514.000 2487.170 514.280 ;
        RECT 2488.010 514.000 2500.050 514.280 ;
        RECT 2500.890 514.000 2507.040 514.280 ;
      LAYER met2 ;
        RECT 906.890 510.000 907.170 514.000 ;
        RECT 1215.090 510.000 1215.370 514.000 ;
        RECT 1660.370 510.000 1660.650 514.000 ;
        RECT 1746.850 510.000 1747.130 514.000 ;
      LAYER via2 ;
        RECT 2014.430 3006.480 2014.710 3006.760 ;
      LAYER met3 ;
        RECT 2014.405 3006.770 2014.735 3006.785 ;
        RECT 2025.190 3006.770 2025.570 3006.780 ;
        RECT 2014.405 3006.470 2025.570 3006.770 ;
        RECT 2014.405 3006.455 2014.735 3006.470 ;
        RECT 2025.190 3006.460 2025.570 3006.470 ;
        RECT 2025.190 2999.660 2025.570 2999.980 ;
        RECT 2025.230 2998.965 2025.530 2999.660 ;
      LAYER met3 ;
        RECT 414.000 2998.480 2506.000 2998.965 ;
        RECT 414.400 2997.080 2506.000 2998.480 ;
        RECT 414.000 2987.600 2506.000 2997.080 ;
        RECT 414.000 2986.200 2505.600 2987.600 ;
        RECT 414.000 2979.440 2506.000 2986.200 ;
        RECT 414.400 2978.040 2506.000 2979.440 ;
        RECT 414.000 2969.920 2506.000 2978.040 ;
        RECT 414.000 2968.520 2505.600 2969.920 ;
        RECT 414.000 2961.760 2506.000 2968.520 ;
        RECT 414.400 2960.360 2506.000 2961.760 ;
        RECT 414.000 2950.880 2506.000 2960.360 ;
        RECT 414.000 2949.480 2505.600 2950.880 ;
        RECT 414.000 2942.720 2506.000 2949.480 ;
        RECT 414.400 2941.320 2506.000 2942.720 ;
        RECT 414.000 2933.200 2506.000 2941.320 ;
        RECT 414.000 2931.800 2505.600 2933.200 ;
        RECT 414.000 2925.040 2506.000 2931.800 ;
      LAYER met3 ;
        RECT 410.000 2924.040 414.000 2924.640 ;
      LAYER met3 ;
        RECT 414.400 2923.640 2506.000 2925.040 ;
        RECT 414.000 2914.160 2506.000 2923.640 ;
        RECT 414.000 2912.760 2505.600 2914.160 ;
        RECT 414.000 2907.360 2506.000 2912.760 ;
        RECT 414.400 2905.960 2506.000 2907.360 ;
        RECT 414.000 2896.480 2506.000 2905.960 ;
        RECT 414.000 2895.080 2505.600 2896.480 ;
        RECT 414.000 2888.320 2506.000 2895.080 ;
        RECT 414.400 2886.920 2506.000 2888.320 ;
        RECT 414.000 2878.800 2506.000 2886.920 ;
        RECT 414.000 2877.400 2505.600 2878.800 ;
        RECT 414.000 2870.640 2506.000 2877.400 ;
        RECT 414.400 2869.240 2506.000 2870.640 ;
        RECT 414.000 2859.760 2506.000 2869.240 ;
        RECT 414.000 2858.360 2505.600 2859.760 ;
        RECT 414.000 2851.600 2506.000 2858.360 ;
        RECT 414.400 2850.200 2506.000 2851.600 ;
        RECT 414.000 2842.080 2506.000 2850.200 ;
        RECT 414.000 2840.680 2505.600 2842.080 ;
        RECT 414.000 2833.920 2506.000 2840.680 ;
        RECT 414.400 2832.520 2506.000 2833.920 ;
        RECT 414.000 2823.040 2506.000 2832.520 ;
        RECT 414.000 2821.640 2505.600 2823.040 ;
        RECT 414.000 2814.880 2506.000 2821.640 ;
        RECT 414.400 2813.480 2506.000 2814.880 ;
        RECT 414.000 2805.360 2506.000 2813.480 ;
        RECT 414.000 2803.960 2505.600 2805.360 ;
        RECT 414.000 2797.200 2506.000 2803.960 ;
        RECT 414.400 2795.800 2506.000 2797.200 ;
        RECT 414.000 2786.320 2506.000 2795.800 ;
        RECT 414.000 2784.920 2505.600 2786.320 ;
        RECT 414.000 2779.520 2506.000 2784.920 ;
        RECT 414.400 2778.120 2506.000 2779.520 ;
        RECT 414.000 2768.640 2506.000 2778.120 ;
        RECT 414.000 2767.240 2505.600 2768.640 ;
        RECT 414.000 2760.480 2506.000 2767.240 ;
        RECT 414.400 2759.080 2506.000 2760.480 ;
        RECT 414.000 2750.960 2506.000 2759.080 ;
        RECT 414.000 2749.560 2505.600 2750.960 ;
        RECT 414.000 2742.800 2506.000 2749.560 ;
        RECT 414.400 2741.400 2506.000 2742.800 ;
        RECT 414.000 2731.920 2506.000 2741.400 ;
        RECT 414.000 2730.520 2505.600 2731.920 ;
        RECT 414.000 2723.760 2506.000 2730.520 ;
        RECT 414.400 2722.360 2506.000 2723.760 ;
        RECT 414.000 2714.240 2506.000 2722.360 ;
        RECT 414.000 2712.840 2505.600 2714.240 ;
        RECT 414.000 2706.080 2506.000 2712.840 ;
        RECT 414.400 2704.680 2506.000 2706.080 ;
        RECT 414.000 2695.200 2506.000 2704.680 ;
        RECT 414.000 2693.800 2505.600 2695.200 ;
        RECT 414.000 2687.040 2506.000 2693.800 ;
        RECT 414.400 2685.640 2506.000 2687.040 ;
        RECT 414.000 2677.520 2506.000 2685.640 ;
        RECT 414.000 2676.120 2505.600 2677.520 ;
        RECT 414.000 2669.360 2506.000 2676.120 ;
        RECT 414.400 2667.960 2506.000 2669.360 ;
        RECT 414.000 2658.480 2506.000 2667.960 ;
        RECT 414.000 2657.080 2505.600 2658.480 ;
        RECT 414.000 2651.680 2506.000 2657.080 ;
        RECT 414.400 2650.280 2506.000 2651.680 ;
        RECT 414.000 2640.800 2506.000 2650.280 ;
        RECT 414.000 2639.400 2505.600 2640.800 ;
      LAYER met3 ;
        RECT 2506.000 2639.800 2510.000 2640.400 ;
      LAYER met3 ;
        RECT 414.000 2632.640 2506.000 2639.400 ;
        RECT 414.400 2631.240 2506.000 2632.640 ;
        RECT 414.000 2623.120 2506.000 2631.240 ;
        RECT 414.000 2621.720 2505.600 2623.120 ;
        RECT 414.000 2614.960 2506.000 2621.720 ;
        RECT 414.400 2613.560 2506.000 2614.960 ;
        RECT 414.000 2604.080 2506.000 2613.560 ;
        RECT 414.000 2602.680 2505.600 2604.080 ;
        RECT 414.000 2595.920 2506.000 2602.680 ;
        RECT 414.400 2594.520 2506.000 2595.920 ;
        RECT 414.000 2586.400 2506.000 2594.520 ;
        RECT 414.000 2585.000 2505.600 2586.400 ;
        RECT 414.000 2578.240 2506.000 2585.000 ;
        RECT 414.400 2576.840 2506.000 2578.240 ;
        RECT 414.000 2567.360 2506.000 2576.840 ;
        RECT 414.000 2565.960 2505.600 2567.360 ;
        RECT 414.000 2559.200 2506.000 2565.960 ;
        RECT 414.400 2557.800 2506.000 2559.200 ;
        RECT 414.000 2549.680 2506.000 2557.800 ;
        RECT 414.000 2548.280 2505.600 2549.680 ;
        RECT 414.000 2541.520 2506.000 2548.280 ;
        RECT 414.400 2540.120 2506.000 2541.520 ;
        RECT 414.000 2530.640 2506.000 2540.120 ;
        RECT 414.000 2529.240 2505.600 2530.640 ;
        RECT 414.000 2523.840 2506.000 2529.240 ;
        RECT 414.400 2522.440 2506.000 2523.840 ;
        RECT 414.000 2512.960 2506.000 2522.440 ;
        RECT 414.000 2511.560 2505.600 2512.960 ;
        RECT 414.000 2504.800 2506.000 2511.560 ;
        RECT 414.400 2503.400 2506.000 2504.800 ;
        RECT 414.000 2495.280 2506.000 2503.400 ;
        RECT 414.000 2493.880 2505.600 2495.280 ;
        RECT 414.000 2487.120 2506.000 2493.880 ;
        RECT 414.400 2485.720 2506.000 2487.120 ;
        RECT 414.000 2476.240 2506.000 2485.720 ;
        RECT 414.000 2474.840 2505.600 2476.240 ;
        RECT 414.000 2468.080 2506.000 2474.840 ;
        RECT 414.400 2466.680 2506.000 2468.080 ;
        RECT 414.000 2458.560 2506.000 2466.680 ;
        RECT 414.000 2457.160 2505.600 2458.560 ;
        RECT 414.000 2450.400 2506.000 2457.160 ;
        RECT 414.400 2449.000 2506.000 2450.400 ;
        RECT 414.000 2439.520 2506.000 2449.000 ;
        RECT 414.000 2438.120 2505.600 2439.520 ;
        RECT 414.000 2431.360 2506.000 2438.120 ;
        RECT 414.400 2429.960 2506.000 2431.360 ;
        RECT 414.000 2421.840 2506.000 2429.960 ;
        RECT 414.000 2420.440 2505.600 2421.840 ;
        RECT 414.000 2413.680 2506.000 2420.440 ;
        RECT 414.400 2412.280 2506.000 2413.680 ;
        RECT 414.000 2402.800 2506.000 2412.280 ;
        RECT 414.000 2401.400 2505.600 2402.800 ;
        RECT 414.000 2396.000 2506.000 2401.400 ;
        RECT 414.400 2394.600 2506.000 2396.000 ;
        RECT 414.000 2385.120 2506.000 2394.600 ;
        RECT 414.000 2383.720 2505.600 2385.120 ;
        RECT 414.000 2376.960 2506.000 2383.720 ;
        RECT 414.400 2375.560 2506.000 2376.960 ;
        RECT 414.000 2367.440 2506.000 2375.560 ;
        RECT 414.000 2366.040 2505.600 2367.440 ;
        RECT 414.000 2359.280 2506.000 2366.040 ;
        RECT 414.400 2357.880 2506.000 2359.280 ;
        RECT 414.000 2348.400 2506.000 2357.880 ;
        RECT 414.000 2347.000 2505.600 2348.400 ;
        RECT 414.000 2340.240 2506.000 2347.000 ;
        RECT 414.400 2338.840 2506.000 2340.240 ;
        RECT 414.000 2330.720 2506.000 2338.840 ;
        RECT 414.000 2329.320 2505.600 2330.720 ;
        RECT 414.000 2322.560 2506.000 2329.320 ;
        RECT 414.400 2321.160 2506.000 2322.560 ;
        RECT 414.000 2311.680 2506.000 2321.160 ;
        RECT 414.000 2310.280 2505.600 2311.680 ;
        RECT 414.000 2303.520 2506.000 2310.280 ;
        RECT 414.400 2302.120 2506.000 2303.520 ;
        RECT 414.000 2294.000 2506.000 2302.120 ;
        RECT 414.000 2292.600 2505.600 2294.000 ;
        RECT 414.000 2285.840 2506.000 2292.600 ;
        RECT 414.400 2284.440 2506.000 2285.840 ;
        RECT 414.000 2274.960 2506.000 2284.440 ;
        RECT 414.000 2273.560 2505.600 2274.960 ;
        RECT 414.000 2268.160 2506.000 2273.560 ;
        RECT 414.400 2266.760 2506.000 2268.160 ;
        RECT 414.000 2257.280 2506.000 2266.760 ;
        RECT 414.000 2255.880 2505.600 2257.280 ;
        RECT 414.000 2249.120 2506.000 2255.880 ;
        RECT 414.400 2247.720 2506.000 2249.120 ;
        RECT 414.000 2239.600 2506.000 2247.720 ;
        RECT 414.000 2238.200 2505.600 2239.600 ;
        RECT 414.000 2231.440 2506.000 2238.200 ;
        RECT 414.400 2230.040 2506.000 2231.440 ;
        RECT 414.000 2220.560 2506.000 2230.040 ;
        RECT 414.000 2219.160 2505.600 2220.560 ;
        RECT 414.000 2212.400 2506.000 2219.160 ;
        RECT 414.400 2211.000 2506.000 2212.400 ;
        RECT 414.000 2202.880 2506.000 2211.000 ;
        RECT 414.000 2201.480 2505.600 2202.880 ;
        RECT 414.000 2194.720 2506.000 2201.480 ;
        RECT 414.400 2193.320 2506.000 2194.720 ;
        RECT 414.000 2183.840 2506.000 2193.320 ;
        RECT 414.000 2182.440 2505.600 2183.840 ;
        RECT 414.000 2175.680 2506.000 2182.440 ;
        RECT 414.400 2174.280 2506.000 2175.680 ;
        RECT 414.000 2166.160 2506.000 2174.280 ;
        RECT 414.000 2164.760 2505.600 2166.160 ;
        RECT 414.000 2158.000 2506.000 2164.760 ;
        RECT 414.400 2156.600 2506.000 2158.000 ;
        RECT 414.000 2147.120 2506.000 2156.600 ;
        RECT 414.000 2145.720 2505.600 2147.120 ;
        RECT 414.000 2140.320 2506.000 2145.720 ;
        RECT 414.400 2138.920 2506.000 2140.320 ;
        RECT 414.000 2129.440 2506.000 2138.920 ;
        RECT 414.000 2128.040 2505.600 2129.440 ;
        RECT 414.000 2121.280 2506.000 2128.040 ;
        RECT 414.400 2119.880 2506.000 2121.280 ;
        RECT 414.000 2111.760 2506.000 2119.880 ;
        RECT 414.000 2110.360 2505.600 2111.760 ;
        RECT 414.000 2103.600 2506.000 2110.360 ;
        RECT 414.400 2102.200 2506.000 2103.600 ;
        RECT 414.000 2092.720 2506.000 2102.200 ;
        RECT 414.000 2091.320 2505.600 2092.720 ;
        RECT 414.000 2084.560 2506.000 2091.320 ;
        RECT 414.400 2083.160 2506.000 2084.560 ;
        RECT 414.000 2075.040 2506.000 2083.160 ;
        RECT 414.000 2073.640 2505.600 2075.040 ;
        RECT 414.000 2066.880 2506.000 2073.640 ;
        RECT 414.400 2065.480 2506.000 2066.880 ;
        RECT 414.000 2056.000 2506.000 2065.480 ;
        RECT 414.000 2054.600 2505.600 2056.000 ;
        RECT 414.000 2047.840 2506.000 2054.600 ;
        RECT 414.400 2046.440 2506.000 2047.840 ;
        RECT 414.000 2038.320 2506.000 2046.440 ;
        RECT 414.000 2036.920 2505.600 2038.320 ;
        RECT 414.000 2030.160 2506.000 2036.920 ;
        RECT 414.400 2028.760 2506.000 2030.160 ;
        RECT 414.000 2019.280 2506.000 2028.760 ;
        RECT 414.000 2017.880 2505.600 2019.280 ;
        RECT 414.000 2012.480 2506.000 2017.880 ;
        RECT 414.400 2011.080 2506.000 2012.480 ;
        RECT 414.000 2001.600 2506.000 2011.080 ;
        RECT 414.000 2000.200 2505.600 2001.600 ;
        RECT 414.000 1993.440 2506.000 2000.200 ;
        RECT 414.400 1992.040 2506.000 1993.440 ;
        RECT 414.000 1983.920 2506.000 1992.040 ;
        RECT 414.000 1982.520 2505.600 1983.920 ;
        RECT 414.000 1975.760 2506.000 1982.520 ;
        RECT 414.400 1974.360 2506.000 1975.760 ;
        RECT 414.000 1964.880 2506.000 1974.360 ;
        RECT 414.000 1963.480 2505.600 1964.880 ;
        RECT 414.000 1956.720 2506.000 1963.480 ;
        RECT 414.400 1955.320 2506.000 1956.720 ;
        RECT 414.000 1947.200 2506.000 1955.320 ;
        RECT 414.000 1945.800 2505.600 1947.200 ;
        RECT 414.000 1939.040 2506.000 1945.800 ;
        RECT 414.400 1937.640 2506.000 1939.040 ;
        RECT 414.000 1928.160 2506.000 1937.640 ;
        RECT 414.000 1926.760 2505.600 1928.160 ;
        RECT 414.000 1920.000 2506.000 1926.760 ;
        RECT 414.400 1918.600 2506.000 1920.000 ;
        RECT 414.000 1910.480 2506.000 1918.600 ;
        RECT 414.000 1909.080 2505.600 1910.480 ;
        RECT 414.000 1902.320 2506.000 1909.080 ;
        RECT 414.400 1900.920 2506.000 1902.320 ;
        RECT 414.000 1891.440 2506.000 1900.920 ;
        RECT 414.000 1890.040 2505.600 1891.440 ;
        RECT 414.000 1884.640 2506.000 1890.040 ;
        RECT 414.400 1883.240 2506.000 1884.640 ;
        RECT 414.000 1873.760 2506.000 1883.240 ;
        RECT 414.000 1872.360 2505.600 1873.760 ;
        RECT 414.000 1865.600 2506.000 1872.360 ;
        RECT 414.400 1864.200 2506.000 1865.600 ;
        RECT 414.000 1856.080 2506.000 1864.200 ;
        RECT 414.000 1854.680 2505.600 1856.080 ;
        RECT 414.000 1847.920 2506.000 1854.680 ;
        RECT 414.400 1846.520 2506.000 1847.920 ;
        RECT 414.000 1837.040 2506.000 1846.520 ;
        RECT 414.000 1835.640 2505.600 1837.040 ;
        RECT 414.000 1828.880 2506.000 1835.640 ;
        RECT 414.400 1827.480 2506.000 1828.880 ;
        RECT 414.000 1819.360 2506.000 1827.480 ;
        RECT 414.000 1817.960 2505.600 1819.360 ;
        RECT 414.000 1811.200 2506.000 1817.960 ;
        RECT 414.400 1809.800 2506.000 1811.200 ;
        RECT 414.000 1800.320 2506.000 1809.800 ;
        RECT 414.000 1798.920 2505.600 1800.320 ;
        RECT 414.000 1792.160 2506.000 1798.920 ;
        RECT 414.400 1790.760 2506.000 1792.160 ;
        RECT 414.000 1782.640 2506.000 1790.760 ;
        RECT 414.000 1781.240 2505.600 1782.640 ;
        RECT 414.000 1774.480 2506.000 1781.240 ;
      LAYER met3 ;
        RECT 410.000 1773.480 414.000 1774.080 ;
      LAYER met3 ;
        RECT 414.400 1773.080 2506.000 1774.480 ;
        RECT 414.000 1763.600 2506.000 1773.080 ;
        RECT 414.000 1762.200 2505.600 1763.600 ;
        RECT 414.000 1756.800 2506.000 1762.200 ;
        RECT 414.400 1755.400 2506.000 1756.800 ;
        RECT 414.000 1745.920 2506.000 1755.400 ;
        RECT 414.000 1744.520 2505.600 1745.920 ;
        RECT 414.000 1737.760 2506.000 1744.520 ;
        RECT 414.400 1736.360 2506.000 1737.760 ;
        RECT 414.000 1728.240 2506.000 1736.360 ;
        RECT 414.000 1726.840 2505.600 1728.240 ;
        RECT 414.000 1720.080 2506.000 1726.840 ;
        RECT 414.400 1718.680 2506.000 1720.080 ;
        RECT 414.000 1709.200 2506.000 1718.680 ;
        RECT 414.000 1707.800 2505.600 1709.200 ;
        RECT 414.000 1701.040 2506.000 1707.800 ;
        RECT 414.400 1699.640 2506.000 1701.040 ;
        RECT 414.000 1691.520 2506.000 1699.640 ;
        RECT 414.000 1690.120 2505.600 1691.520 ;
        RECT 414.000 1683.360 2506.000 1690.120 ;
        RECT 414.400 1681.960 2506.000 1683.360 ;
        RECT 414.000 1672.480 2506.000 1681.960 ;
        RECT 414.000 1671.080 2505.600 1672.480 ;
        RECT 414.000 1664.320 2506.000 1671.080 ;
        RECT 414.400 1662.920 2506.000 1664.320 ;
        RECT 414.000 1654.800 2506.000 1662.920 ;
        RECT 414.000 1653.400 2505.600 1654.800 ;
        RECT 414.000 1646.640 2506.000 1653.400 ;
        RECT 414.400 1645.240 2506.000 1646.640 ;
        RECT 414.000 1635.760 2506.000 1645.240 ;
        RECT 414.000 1634.360 2505.600 1635.760 ;
        RECT 414.000 1628.960 2506.000 1634.360 ;
        RECT 414.400 1627.560 2506.000 1628.960 ;
        RECT 414.000 1618.080 2506.000 1627.560 ;
        RECT 414.000 1616.680 2505.600 1618.080 ;
        RECT 414.000 1609.920 2506.000 1616.680 ;
        RECT 414.400 1608.520 2506.000 1609.920 ;
        RECT 414.000 1600.400 2506.000 1608.520 ;
        RECT 414.000 1599.000 2505.600 1600.400 ;
        RECT 414.000 1592.240 2506.000 1599.000 ;
        RECT 414.400 1590.840 2506.000 1592.240 ;
        RECT 414.000 1581.360 2506.000 1590.840 ;
        RECT 414.000 1579.960 2505.600 1581.360 ;
        RECT 414.000 1573.200 2506.000 1579.960 ;
        RECT 414.400 1571.800 2506.000 1573.200 ;
        RECT 414.000 1563.680 2506.000 1571.800 ;
        RECT 414.000 1562.280 2505.600 1563.680 ;
        RECT 414.000 1555.520 2506.000 1562.280 ;
        RECT 414.400 1554.120 2506.000 1555.520 ;
        RECT 414.000 1544.640 2506.000 1554.120 ;
        RECT 414.000 1543.240 2505.600 1544.640 ;
        RECT 414.000 1536.480 2506.000 1543.240 ;
        RECT 414.400 1535.080 2506.000 1536.480 ;
        RECT 414.000 1526.960 2506.000 1535.080 ;
        RECT 414.000 1525.560 2505.600 1526.960 ;
        RECT 414.000 1518.800 2506.000 1525.560 ;
        RECT 414.400 1517.400 2506.000 1518.800 ;
        RECT 414.000 1507.920 2506.000 1517.400 ;
        RECT 414.000 1506.520 2505.600 1507.920 ;
        RECT 414.000 1501.120 2506.000 1506.520 ;
        RECT 414.400 1499.720 2506.000 1501.120 ;
        RECT 414.000 1490.240 2506.000 1499.720 ;
        RECT 414.000 1488.840 2505.600 1490.240 ;
        RECT 414.000 1482.080 2506.000 1488.840 ;
        RECT 414.400 1480.680 2506.000 1482.080 ;
        RECT 414.000 1472.560 2506.000 1480.680 ;
        RECT 414.000 1471.160 2505.600 1472.560 ;
        RECT 414.000 1464.400 2506.000 1471.160 ;
        RECT 414.400 1463.000 2506.000 1464.400 ;
        RECT 414.000 1453.520 2506.000 1463.000 ;
        RECT 414.000 1452.120 2505.600 1453.520 ;
        RECT 414.000 1445.360 2506.000 1452.120 ;
        RECT 414.400 1443.960 2506.000 1445.360 ;
        RECT 414.000 1435.840 2506.000 1443.960 ;
        RECT 414.000 1434.440 2505.600 1435.840 ;
        RECT 414.000 1427.680 2506.000 1434.440 ;
        RECT 414.400 1426.280 2506.000 1427.680 ;
        RECT 414.000 1416.800 2506.000 1426.280 ;
        RECT 414.000 1415.400 2505.600 1416.800 ;
        RECT 414.000 1408.640 2506.000 1415.400 ;
        RECT 414.400 1407.240 2506.000 1408.640 ;
        RECT 414.000 1399.120 2506.000 1407.240 ;
        RECT 414.000 1397.720 2505.600 1399.120 ;
        RECT 414.000 1390.960 2506.000 1397.720 ;
        RECT 414.400 1389.560 2506.000 1390.960 ;
        RECT 414.000 1380.080 2506.000 1389.560 ;
        RECT 414.000 1378.680 2505.600 1380.080 ;
        RECT 414.000 1373.280 2506.000 1378.680 ;
        RECT 414.400 1371.880 2506.000 1373.280 ;
        RECT 414.000 1362.400 2506.000 1371.880 ;
        RECT 414.000 1361.000 2505.600 1362.400 ;
        RECT 414.000 1354.240 2506.000 1361.000 ;
        RECT 414.400 1352.840 2506.000 1354.240 ;
        RECT 414.000 1344.720 2506.000 1352.840 ;
        RECT 414.000 1343.320 2505.600 1344.720 ;
        RECT 414.000 1336.560 2506.000 1343.320 ;
        RECT 414.400 1335.160 2506.000 1336.560 ;
        RECT 414.000 1325.680 2506.000 1335.160 ;
        RECT 414.000 1324.280 2505.600 1325.680 ;
        RECT 414.000 1317.520 2506.000 1324.280 ;
        RECT 414.400 1316.120 2506.000 1317.520 ;
        RECT 414.000 1308.000 2506.000 1316.120 ;
        RECT 414.000 1306.600 2505.600 1308.000 ;
        RECT 414.000 1299.840 2506.000 1306.600 ;
        RECT 414.400 1298.440 2506.000 1299.840 ;
        RECT 414.000 1288.960 2506.000 1298.440 ;
        RECT 414.000 1287.560 2505.600 1288.960 ;
        RECT 414.000 1280.800 2506.000 1287.560 ;
        RECT 414.400 1279.400 2506.000 1280.800 ;
        RECT 414.000 1271.280 2506.000 1279.400 ;
        RECT 414.000 1269.880 2505.600 1271.280 ;
        RECT 414.000 1263.120 2506.000 1269.880 ;
        RECT 414.400 1261.720 2506.000 1263.120 ;
        RECT 414.000 1252.240 2506.000 1261.720 ;
        RECT 414.000 1250.840 2505.600 1252.240 ;
        RECT 414.000 1245.440 2506.000 1250.840 ;
        RECT 414.400 1244.040 2506.000 1245.440 ;
        RECT 414.000 1234.560 2506.000 1244.040 ;
        RECT 414.000 1233.160 2505.600 1234.560 ;
        RECT 414.000 1226.400 2506.000 1233.160 ;
        RECT 414.400 1225.000 2506.000 1226.400 ;
        RECT 414.000 1216.880 2506.000 1225.000 ;
        RECT 414.000 1215.480 2505.600 1216.880 ;
        RECT 414.000 1208.720 2506.000 1215.480 ;
        RECT 414.400 1207.320 2506.000 1208.720 ;
        RECT 414.000 1197.840 2506.000 1207.320 ;
        RECT 414.000 1196.440 2505.600 1197.840 ;
        RECT 414.000 1189.680 2506.000 1196.440 ;
        RECT 414.400 1188.280 2506.000 1189.680 ;
        RECT 414.000 1180.160 2506.000 1188.280 ;
        RECT 414.000 1178.760 2505.600 1180.160 ;
        RECT 414.000 1172.000 2506.000 1178.760 ;
        RECT 414.400 1170.600 2506.000 1172.000 ;
        RECT 414.000 1161.120 2506.000 1170.600 ;
        RECT 414.000 1159.720 2505.600 1161.120 ;
        RECT 414.000 1152.960 2506.000 1159.720 ;
        RECT 414.400 1151.560 2506.000 1152.960 ;
        RECT 414.000 1143.440 2506.000 1151.560 ;
        RECT 414.000 1142.040 2505.600 1143.440 ;
        RECT 414.000 1135.280 2506.000 1142.040 ;
        RECT 414.400 1133.880 2506.000 1135.280 ;
        RECT 414.000 1124.400 2506.000 1133.880 ;
        RECT 414.000 1123.000 2505.600 1124.400 ;
        RECT 414.000 1117.600 2506.000 1123.000 ;
        RECT 414.400 1116.200 2506.000 1117.600 ;
        RECT 414.000 1106.720 2506.000 1116.200 ;
        RECT 414.000 1105.320 2505.600 1106.720 ;
        RECT 414.000 1098.560 2506.000 1105.320 ;
        RECT 414.400 1097.160 2506.000 1098.560 ;
        RECT 414.000 1089.040 2506.000 1097.160 ;
        RECT 414.000 1087.640 2505.600 1089.040 ;
        RECT 414.000 1080.880 2506.000 1087.640 ;
        RECT 414.400 1079.480 2506.000 1080.880 ;
        RECT 414.000 1070.000 2506.000 1079.480 ;
        RECT 414.000 1068.600 2505.600 1070.000 ;
        RECT 414.000 1061.840 2506.000 1068.600 ;
        RECT 414.400 1060.440 2506.000 1061.840 ;
        RECT 414.000 1052.320 2506.000 1060.440 ;
        RECT 414.000 1050.920 2505.600 1052.320 ;
        RECT 414.000 1044.160 2506.000 1050.920 ;
        RECT 414.400 1042.760 2506.000 1044.160 ;
        RECT 414.000 1033.280 2506.000 1042.760 ;
        RECT 414.000 1031.880 2505.600 1033.280 ;
        RECT 414.000 1025.120 2506.000 1031.880 ;
        RECT 414.400 1023.720 2506.000 1025.120 ;
        RECT 414.000 1015.600 2506.000 1023.720 ;
        RECT 414.000 1014.200 2505.600 1015.600 ;
        RECT 414.000 1007.440 2506.000 1014.200 ;
        RECT 414.400 1006.040 2506.000 1007.440 ;
        RECT 414.000 996.560 2506.000 1006.040 ;
        RECT 414.000 995.160 2505.600 996.560 ;
        RECT 414.000 989.760 2506.000 995.160 ;
        RECT 414.400 988.360 2506.000 989.760 ;
        RECT 414.000 978.880 2506.000 988.360 ;
        RECT 414.000 977.480 2505.600 978.880 ;
        RECT 414.000 970.720 2506.000 977.480 ;
        RECT 414.400 969.320 2506.000 970.720 ;
        RECT 414.000 961.200 2506.000 969.320 ;
        RECT 414.000 959.800 2505.600 961.200 ;
        RECT 414.000 953.040 2506.000 959.800 ;
        RECT 414.400 951.640 2506.000 953.040 ;
        RECT 414.000 942.160 2506.000 951.640 ;
        RECT 414.000 940.760 2505.600 942.160 ;
        RECT 414.000 934.000 2506.000 940.760 ;
        RECT 414.400 932.600 2506.000 934.000 ;
        RECT 414.000 924.480 2506.000 932.600 ;
        RECT 414.000 923.080 2505.600 924.480 ;
        RECT 414.000 916.320 2506.000 923.080 ;
        RECT 414.400 914.920 2506.000 916.320 ;
        RECT 414.000 905.440 2506.000 914.920 ;
        RECT 414.000 904.040 2505.600 905.440 ;
        RECT 414.000 897.280 2506.000 904.040 ;
        RECT 414.400 895.880 2506.000 897.280 ;
        RECT 414.000 887.760 2506.000 895.880 ;
        RECT 414.000 886.360 2505.600 887.760 ;
        RECT 414.000 879.600 2506.000 886.360 ;
        RECT 414.400 878.200 2506.000 879.600 ;
        RECT 414.000 868.720 2506.000 878.200 ;
        RECT 414.000 867.320 2505.600 868.720 ;
        RECT 414.000 861.920 2506.000 867.320 ;
        RECT 414.400 860.520 2506.000 861.920 ;
        RECT 414.000 851.040 2506.000 860.520 ;
        RECT 414.000 849.640 2505.600 851.040 ;
        RECT 414.000 842.880 2506.000 849.640 ;
        RECT 414.400 841.480 2506.000 842.880 ;
        RECT 414.000 833.360 2506.000 841.480 ;
        RECT 414.000 831.960 2505.600 833.360 ;
        RECT 414.000 825.200 2506.000 831.960 ;
        RECT 414.400 823.800 2506.000 825.200 ;
        RECT 414.000 814.320 2506.000 823.800 ;
        RECT 414.000 812.920 2505.600 814.320 ;
        RECT 414.000 806.160 2506.000 812.920 ;
        RECT 414.400 804.760 2506.000 806.160 ;
        RECT 414.000 796.640 2506.000 804.760 ;
        RECT 414.000 795.240 2505.600 796.640 ;
        RECT 414.000 788.480 2506.000 795.240 ;
        RECT 414.400 787.080 2506.000 788.480 ;
        RECT 414.000 777.600 2506.000 787.080 ;
        RECT 414.000 776.200 2505.600 777.600 ;
        RECT 414.000 769.440 2506.000 776.200 ;
        RECT 414.400 768.040 2506.000 769.440 ;
        RECT 414.000 759.920 2506.000 768.040 ;
        RECT 414.000 758.520 2505.600 759.920 ;
        RECT 414.000 751.760 2506.000 758.520 ;
        RECT 414.400 750.360 2506.000 751.760 ;
        RECT 414.000 740.880 2506.000 750.360 ;
        RECT 414.000 739.480 2505.600 740.880 ;
        RECT 414.000 734.080 2506.000 739.480 ;
        RECT 414.400 732.680 2506.000 734.080 ;
        RECT 414.000 723.200 2506.000 732.680 ;
        RECT 414.000 721.800 2505.600 723.200 ;
        RECT 414.000 715.040 2506.000 721.800 ;
        RECT 414.400 713.640 2506.000 715.040 ;
        RECT 414.000 705.520 2506.000 713.640 ;
        RECT 414.000 704.120 2505.600 705.520 ;
        RECT 414.000 697.360 2506.000 704.120 ;
        RECT 414.400 695.960 2506.000 697.360 ;
        RECT 414.000 686.480 2506.000 695.960 ;
        RECT 414.000 685.080 2505.600 686.480 ;
        RECT 414.000 678.320 2506.000 685.080 ;
        RECT 414.400 676.920 2506.000 678.320 ;
        RECT 414.000 668.800 2506.000 676.920 ;
        RECT 414.000 667.400 2505.600 668.800 ;
        RECT 414.000 660.640 2506.000 667.400 ;
        RECT 414.400 659.240 2506.000 660.640 ;
        RECT 414.000 649.760 2506.000 659.240 ;
        RECT 414.000 648.360 2505.600 649.760 ;
        RECT 414.000 641.600 2506.000 648.360 ;
        RECT 414.400 640.200 2506.000 641.600 ;
        RECT 414.000 632.080 2506.000 640.200 ;
        RECT 414.000 630.680 2505.600 632.080 ;
        RECT 414.000 623.920 2506.000 630.680 ;
        RECT 414.400 622.520 2506.000 623.920 ;
        RECT 414.000 613.040 2506.000 622.520 ;
        RECT 414.000 611.640 2505.600 613.040 ;
        RECT 414.000 606.240 2506.000 611.640 ;
        RECT 414.400 604.840 2506.000 606.240 ;
        RECT 414.000 595.360 2506.000 604.840 ;
        RECT 414.000 593.960 2505.600 595.360 ;
        RECT 414.000 587.200 2506.000 593.960 ;
        RECT 414.400 585.800 2506.000 587.200 ;
        RECT 414.000 577.680 2506.000 585.800 ;
        RECT 414.000 576.280 2505.600 577.680 ;
        RECT 414.000 569.520 2506.000 576.280 ;
        RECT 414.400 568.120 2506.000 569.520 ;
        RECT 414.000 558.640 2506.000 568.120 ;
        RECT 414.000 557.240 2505.600 558.640 ;
        RECT 414.000 550.480 2506.000 557.240 ;
        RECT 414.400 549.080 2506.000 550.480 ;
        RECT 414.000 540.960 2506.000 549.080 ;
        RECT 414.000 539.560 2505.600 540.960 ;
        RECT 414.000 532.800 2506.000 539.560 ;
        RECT 414.400 531.400 2506.000 532.800 ;
        RECT 414.000 521.920 2506.000 531.400 ;
        RECT 414.000 520.520 2505.600 521.920 ;
        RECT 414.000 514.255 2506.000 520.520 ;
      LAYER via3 ;
        RECT 2025.220 3006.460 2025.540 3006.780 ;
        RECT 2025.220 2999.660 2025.540 2999.980 ;
      LAYER met4 ;
        RECT 2025.215 3006.455 2025.545 3006.785 ;
        RECT 2025.230 2999.985 2025.530 3006.455 ;
        RECT 2025.215 2999.655 2025.545 2999.985 ;
      LAYER met4 ;
        RECT 422.255 520.640 430.640 2999.040 ;
      LAYER met4 ;
        RECT 431.040 520.640 432.640 2999.040 ;
      LAYER met4 ;
        RECT 433.040 520.640 507.440 2999.040 ;
      LAYER met4 ;
        RECT 507.840 520.640 509.440 2999.040 ;
      LAYER met4 ;
        RECT 509.840 2997.690 2429.440 2999.040 ;
        RECT 509.840 2996.510 2024.790 2997.690 ;
        RECT 2025.970 2996.510 2429.440 2997.690 ;
        RECT 509.840 520.640 2429.440 2996.510 ;
  END
END user_project_wrapper
END LIBRARY

