VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Ibtida_top_dffram_cv
  CLASS BLOCK ;
  FOREIGN Ibtida_top_dffram_cv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1591.465 BY 1602.185 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 17.720 1591.465 18.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1085.320 1591.465 1085.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1192.080 1591.465 1192.680 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1298.840 1591.465 1299.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1405.600 1591.465 1406.200 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1512.360 1591.465 1512.960 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1561.790 1598.185 1562.070 1602.185 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1385.150 1598.185 1385.430 1602.185 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.050 1598.185 1208.330 1602.185 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.410 1598.185 1031.690 1602.185 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.770 1598.185 855.050 1602.185 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 124.480 1591.465 125.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 677.670 1598.185 677.950 1602.185 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.030 1598.185 501.310 1602.185 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 1598.185 324.210 1602.185 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 1598.185 147.570 1602.185 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1582.400 4.000 1583.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.160 4.000 1468.760 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.920 4.000 1354.520 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 231.240 1591.465 231.840 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 781.360 4.000 781.960 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 338.000 1591.465 338.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 444.760 1591.465 445.360 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 551.520 1591.465 552.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 658.280 1591.465 658.880 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 765.040 1591.465 765.640 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 871.800 1591.465 872.400 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1587.465 978.560 1591.465 979.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 88.440 1591.465 89.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1156.720 1591.465 1157.320 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1263.480 1591.465 1264.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1370.240 1591.465 1370.840 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1477.000 1591.465 1477.600 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1583.760 1591.465 1584.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.030 1598.185 1444.310 1602.185 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1267.390 1598.185 1267.670 1602.185 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1090.290 1598.185 1090.570 1602.185 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.650 1598.185 913.930 1602.185 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 736.550 1598.185 736.830 1602.185 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 195.200 1591.465 195.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.910 1598.185 560.190 1602.185 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.810 1598.185 383.090 1602.185 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.170 1598.185 206.450 1602.185 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.530 1598.185 29.810 1602.185 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.240 4.000 1506.840 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.760 4.000 1278.360 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 301.960 1591.465 302.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 408.720 1591.465 409.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 515.480 1591.465 516.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 622.920 1591.465 623.520 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 729.680 1591.465 730.280 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 836.440 1591.465 837.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 943.200 1591.465 943.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1049.960 1591.465 1050.560 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 53.080 1591.465 53.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1121.360 1591.465 1121.960 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1228.120 1591.465 1228.720 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1334.880 1591.465 1335.480 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1441.640 1591.465 1442.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1548.400 1591.465 1549.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1502.910 1598.185 1503.190 1602.185 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1326.270 1598.185 1326.550 1602.185 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1149.170 1598.185 1149.450 1602.185 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.530 1598.185 972.810 1602.185 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.430 1598.185 795.710 1602.185 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 159.840 1591.465 160.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 618.790 1598.185 619.070 1602.185 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.150 1598.185 442.430 1602.185 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.050 1598.185 265.330 1602.185 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 1598.185 88.690 1602.185 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1544.320 4.000 1544.920 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.080 4.000 1430.680 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.920 4.000 1201.520 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.680 4.000 1087.280 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 266.600 1591.465 267.200 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 373.360 1591.465 373.960 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 480.120 1591.465 480.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 586.880 1591.465 587.480 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 693.640 1591.465 694.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 800.400 1591.465 801.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 907.160 1591.465 907.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1587.465 1013.920 1591.465 1014.520 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1296.370 0.000 1296.650 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1321.210 0.000 1321.490 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.630 0.000 1333.910 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.470 0.000 1358.750 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.850 0.000 1383.130 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.270 0.000 1395.550 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1432.530 0.000 1432.810 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.950 0.000 1445.230 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1457.370 0.000 1457.650 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1469.790 0.000 1470.070 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.750 0.000 1482.030 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.590 0.000 1506.870 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1531.430 0.000 1531.710 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1543.850 0.000 1544.130 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1556.270 0.000 1556.550 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1568.690 0.000 1568.970 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.770 0.000 901.050 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.150 0.000 925.430 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.570 0.000 937.850 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.470 0.000 1036.750 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.890 0.000 1049.170 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.630 0.000 1172.910 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1209.890 0.000 1210.170 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.310 0.000 1222.590 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.730 0.000 1235.010 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1251.290 0.000 1251.570 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.250 0.000 1263.530 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1275.670 0.000 1275.950 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.510 0.000 1300.790 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.930 0.000 1313.210 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1337.770 0.000 1338.050 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1350.190 0.000 1350.470 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1362.610 0.000 1362.890 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1374.570 0.000 1374.850 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1386.990 0.000 1387.270 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1399.410 0.000 1399.690 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1411.830 0.000 1412.110 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1424.250 0.000 1424.530 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1436.670 0.000 1436.950 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1510.730 0.000 1511.010 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1535.570 0.000 1535.850 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1547.990 0.000 1548.270 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1560.410 0.000 1560.690 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1585.250 0.000 1585.530 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1028.190 0.000 1028.470 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.870 0.000 1078.150 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1115.130 0.000 1115.410 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1127.550 0.000 1127.830 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.510 0.000 1139.790 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1238.870 0.000 1239.150 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1254.970 0.000 1255.250 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1267.390 0.000 1267.670 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1279.810 0.000 1280.090 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.230 0.000 1292.510 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.650 0.000 1304.930 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1329.490 0.000 1329.770 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1366.290 0.000 1366.570 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.710 0.000 1378.990 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.970 0.000 1416.250 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1440.810 0.000 1441.090 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.230 0.000 1453.510 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.650 0.000 1465.930 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1502.450 0.000 1502.730 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1514.870 0.000 1515.150 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1527.290 0.000 1527.570 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.970 0.000 1577.250 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.390 0.000 1589.670 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 970.690 0.000 970.970 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.530 0.000 995.810 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.170 0.000 1057.450 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.330 0.000 1193.610 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_rst_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1591.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1591.440 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1585.620 1591.285 ;
      LAYER met1 ;
        RECT 0.070 10.640 1585.620 1597.960 ;
      LAYER met2 ;
        RECT 0.090 1597.905 29.250 1598.185 ;
        RECT 30.090 1597.905 88.130 1598.185 ;
        RECT 88.970 1597.905 147.010 1598.185 ;
        RECT 147.850 1597.905 205.890 1598.185 ;
        RECT 206.730 1597.905 264.770 1598.185 ;
        RECT 265.610 1597.905 323.650 1598.185 ;
        RECT 324.490 1597.905 382.530 1598.185 ;
        RECT 383.370 1597.905 441.870 1598.185 ;
        RECT 442.710 1597.905 500.750 1598.185 ;
        RECT 501.590 1597.905 559.630 1598.185 ;
        RECT 560.470 1597.905 618.510 1598.185 ;
        RECT 619.350 1597.905 677.390 1598.185 ;
        RECT 678.230 1597.905 736.270 1598.185 ;
        RECT 737.110 1597.905 795.150 1598.185 ;
        RECT 795.990 1597.905 854.490 1598.185 ;
        RECT 855.330 1597.905 913.370 1598.185 ;
        RECT 914.210 1597.905 972.250 1598.185 ;
        RECT 973.090 1597.905 1031.130 1598.185 ;
        RECT 1031.970 1597.905 1090.010 1598.185 ;
        RECT 1090.850 1597.905 1148.890 1598.185 ;
        RECT 1149.730 1597.905 1207.770 1598.185 ;
        RECT 1208.610 1597.905 1267.110 1598.185 ;
        RECT 1267.950 1597.905 1325.990 1598.185 ;
        RECT 1326.830 1597.905 1384.870 1598.185 ;
        RECT 1385.710 1597.905 1443.750 1598.185 ;
        RECT 1444.590 1597.905 1502.630 1598.185 ;
        RECT 1503.470 1597.905 1561.510 1598.185 ;
        RECT 1562.350 1597.905 1585.520 1598.185 ;
        RECT 0.090 4.280 1585.520 1597.905 ;
        RECT 0.090 4.000 1.650 4.280 ;
        RECT 2.490 4.000 5.330 4.280 ;
        RECT 6.170 4.000 9.470 4.280 ;
        RECT 10.310 4.000 13.610 4.280 ;
        RECT 14.450 4.000 17.750 4.280 ;
        RECT 18.590 4.000 21.890 4.280 ;
        RECT 22.730 4.000 26.030 4.280 ;
        RECT 26.870 4.000 30.170 4.280 ;
        RECT 31.010 4.000 34.310 4.280 ;
        RECT 35.150 4.000 38.450 4.280 ;
        RECT 39.290 4.000 42.590 4.280 ;
        RECT 43.430 4.000 46.730 4.280 ;
        RECT 47.570 4.000 50.870 4.280 ;
        RECT 51.710 4.000 55.010 4.280 ;
        RECT 55.850 4.000 59.150 4.280 ;
        RECT 59.990 4.000 63.290 4.280 ;
        RECT 64.130 4.000 67.430 4.280 ;
        RECT 68.270 4.000 71.570 4.280 ;
        RECT 72.410 4.000 75.710 4.280 ;
        RECT 76.550 4.000 79.850 4.280 ;
        RECT 80.690 4.000 83.990 4.280 ;
        RECT 84.830 4.000 88.130 4.280 ;
        RECT 88.970 4.000 92.270 4.280 ;
        RECT 93.110 4.000 96.410 4.280 ;
        RECT 97.250 4.000 100.550 4.280 ;
        RECT 101.390 4.000 104.690 4.280 ;
        RECT 105.530 4.000 108.830 4.280 ;
        RECT 109.670 4.000 112.970 4.280 ;
        RECT 113.810 4.000 116.650 4.280 ;
        RECT 117.490 4.000 120.790 4.280 ;
        RECT 121.630 4.000 124.930 4.280 ;
        RECT 125.770 4.000 129.070 4.280 ;
        RECT 129.910 4.000 133.210 4.280 ;
        RECT 134.050 4.000 137.350 4.280 ;
        RECT 138.190 4.000 141.490 4.280 ;
        RECT 142.330 4.000 145.630 4.280 ;
        RECT 146.470 4.000 149.770 4.280 ;
        RECT 150.610 4.000 153.910 4.280 ;
        RECT 154.750 4.000 158.050 4.280 ;
        RECT 158.890 4.000 162.190 4.280 ;
        RECT 163.030 4.000 166.330 4.280 ;
        RECT 167.170 4.000 170.470 4.280 ;
        RECT 171.310 4.000 174.610 4.280 ;
        RECT 175.450 4.000 178.750 4.280 ;
        RECT 179.590 4.000 182.890 4.280 ;
        RECT 183.730 4.000 187.030 4.280 ;
        RECT 187.870 4.000 191.170 4.280 ;
        RECT 192.010 4.000 195.310 4.280 ;
        RECT 196.150 4.000 199.450 4.280 ;
        RECT 200.290 4.000 203.590 4.280 ;
        RECT 204.430 4.000 207.730 4.280 ;
        RECT 208.570 4.000 211.870 4.280 ;
        RECT 212.710 4.000 216.010 4.280 ;
        RECT 216.850 4.000 220.150 4.280 ;
        RECT 220.990 4.000 224.290 4.280 ;
        RECT 225.130 4.000 228.430 4.280 ;
        RECT 229.270 4.000 232.110 4.280 ;
        RECT 232.950 4.000 236.250 4.280 ;
        RECT 237.090 4.000 240.390 4.280 ;
        RECT 241.230 4.000 244.530 4.280 ;
        RECT 245.370 4.000 248.670 4.280 ;
        RECT 249.510 4.000 252.810 4.280 ;
        RECT 253.650 4.000 256.950 4.280 ;
        RECT 257.790 4.000 261.090 4.280 ;
        RECT 261.930 4.000 265.230 4.280 ;
        RECT 266.070 4.000 269.370 4.280 ;
        RECT 270.210 4.000 273.510 4.280 ;
        RECT 274.350 4.000 277.650 4.280 ;
        RECT 278.490 4.000 281.790 4.280 ;
        RECT 282.630 4.000 285.930 4.280 ;
        RECT 286.770 4.000 290.070 4.280 ;
        RECT 290.910 4.000 294.210 4.280 ;
        RECT 295.050 4.000 298.350 4.280 ;
        RECT 299.190 4.000 302.490 4.280 ;
        RECT 303.330 4.000 306.630 4.280 ;
        RECT 307.470 4.000 310.770 4.280 ;
        RECT 311.610 4.000 314.910 4.280 ;
        RECT 315.750 4.000 319.050 4.280 ;
        RECT 319.890 4.000 323.190 4.280 ;
        RECT 324.030 4.000 327.330 4.280 ;
        RECT 328.170 4.000 331.470 4.280 ;
        RECT 332.310 4.000 335.610 4.280 ;
        RECT 336.450 4.000 339.750 4.280 ;
        RECT 340.590 4.000 343.430 4.280 ;
        RECT 344.270 4.000 347.570 4.280 ;
        RECT 348.410 4.000 351.710 4.280 ;
        RECT 352.550 4.000 355.850 4.280 ;
        RECT 356.690 4.000 359.990 4.280 ;
        RECT 360.830 4.000 364.130 4.280 ;
        RECT 364.970 4.000 368.270 4.280 ;
        RECT 369.110 4.000 372.410 4.280 ;
        RECT 373.250 4.000 376.550 4.280 ;
        RECT 377.390 4.000 380.690 4.280 ;
        RECT 381.530 4.000 384.830 4.280 ;
        RECT 385.670 4.000 388.970 4.280 ;
        RECT 389.810 4.000 393.110 4.280 ;
        RECT 393.950 4.000 397.250 4.280 ;
        RECT 398.090 4.000 401.390 4.280 ;
        RECT 402.230 4.000 405.530 4.280 ;
        RECT 406.370 4.000 409.670 4.280 ;
        RECT 410.510 4.000 413.810 4.280 ;
        RECT 414.650 4.000 417.950 4.280 ;
        RECT 418.790 4.000 422.090 4.280 ;
        RECT 422.930 4.000 426.230 4.280 ;
        RECT 427.070 4.000 430.370 4.280 ;
        RECT 431.210 4.000 434.510 4.280 ;
        RECT 435.350 4.000 438.650 4.280 ;
        RECT 439.490 4.000 442.790 4.280 ;
        RECT 443.630 4.000 446.930 4.280 ;
        RECT 447.770 4.000 451.070 4.280 ;
        RECT 451.910 4.000 455.210 4.280 ;
        RECT 456.050 4.000 458.890 4.280 ;
        RECT 459.730 4.000 463.030 4.280 ;
        RECT 463.870 4.000 467.170 4.280 ;
        RECT 468.010 4.000 471.310 4.280 ;
        RECT 472.150 4.000 475.450 4.280 ;
        RECT 476.290 4.000 479.590 4.280 ;
        RECT 480.430 4.000 483.730 4.280 ;
        RECT 484.570 4.000 487.870 4.280 ;
        RECT 488.710 4.000 492.010 4.280 ;
        RECT 492.850 4.000 496.150 4.280 ;
        RECT 496.990 4.000 500.290 4.280 ;
        RECT 501.130 4.000 504.430 4.280 ;
        RECT 505.270 4.000 508.570 4.280 ;
        RECT 509.410 4.000 512.710 4.280 ;
        RECT 513.550 4.000 516.850 4.280 ;
        RECT 517.690 4.000 520.990 4.280 ;
        RECT 521.830 4.000 525.130 4.280 ;
        RECT 525.970 4.000 529.270 4.280 ;
        RECT 530.110 4.000 533.410 4.280 ;
        RECT 534.250 4.000 537.550 4.280 ;
        RECT 538.390 4.000 541.690 4.280 ;
        RECT 542.530 4.000 545.830 4.280 ;
        RECT 546.670 4.000 549.970 4.280 ;
        RECT 550.810 4.000 554.110 4.280 ;
        RECT 554.950 4.000 558.250 4.280 ;
        RECT 559.090 4.000 562.390 4.280 ;
        RECT 563.230 4.000 566.530 4.280 ;
        RECT 567.370 4.000 570.210 4.280 ;
        RECT 571.050 4.000 574.350 4.280 ;
        RECT 575.190 4.000 578.490 4.280 ;
        RECT 579.330 4.000 582.630 4.280 ;
        RECT 583.470 4.000 586.770 4.280 ;
        RECT 587.610 4.000 590.910 4.280 ;
        RECT 591.750 4.000 595.050 4.280 ;
        RECT 595.890 4.000 599.190 4.280 ;
        RECT 600.030 4.000 603.330 4.280 ;
        RECT 604.170 4.000 607.470 4.280 ;
        RECT 608.310 4.000 611.610 4.280 ;
        RECT 612.450 4.000 615.750 4.280 ;
        RECT 616.590 4.000 619.890 4.280 ;
        RECT 620.730 4.000 624.030 4.280 ;
        RECT 624.870 4.000 628.170 4.280 ;
        RECT 629.010 4.000 632.310 4.280 ;
        RECT 633.150 4.000 636.450 4.280 ;
        RECT 637.290 4.000 640.590 4.280 ;
        RECT 641.430 4.000 644.730 4.280 ;
        RECT 645.570 4.000 648.870 4.280 ;
        RECT 649.710 4.000 653.010 4.280 ;
        RECT 653.850 4.000 657.150 4.280 ;
        RECT 657.990 4.000 661.290 4.280 ;
        RECT 662.130 4.000 665.430 4.280 ;
        RECT 666.270 4.000 669.570 4.280 ;
        RECT 670.410 4.000 673.710 4.280 ;
        RECT 674.550 4.000 677.850 4.280 ;
        RECT 678.690 4.000 681.990 4.280 ;
        RECT 682.830 4.000 685.670 4.280 ;
        RECT 686.510 4.000 689.810 4.280 ;
        RECT 690.650 4.000 693.950 4.280 ;
        RECT 694.790 4.000 698.090 4.280 ;
        RECT 698.930 4.000 702.230 4.280 ;
        RECT 703.070 4.000 706.370 4.280 ;
        RECT 707.210 4.000 710.510 4.280 ;
        RECT 711.350 4.000 714.650 4.280 ;
        RECT 715.490 4.000 718.790 4.280 ;
        RECT 719.630 4.000 722.930 4.280 ;
        RECT 723.770 4.000 727.070 4.280 ;
        RECT 727.910 4.000 731.210 4.280 ;
        RECT 732.050 4.000 735.350 4.280 ;
        RECT 736.190 4.000 739.490 4.280 ;
        RECT 740.330 4.000 743.630 4.280 ;
        RECT 744.470 4.000 747.770 4.280 ;
        RECT 748.610 4.000 751.910 4.280 ;
        RECT 752.750 4.000 756.050 4.280 ;
        RECT 756.890 4.000 760.190 4.280 ;
        RECT 761.030 4.000 764.330 4.280 ;
        RECT 765.170 4.000 768.470 4.280 ;
        RECT 769.310 4.000 772.610 4.280 ;
        RECT 773.450 4.000 776.750 4.280 ;
        RECT 777.590 4.000 780.890 4.280 ;
        RECT 781.730 4.000 785.030 4.280 ;
        RECT 785.870 4.000 789.170 4.280 ;
        RECT 790.010 4.000 793.310 4.280 ;
        RECT 794.150 4.000 797.450 4.280 ;
        RECT 798.290 4.000 801.130 4.280 ;
        RECT 801.970 4.000 805.270 4.280 ;
        RECT 806.110 4.000 809.410 4.280 ;
        RECT 810.250 4.000 813.550 4.280 ;
        RECT 814.390 4.000 817.690 4.280 ;
        RECT 818.530 4.000 821.830 4.280 ;
        RECT 822.670 4.000 825.970 4.280 ;
        RECT 826.810 4.000 830.110 4.280 ;
        RECT 830.950 4.000 834.250 4.280 ;
        RECT 835.090 4.000 838.390 4.280 ;
        RECT 839.230 4.000 842.530 4.280 ;
        RECT 843.370 4.000 846.670 4.280 ;
        RECT 847.510 4.000 850.810 4.280 ;
        RECT 851.650 4.000 854.950 4.280 ;
        RECT 855.790 4.000 859.090 4.280 ;
        RECT 859.930 4.000 863.230 4.280 ;
        RECT 864.070 4.000 867.370 4.280 ;
        RECT 868.210 4.000 871.510 4.280 ;
        RECT 872.350 4.000 875.650 4.280 ;
        RECT 876.490 4.000 879.790 4.280 ;
        RECT 880.630 4.000 883.930 4.280 ;
        RECT 884.770 4.000 888.070 4.280 ;
        RECT 888.910 4.000 892.210 4.280 ;
        RECT 893.050 4.000 896.350 4.280 ;
        RECT 897.190 4.000 900.490 4.280 ;
        RECT 901.330 4.000 904.630 4.280 ;
        RECT 905.470 4.000 908.770 4.280 ;
        RECT 909.610 4.000 912.450 4.280 ;
        RECT 913.290 4.000 916.590 4.280 ;
        RECT 917.430 4.000 920.730 4.280 ;
        RECT 921.570 4.000 924.870 4.280 ;
        RECT 925.710 4.000 929.010 4.280 ;
        RECT 929.850 4.000 933.150 4.280 ;
        RECT 933.990 4.000 937.290 4.280 ;
        RECT 938.130 4.000 941.430 4.280 ;
        RECT 942.270 4.000 945.570 4.280 ;
        RECT 946.410 4.000 949.710 4.280 ;
        RECT 950.550 4.000 953.850 4.280 ;
        RECT 954.690 4.000 957.990 4.280 ;
        RECT 958.830 4.000 962.130 4.280 ;
        RECT 962.970 4.000 966.270 4.280 ;
        RECT 967.110 4.000 970.410 4.280 ;
        RECT 971.250 4.000 974.550 4.280 ;
        RECT 975.390 4.000 978.690 4.280 ;
        RECT 979.530 4.000 982.830 4.280 ;
        RECT 983.670 4.000 986.970 4.280 ;
        RECT 987.810 4.000 991.110 4.280 ;
        RECT 991.950 4.000 995.250 4.280 ;
        RECT 996.090 4.000 999.390 4.280 ;
        RECT 1000.230 4.000 1003.530 4.280 ;
        RECT 1004.370 4.000 1007.670 4.280 ;
        RECT 1008.510 4.000 1011.810 4.280 ;
        RECT 1012.650 4.000 1015.950 4.280 ;
        RECT 1016.790 4.000 1020.090 4.280 ;
        RECT 1020.930 4.000 1024.230 4.280 ;
        RECT 1025.070 4.000 1027.910 4.280 ;
        RECT 1028.750 4.000 1032.050 4.280 ;
        RECT 1032.890 4.000 1036.190 4.280 ;
        RECT 1037.030 4.000 1040.330 4.280 ;
        RECT 1041.170 4.000 1044.470 4.280 ;
        RECT 1045.310 4.000 1048.610 4.280 ;
        RECT 1049.450 4.000 1052.750 4.280 ;
        RECT 1053.590 4.000 1056.890 4.280 ;
        RECT 1057.730 4.000 1061.030 4.280 ;
        RECT 1061.870 4.000 1065.170 4.280 ;
        RECT 1066.010 4.000 1069.310 4.280 ;
        RECT 1070.150 4.000 1073.450 4.280 ;
        RECT 1074.290 4.000 1077.590 4.280 ;
        RECT 1078.430 4.000 1081.730 4.280 ;
        RECT 1082.570 4.000 1085.870 4.280 ;
        RECT 1086.710 4.000 1090.010 4.280 ;
        RECT 1090.850 4.000 1094.150 4.280 ;
        RECT 1094.990 4.000 1098.290 4.280 ;
        RECT 1099.130 4.000 1102.430 4.280 ;
        RECT 1103.270 4.000 1106.570 4.280 ;
        RECT 1107.410 4.000 1110.710 4.280 ;
        RECT 1111.550 4.000 1114.850 4.280 ;
        RECT 1115.690 4.000 1118.990 4.280 ;
        RECT 1119.830 4.000 1123.130 4.280 ;
        RECT 1123.970 4.000 1127.270 4.280 ;
        RECT 1128.110 4.000 1131.410 4.280 ;
        RECT 1132.250 4.000 1135.550 4.280 ;
        RECT 1136.390 4.000 1139.230 4.280 ;
        RECT 1140.070 4.000 1143.370 4.280 ;
        RECT 1144.210 4.000 1147.510 4.280 ;
        RECT 1148.350 4.000 1151.650 4.280 ;
        RECT 1152.490 4.000 1155.790 4.280 ;
        RECT 1156.630 4.000 1159.930 4.280 ;
        RECT 1160.770 4.000 1164.070 4.280 ;
        RECT 1164.910 4.000 1168.210 4.280 ;
        RECT 1169.050 4.000 1172.350 4.280 ;
        RECT 1173.190 4.000 1176.490 4.280 ;
        RECT 1177.330 4.000 1180.630 4.280 ;
        RECT 1181.470 4.000 1184.770 4.280 ;
        RECT 1185.610 4.000 1188.910 4.280 ;
        RECT 1189.750 4.000 1193.050 4.280 ;
        RECT 1193.890 4.000 1197.190 4.280 ;
        RECT 1198.030 4.000 1201.330 4.280 ;
        RECT 1202.170 4.000 1205.470 4.280 ;
        RECT 1206.310 4.000 1209.610 4.280 ;
        RECT 1210.450 4.000 1213.750 4.280 ;
        RECT 1214.590 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1222.030 4.280 ;
        RECT 1222.870 4.000 1226.170 4.280 ;
        RECT 1227.010 4.000 1230.310 4.280 ;
        RECT 1231.150 4.000 1234.450 4.280 ;
        RECT 1235.290 4.000 1238.590 4.280 ;
        RECT 1239.430 4.000 1242.730 4.280 ;
        RECT 1243.570 4.000 1246.870 4.280 ;
        RECT 1247.710 4.000 1251.010 4.280 ;
        RECT 1251.850 4.000 1254.690 4.280 ;
        RECT 1255.530 4.000 1258.830 4.280 ;
        RECT 1259.670 4.000 1262.970 4.280 ;
        RECT 1263.810 4.000 1267.110 4.280 ;
        RECT 1267.950 4.000 1271.250 4.280 ;
        RECT 1272.090 4.000 1275.390 4.280 ;
        RECT 1276.230 4.000 1279.530 4.280 ;
        RECT 1280.370 4.000 1283.670 4.280 ;
        RECT 1284.510 4.000 1287.810 4.280 ;
        RECT 1288.650 4.000 1291.950 4.280 ;
        RECT 1292.790 4.000 1296.090 4.280 ;
        RECT 1296.930 4.000 1300.230 4.280 ;
        RECT 1301.070 4.000 1304.370 4.280 ;
        RECT 1305.210 4.000 1308.510 4.280 ;
        RECT 1309.350 4.000 1312.650 4.280 ;
        RECT 1313.490 4.000 1316.790 4.280 ;
        RECT 1317.630 4.000 1320.930 4.280 ;
        RECT 1321.770 4.000 1325.070 4.280 ;
        RECT 1325.910 4.000 1329.210 4.280 ;
        RECT 1330.050 4.000 1333.350 4.280 ;
        RECT 1334.190 4.000 1337.490 4.280 ;
        RECT 1338.330 4.000 1341.630 4.280 ;
        RECT 1342.470 4.000 1345.770 4.280 ;
        RECT 1346.610 4.000 1349.910 4.280 ;
        RECT 1350.750 4.000 1354.050 4.280 ;
        RECT 1354.890 4.000 1358.190 4.280 ;
        RECT 1359.030 4.000 1362.330 4.280 ;
        RECT 1363.170 4.000 1366.010 4.280 ;
        RECT 1366.850 4.000 1370.150 4.280 ;
        RECT 1370.990 4.000 1374.290 4.280 ;
        RECT 1375.130 4.000 1378.430 4.280 ;
        RECT 1379.270 4.000 1382.570 4.280 ;
        RECT 1383.410 4.000 1386.710 4.280 ;
        RECT 1387.550 4.000 1390.850 4.280 ;
        RECT 1391.690 4.000 1394.990 4.280 ;
        RECT 1395.830 4.000 1399.130 4.280 ;
        RECT 1399.970 4.000 1403.270 4.280 ;
        RECT 1404.110 4.000 1407.410 4.280 ;
        RECT 1408.250 4.000 1411.550 4.280 ;
        RECT 1412.390 4.000 1415.690 4.280 ;
        RECT 1416.530 4.000 1419.830 4.280 ;
        RECT 1420.670 4.000 1423.970 4.280 ;
        RECT 1424.810 4.000 1428.110 4.280 ;
        RECT 1428.950 4.000 1432.250 4.280 ;
        RECT 1433.090 4.000 1436.390 4.280 ;
        RECT 1437.230 4.000 1440.530 4.280 ;
        RECT 1441.370 4.000 1444.670 4.280 ;
        RECT 1445.510 4.000 1448.810 4.280 ;
        RECT 1449.650 4.000 1452.950 4.280 ;
        RECT 1453.790 4.000 1457.090 4.280 ;
        RECT 1457.930 4.000 1461.230 4.280 ;
        RECT 1462.070 4.000 1465.370 4.280 ;
        RECT 1466.210 4.000 1469.510 4.280 ;
        RECT 1470.350 4.000 1473.650 4.280 ;
        RECT 1474.490 4.000 1477.790 4.280 ;
        RECT 1478.630 4.000 1481.470 4.280 ;
        RECT 1482.310 4.000 1485.610 4.280 ;
        RECT 1486.450 4.000 1489.750 4.280 ;
        RECT 1490.590 4.000 1493.890 4.280 ;
        RECT 1494.730 4.000 1498.030 4.280 ;
        RECT 1498.870 4.000 1502.170 4.280 ;
        RECT 1503.010 4.000 1506.310 4.280 ;
        RECT 1507.150 4.000 1510.450 4.280 ;
        RECT 1511.290 4.000 1514.590 4.280 ;
        RECT 1515.430 4.000 1518.730 4.280 ;
        RECT 1519.570 4.000 1522.870 4.280 ;
        RECT 1523.710 4.000 1527.010 4.280 ;
        RECT 1527.850 4.000 1531.150 4.280 ;
        RECT 1531.990 4.000 1535.290 4.280 ;
        RECT 1536.130 4.000 1539.430 4.280 ;
        RECT 1540.270 4.000 1543.570 4.280 ;
        RECT 1544.410 4.000 1547.710 4.280 ;
        RECT 1548.550 4.000 1551.850 4.280 ;
        RECT 1552.690 4.000 1555.990 4.280 ;
        RECT 1556.830 4.000 1560.130 4.280 ;
        RECT 1560.970 4.000 1564.270 4.280 ;
        RECT 1565.110 4.000 1568.410 4.280 ;
        RECT 1569.250 4.000 1572.550 4.280 ;
        RECT 1573.390 4.000 1576.690 4.280 ;
        RECT 1577.530 4.000 1580.830 4.280 ;
        RECT 1581.670 4.000 1584.970 4.280 ;
      LAYER met3 ;
        RECT 0.065 1584.760 1587.610 1591.365 ;
        RECT 0.065 1583.400 1587.065 1584.760 ;
        RECT 4.400 1583.360 1587.065 1583.400 ;
        RECT 4.400 1582.000 1587.610 1583.360 ;
        RECT 0.065 1549.400 1587.610 1582.000 ;
        RECT 0.065 1548.000 1587.065 1549.400 ;
        RECT 0.065 1545.320 1587.610 1548.000 ;
        RECT 4.400 1543.920 1587.610 1545.320 ;
        RECT 0.065 1513.360 1587.610 1543.920 ;
        RECT 0.065 1511.960 1587.065 1513.360 ;
        RECT 0.065 1507.240 1587.610 1511.960 ;
        RECT 4.400 1505.840 1587.610 1507.240 ;
        RECT 0.065 1478.000 1587.610 1505.840 ;
        RECT 0.065 1476.600 1587.065 1478.000 ;
        RECT 0.065 1469.160 1587.610 1476.600 ;
        RECT 4.400 1467.760 1587.610 1469.160 ;
        RECT 0.065 1442.640 1587.610 1467.760 ;
        RECT 0.065 1441.240 1587.065 1442.640 ;
        RECT 0.065 1431.080 1587.610 1441.240 ;
        RECT 4.400 1429.680 1587.610 1431.080 ;
        RECT 0.065 1406.600 1587.610 1429.680 ;
        RECT 0.065 1405.200 1587.065 1406.600 ;
        RECT 0.065 1393.000 1587.610 1405.200 ;
        RECT 4.400 1391.600 1587.610 1393.000 ;
        RECT 0.065 1371.240 1587.610 1391.600 ;
        RECT 0.065 1369.840 1587.065 1371.240 ;
        RECT 0.065 1354.920 1587.610 1369.840 ;
        RECT 4.400 1353.520 1587.610 1354.920 ;
        RECT 0.065 1335.880 1587.610 1353.520 ;
        RECT 0.065 1334.480 1587.065 1335.880 ;
        RECT 0.065 1316.840 1587.610 1334.480 ;
        RECT 4.400 1315.440 1587.610 1316.840 ;
        RECT 0.065 1299.840 1587.610 1315.440 ;
        RECT 0.065 1298.440 1587.065 1299.840 ;
        RECT 0.065 1278.760 1587.610 1298.440 ;
        RECT 4.400 1277.360 1587.610 1278.760 ;
        RECT 0.065 1264.480 1587.610 1277.360 ;
        RECT 0.065 1263.080 1587.065 1264.480 ;
        RECT 0.065 1240.680 1587.610 1263.080 ;
        RECT 4.400 1239.280 1587.610 1240.680 ;
        RECT 0.065 1229.120 1587.610 1239.280 ;
        RECT 0.065 1227.720 1587.065 1229.120 ;
        RECT 0.065 1201.920 1587.610 1227.720 ;
        RECT 4.400 1200.520 1587.610 1201.920 ;
        RECT 0.065 1193.080 1587.610 1200.520 ;
        RECT 0.065 1191.680 1587.065 1193.080 ;
        RECT 0.065 1163.840 1587.610 1191.680 ;
        RECT 4.400 1162.440 1587.610 1163.840 ;
        RECT 0.065 1157.720 1587.610 1162.440 ;
        RECT 0.065 1156.320 1587.065 1157.720 ;
        RECT 0.065 1125.760 1587.610 1156.320 ;
        RECT 4.400 1124.360 1587.610 1125.760 ;
        RECT 0.065 1122.360 1587.610 1124.360 ;
        RECT 0.065 1120.960 1587.065 1122.360 ;
        RECT 0.065 1087.680 1587.610 1120.960 ;
        RECT 4.400 1086.320 1587.610 1087.680 ;
        RECT 4.400 1086.280 1587.065 1086.320 ;
        RECT 0.065 1084.920 1587.065 1086.280 ;
        RECT 0.065 1050.960 1587.610 1084.920 ;
        RECT 0.065 1049.600 1587.065 1050.960 ;
        RECT 4.400 1049.560 1587.065 1049.600 ;
        RECT 4.400 1048.200 1587.610 1049.560 ;
        RECT 0.065 1014.920 1587.610 1048.200 ;
        RECT 0.065 1013.520 1587.065 1014.920 ;
        RECT 0.065 1011.520 1587.610 1013.520 ;
        RECT 4.400 1010.120 1587.610 1011.520 ;
        RECT 0.065 979.560 1587.610 1010.120 ;
        RECT 0.065 978.160 1587.065 979.560 ;
        RECT 0.065 973.440 1587.610 978.160 ;
        RECT 4.400 972.040 1587.610 973.440 ;
        RECT 0.065 944.200 1587.610 972.040 ;
        RECT 0.065 942.800 1587.065 944.200 ;
        RECT 0.065 935.360 1587.610 942.800 ;
        RECT 4.400 933.960 1587.610 935.360 ;
        RECT 0.065 908.160 1587.610 933.960 ;
        RECT 0.065 906.760 1587.065 908.160 ;
        RECT 0.065 897.280 1587.610 906.760 ;
        RECT 4.400 895.880 1587.610 897.280 ;
        RECT 0.065 872.800 1587.610 895.880 ;
        RECT 0.065 871.400 1587.065 872.800 ;
        RECT 0.065 859.200 1587.610 871.400 ;
        RECT 4.400 857.800 1587.610 859.200 ;
        RECT 0.065 837.440 1587.610 857.800 ;
        RECT 0.065 836.040 1587.065 837.440 ;
        RECT 0.065 821.120 1587.610 836.040 ;
        RECT 4.400 819.720 1587.610 821.120 ;
        RECT 0.065 801.400 1587.610 819.720 ;
        RECT 0.065 800.000 1587.065 801.400 ;
        RECT 0.065 782.360 1587.610 800.000 ;
        RECT 4.400 780.960 1587.610 782.360 ;
        RECT 0.065 766.040 1587.610 780.960 ;
        RECT 0.065 764.640 1587.065 766.040 ;
        RECT 0.065 744.280 1587.610 764.640 ;
        RECT 4.400 742.880 1587.610 744.280 ;
        RECT 0.065 730.680 1587.610 742.880 ;
        RECT 0.065 729.280 1587.065 730.680 ;
        RECT 0.065 706.200 1587.610 729.280 ;
        RECT 4.400 704.800 1587.610 706.200 ;
        RECT 0.065 694.640 1587.610 704.800 ;
        RECT 0.065 693.240 1587.065 694.640 ;
        RECT 0.065 668.120 1587.610 693.240 ;
        RECT 4.400 666.720 1587.610 668.120 ;
        RECT 0.065 659.280 1587.610 666.720 ;
        RECT 0.065 657.880 1587.065 659.280 ;
        RECT 0.065 630.040 1587.610 657.880 ;
        RECT 4.400 628.640 1587.610 630.040 ;
        RECT 0.065 623.920 1587.610 628.640 ;
        RECT 0.065 622.520 1587.065 623.920 ;
        RECT 0.065 591.960 1587.610 622.520 ;
        RECT 4.400 590.560 1587.610 591.960 ;
        RECT 0.065 587.880 1587.610 590.560 ;
        RECT 0.065 586.480 1587.065 587.880 ;
        RECT 0.065 553.880 1587.610 586.480 ;
        RECT 4.400 552.520 1587.610 553.880 ;
        RECT 4.400 552.480 1587.065 552.520 ;
        RECT 0.065 551.120 1587.065 552.480 ;
        RECT 0.065 516.480 1587.610 551.120 ;
        RECT 0.065 515.800 1587.065 516.480 ;
        RECT 4.400 515.080 1587.065 515.800 ;
        RECT 4.400 514.400 1587.610 515.080 ;
        RECT 0.065 481.120 1587.610 514.400 ;
        RECT 0.065 479.720 1587.065 481.120 ;
        RECT 0.065 477.720 1587.610 479.720 ;
        RECT 4.400 476.320 1587.610 477.720 ;
        RECT 0.065 445.760 1587.610 476.320 ;
        RECT 0.065 444.360 1587.065 445.760 ;
        RECT 0.065 439.640 1587.610 444.360 ;
        RECT 4.400 438.240 1587.610 439.640 ;
        RECT 0.065 409.720 1587.610 438.240 ;
        RECT 0.065 408.320 1587.065 409.720 ;
        RECT 0.065 400.880 1587.610 408.320 ;
        RECT 4.400 399.480 1587.610 400.880 ;
        RECT 0.065 374.360 1587.610 399.480 ;
        RECT 0.065 372.960 1587.065 374.360 ;
        RECT 0.065 362.800 1587.610 372.960 ;
        RECT 4.400 361.400 1587.610 362.800 ;
        RECT 0.065 339.000 1587.610 361.400 ;
        RECT 0.065 337.600 1587.065 339.000 ;
        RECT 0.065 324.720 1587.610 337.600 ;
        RECT 4.400 323.320 1587.610 324.720 ;
        RECT 0.065 302.960 1587.610 323.320 ;
        RECT 0.065 301.560 1587.065 302.960 ;
        RECT 0.065 286.640 1587.610 301.560 ;
        RECT 4.400 285.240 1587.610 286.640 ;
        RECT 0.065 267.600 1587.610 285.240 ;
        RECT 0.065 266.200 1587.065 267.600 ;
        RECT 0.065 248.560 1587.610 266.200 ;
        RECT 4.400 247.160 1587.610 248.560 ;
        RECT 0.065 232.240 1587.610 247.160 ;
        RECT 0.065 230.840 1587.065 232.240 ;
        RECT 0.065 210.480 1587.610 230.840 ;
        RECT 4.400 209.080 1587.610 210.480 ;
        RECT 0.065 196.200 1587.610 209.080 ;
        RECT 0.065 194.800 1587.065 196.200 ;
        RECT 0.065 172.400 1587.610 194.800 ;
        RECT 4.400 171.000 1587.610 172.400 ;
        RECT 0.065 160.840 1587.610 171.000 ;
        RECT 0.065 159.440 1587.065 160.840 ;
        RECT 0.065 134.320 1587.610 159.440 ;
        RECT 4.400 132.920 1587.610 134.320 ;
        RECT 0.065 125.480 1587.610 132.920 ;
        RECT 0.065 124.080 1587.065 125.480 ;
        RECT 0.065 96.240 1587.610 124.080 ;
        RECT 4.400 94.840 1587.610 96.240 ;
        RECT 0.065 89.440 1587.610 94.840 ;
        RECT 0.065 88.040 1587.065 89.440 ;
        RECT 0.065 58.160 1587.610 88.040 ;
        RECT 4.400 56.760 1587.610 58.160 ;
        RECT 0.065 54.080 1587.610 56.760 ;
        RECT 0.065 52.680 1587.065 54.080 ;
        RECT 0.065 20.080 1587.610 52.680 ;
        RECT 4.400 18.720 1587.610 20.080 ;
        RECT 4.400 18.680 1587.065 18.720 ;
        RECT 0.065 17.320 1587.065 18.680 ;
        RECT 0.065 10.715 1587.610 17.320 ;
      LAYER met4 ;
        RECT 11.335 10.640 20.640 1591.440 ;
        RECT 23.040 10.640 97.440 1591.440 ;
        RECT 99.840 10.640 1558.640 1591.440 ;
  END
END Ibtida_top_dffram_cv
END LIBRARY

