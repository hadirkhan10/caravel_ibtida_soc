magic
tech sky130A
magscale 1 2
timestamp 1607354317
<< obsli1 >>
rect 1104 2159 418876 497777
<< obsm1 >>
rect 1104 892 419414 497808
<< metal2 >>
rect 1858 499200 1914 500000
rect 4434 499200 4490 500000
rect 6826 499200 6882 500000
rect 9218 499200 9274 500000
rect 11794 499200 11850 500000
rect 14186 499200 14242 500000
rect 16762 499200 16818 500000
rect 19154 499200 19210 500000
rect 21730 499200 21786 500000
rect 24122 499200 24178 500000
rect 26514 499200 26570 500000
rect 29090 499200 29146 500000
rect 31482 499200 31538 500000
rect 34058 499200 34114 500000
rect 36450 499200 36506 500000
rect 39026 499200 39082 500000
rect 41418 499200 41474 500000
rect 43810 499200 43866 500000
rect 46386 499200 46442 500000
rect 48778 499200 48834 500000
rect 51354 499200 51410 500000
rect 53746 499200 53802 500000
rect 56322 499200 56378 500000
rect 58714 499200 58770 500000
rect 61106 499200 61162 500000
rect 63682 499200 63738 500000
rect 66074 499200 66130 500000
rect 68650 499200 68706 500000
rect 71042 499200 71098 500000
rect 73618 499200 73674 500000
rect 76010 499200 76066 500000
rect 78402 499200 78458 500000
rect 80978 499200 81034 500000
rect 83370 499200 83426 500000
rect 85946 499200 86002 500000
rect 88338 499200 88394 500000
rect 90914 499200 90970 500000
rect 93306 499200 93362 500000
rect 95698 499200 95754 500000
rect 98274 499200 98330 500000
rect 100666 499200 100722 500000
rect 103242 499200 103298 500000
rect 105634 499200 105690 500000
rect 108210 499200 108266 500000
rect 110602 499200 110658 500000
rect 112994 499200 113050 500000
rect 115570 499200 115626 500000
rect 117962 499200 118018 500000
rect 120538 499200 120594 500000
rect 122930 499200 122986 500000
rect 125506 499200 125562 500000
rect 127898 499200 127954 500000
rect 130290 499200 130346 500000
rect 132866 499200 132922 500000
rect 135258 499200 135314 500000
rect 137834 499200 137890 500000
rect 140226 499200 140282 500000
rect 142802 499200 142858 500000
rect 145194 499200 145250 500000
rect 147586 499200 147642 500000
rect 150162 499200 150218 500000
rect 152554 499200 152610 500000
rect 155130 499200 155186 500000
rect 157522 499200 157578 500000
rect 160098 499200 160154 500000
rect 162490 499200 162546 500000
rect 164882 499200 164938 500000
rect 167458 499200 167514 500000
rect 169850 499200 169906 500000
rect 172426 499200 172482 500000
rect 174818 499200 174874 500000
rect 177394 499200 177450 500000
rect 179786 499200 179842 500000
rect 182178 499200 182234 500000
rect 184754 499200 184810 500000
rect 187146 499200 187202 500000
rect 189722 499200 189778 500000
rect 192114 499200 192170 500000
rect 194690 499200 194746 500000
rect 197082 499200 197138 500000
rect 199474 499200 199530 500000
rect 202050 499200 202106 500000
rect 204442 499200 204498 500000
rect 207018 499200 207074 500000
rect 209410 499200 209466 500000
rect 211986 499200 212042 500000
rect 214378 499200 214434 500000
rect 216770 499200 216826 500000
rect 219346 499200 219402 500000
rect 221738 499200 221794 500000
rect 224314 499200 224370 500000
rect 226706 499200 226762 500000
rect 229282 499200 229338 500000
rect 231674 499200 231730 500000
rect 234066 499200 234122 500000
rect 236642 499200 236698 500000
rect 239034 499200 239090 500000
rect 241610 499200 241666 500000
rect 244002 499200 244058 500000
rect 246578 499200 246634 500000
rect 248970 499200 249026 500000
rect 251362 499200 251418 500000
rect 253938 499200 253994 500000
rect 256330 499200 256386 500000
rect 258906 499200 258962 500000
rect 261298 499200 261354 500000
rect 263874 499200 263930 500000
rect 266266 499200 266322 500000
rect 268658 499200 268714 500000
rect 271234 499200 271290 500000
rect 273626 499200 273682 500000
rect 276202 499200 276258 500000
rect 278594 499200 278650 500000
rect 281170 499200 281226 500000
rect 283562 499200 283618 500000
rect 285954 499200 286010 500000
rect 288530 499200 288586 500000
rect 290922 499200 290978 500000
rect 293498 499200 293554 500000
rect 295890 499200 295946 500000
rect 298466 499200 298522 500000
rect 300858 499200 300914 500000
rect 303250 499200 303306 500000
rect 305826 499200 305882 500000
rect 308218 499200 308274 500000
rect 310794 499200 310850 500000
rect 313186 499200 313242 500000
rect 315762 499200 315818 500000
rect 318154 499200 318210 500000
rect 320546 499200 320602 500000
rect 323122 499200 323178 500000
rect 325514 499200 325570 500000
rect 328090 499200 328146 500000
rect 330482 499200 330538 500000
rect 333058 499200 333114 500000
rect 335450 499200 335506 500000
rect 337842 499200 337898 500000
rect 340418 499200 340474 500000
rect 342810 499200 342866 500000
rect 345386 499200 345442 500000
rect 347778 499200 347834 500000
rect 350354 499200 350410 500000
rect 352746 499200 352802 500000
rect 355138 499200 355194 500000
rect 357714 499200 357770 500000
rect 360106 499200 360162 500000
rect 362682 499200 362738 500000
rect 365074 499200 365130 500000
rect 367650 499200 367706 500000
rect 370042 499200 370098 500000
rect 372434 499200 372490 500000
rect 375010 499200 375066 500000
rect 377402 499200 377458 500000
rect 379978 499200 380034 500000
rect 382370 499200 382426 500000
rect 384946 499200 385002 500000
rect 387338 499200 387394 500000
rect 389730 499200 389786 500000
rect 392306 499200 392362 500000
rect 394698 499200 394754 500000
rect 397274 499200 397330 500000
rect 399666 499200 399722 500000
rect 402242 499200 402298 500000
rect 404634 499200 404690 500000
rect 407026 499200 407082 500000
rect 409602 499200 409658 500000
rect 411994 499200 412050 500000
rect 414570 499200 414626 500000
rect 416962 499200 417018 500000
rect 419354 499200 419410 500000
rect 570 0 626 800
rect 2962 0 3018 800
rect 5354 0 5410 800
rect 7930 0 7986 800
rect 10322 0 10378 800
rect 12898 0 12954 800
rect 15290 0 15346 800
rect 17682 0 17738 800
rect 20258 0 20314 800
rect 22650 0 22706 800
rect 25226 0 25282 800
rect 27618 0 27674 800
rect 30194 0 30250 800
rect 32586 0 32642 800
rect 34978 0 35034 800
rect 37554 0 37610 800
rect 39946 0 40002 800
rect 42522 0 42578 800
rect 44914 0 44970 800
rect 47490 0 47546 800
rect 49882 0 49938 800
rect 52274 0 52330 800
rect 54850 0 54906 800
rect 57242 0 57298 800
rect 59818 0 59874 800
rect 62210 0 62266 800
rect 64786 0 64842 800
rect 67178 0 67234 800
rect 69570 0 69626 800
rect 72146 0 72202 800
rect 74538 0 74594 800
rect 77114 0 77170 800
rect 79506 0 79562 800
rect 82082 0 82138 800
rect 84474 0 84530 800
rect 86866 0 86922 800
rect 89442 0 89498 800
rect 91834 0 91890 800
rect 94410 0 94466 800
rect 96802 0 96858 800
rect 99378 0 99434 800
rect 101770 0 101826 800
rect 104162 0 104218 800
rect 106738 0 106794 800
rect 109130 0 109186 800
rect 111706 0 111762 800
rect 114098 0 114154 800
rect 116674 0 116730 800
rect 119066 0 119122 800
rect 121458 0 121514 800
rect 124034 0 124090 800
rect 126426 0 126482 800
rect 129002 0 129058 800
rect 131394 0 131450 800
rect 133970 0 134026 800
rect 136362 0 136418 800
rect 138754 0 138810 800
rect 141330 0 141386 800
rect 143722 0 143778 800
rect 146298 0 146354 800
rect 148690 0 148746 800
rect 151266 0 151322 800
rect 153658 0 153714 800
rect 156050 0 156106 800
rect 158626 0 158682 800
rect 161018 0 161074 800
rect 163594 0 163650 800
rect 165986 0 166042 800
rect 168562 0 168618 800
rect 170954 0 171010 800
rect 173346 0 173402 800
rect 175922 0 175978 800
rect 178314 0 178370 800
rect 180890 0 180946 800
rect 183282 0 183338 800
rect 185858 0 185914 800
rect 188250 0 188306 800
rect 190642 0 190698 800
rect 193218 0 193274 800
rect 195610 0 195666 800
rect 198186 0 198242 800
rect 200578 0 200634 800
rect 203154 0 203210 800
rect 205546 0 205602 800
rect 207938 0 207994 800
rect 210514 0 210570 800
rect 212906 0 212962 800
rect 215482 0 215538 800
rect 217874 0 217930 800
rect 220450 0 220506 800
rect 222842 0 222898 800
rect 225234 0 225290 800
rect 227810 0 227866 800
rect 230202 0 230258 800
rect 232778 0 232834 800
rect 235170 0 235226 800
rect 237746 0 237802 800
rect 240138 0 240194 800
rect 242530 0 242586 800
rect 245106 0 245162 800
rect 247498 0 247554 800
rect 250074 0 250130 800
rect 252466 0 252522 800
rect 255042 0 255098 800
rect 257434 0 257490 800
rect 259826 0 259882 800
rect 262402 0 262458 800
rect 264794 0 264850 800
rect 267370 0 267426 800
rect 269762 0 269818 800
rect 272338 0 272394 800
rect 274730 0 274786 800
rect 277122 0 277178 800
rect 279698 0 279754 800
rect 282090 0 282146 800
rect 284666 0 284722 800
rect 287058 0 287114 800
rect 289634 0 289690 800
rect 292026 0 292082 800
rect 294418 0 294474 800
rect 296994 0 297050 800
rect 299386 0 299442 800
rect 301962 0 302018 800
rect 304354 0 304410 800
rect 306930 0 306986 800
rect 309322 0 309378 800
rect 311714 0 311770 800
rect 314290 0 314346 800
rect 316682 0 316738 800
rect 319258 0 319314 800
rect 321650 0 321706 800
rect 324226 0 324282 800
rect 326618 0 326674 800
rect 329010 0 329066 800
rect 331586 0 331642 800
rect 333978 0 334034 800
rect 336554 0 336610 800
rect 338946 0 339002 800
rect 341522 0 341578 800
rect 343914 0 343970 800
rect 346306 0 346362 800
rect 348882 0 348938 800
rect 351274 0 351330 800
rect 353850 0 353906 800
rect 356242 0 356298 800
rect 358818 0 358874 800
rect 361210 0 361266 800
rect 363602 0 363658 800
rect 366178 0 366234 800
rect 368570 0 368626 800
rect 371146 0 371202 800
rect 373538 0 373594 800
rect 376114 0 376170 800
rect 378506 0 378562 800
rect 380898 0 380954 800
rect 383474 0 383530 800
rect 385866 0 385922 800
rect 388442 0 388498 800
rect 390834 0 390890 800
rect 393410 0 393466 800
rect 395802 0 395858 800
rect 398194 0 398250 800
rect 400770 0 400826 800
rect 403162 0 403218 800
rect 405738 0 405794 800
rect 408130 0 408186 800
rect 410706 0 410762 800
rect 413098 0 413154 800
rect 415490 0 415546 800
rect 418066 0 418122 800
<< obsm2 >>
rect 1768 499144 1802 499202
rect 1970 499144 4378 499202
rect 4546 499144 6770 499202
rect 6938 499144 9162 499202
rect 9330 499144 11738 499202
rect 11906 499144 14130 499202
rect 14298 499144 16706 499202
rect 16874 499144 19098 499202
rect 19266 499144 21674 499202
rect 21842 499144 24066 499202
rect 24234 499144 26458 499202
rect 26626 499144 29034 499202
rect 29202 499144 31426 499202
rect 31594 499144 34002 499202
rect 34170 499144 36394 499202
rect 36562 499144 38970 499202
rect 39138 499144 41362 499202
rect 41530 499144 43754 499202
rect 43922 499144 46330 499202
rect 46498 499144 48722 499202
rect 48890 499144 51298 499202
rect 51466 499144 53690 499202
rect 53858 499144 56266 499202
rect 56434 499144 58658 499202
rect 58826 499144 61050 499202
rect 61218 499144 63626 499202
rect 63794 499144 66018 499202
rect 66186 499144 68594 499202
rect 68762 499144 70986 499202
rect 71154 499144 73562 499202
rect 73730 499144 75954 499202
rect 76122 499144 78346 499202
rect 78514 499144 80922 499202
rect 81090 499144 83314 499202
rect 83482 499144 85890 499202
rect 86058 499144 88282 499202
rect 88450 499144 90858 499202
rect 91026 499144 93250 499202
rect 93418 499144 95642 499202
rect 95810 499144 98218 499202
rect 98386 499144 100610 499202
rect 100778 499144 103186 499202
rect 103354 499144 105578 499202
rect 105746 499144 108154 499202
rect 108322 499144 110546 499202
rect 110714 499144 112938 499202
rect 113106 499144 115514 499202
rect 115682 499144 117906 499202
rect 118074 499144 120482 499202
rect 120650 499144 122874 499202
rect 123042 499144 125450 499202
rect 125618 499144 127842 499202
rect 128010 499144 130234 499202
rect 130402 499144 132810 499202
rect 132978 499144 135202 499202
rect 135370 499144 137778 499202
rect 137946 499144 140170 499202
rect 140338 499144 142746 499202
rect 142914 499144 145138 499202
rect 145306 499144 147530 499202
rect 147698 499144 150106 499202
rect 150274 499144 152498 499202
rect 152666 499144 155074 499202
rect 155242 499144 157466 499202
rect 157634 499144 160042 499202
rect 160210 499144 162434 499202
rect 162602 499144 164826 499202
rect 164994 499144 167402 499202
rect 167570 499144 169794 499202
rect 169962 499144 172370 499202
rect 172538 499144 174762 499202
rect 174930 499144 177338 499202
rect 177506 499144 179730 499202
rect 179898 499144 182122 499202
rect 182290 499144 184698 499202
rect 184866 499144 187090 499202
rect 187258 499144 189666 499202
rect 189834 499144 192058 499202
rect 192226 499144 194634 499202
rect 194802 499144 197026 499202
rect 197194 499144 199418 499202
rect 199586 499144 201994 499202
rect 202162 499144 204386 499202
rect 204554 499144 206962 499202
rect 207130 499144 209354 499202
rect 209522 499144 211930 499202
rect 212098 499144 214322 499202
rect 214490 499144 216714 499202
rect 216882 499144 219290 499202
rect 219458 499144 221682 499202
rect 221850 499144 224258 499202
rect 224426 499144 226650 499202
rect 226818 499144 229226 499202
rect 229394 499144 231618 499202
rect 231786 499144 234010 499202
rect 234178 499144 236586 499202
rect 236754 499144 238978 499202
rect 239146 499144 241554 499202
rect 241722 499144 243946 499202
rect 244114 499144 246522 499202
rect 246690 499144 248914 499202
rect 249082 499144 251306 499202
rect 251474 499144 253882 499202
rect 254050 499144 256274 499202
rect 256442 499144 258850 499202
rect 259018 499144 261242 499202
rect 261410 499144 263818 499202
rect 263986 499144 266210 499202
rect 266378 499144 268602 499202
rect 268770 499144 271178 499202
rect 271346 499144 273570 499202
rect 273738 499144 276146 499202
rect 276314 499144 278538 499202
rect 278706 499144 281114 499202
rect 281282 499144 283506 499202
rect 283674 499144 285898 499202
rect 286066 499144 288474 499202
rect 288642 499144 290866 499202
rect 291034 499144 293442 499202
rect 293610 499144 295834 499202
rect 296002 499144 298410 499202
rect 298578 499144 300802 499202
rect 300970 499144 303194 499202
rect 303362 499144 305770 499202
rect 305938 499144 308162 499202
rect 308330 499144 310738 499202
rect 310906 499144 313130 499202
rect 313298 499144 315706 499202
rect 315874 499144 318098 499202
rect 318266 499144 320490 499202
rect 320658 499144 323066 499202
rect 323234 499144 325458 499202
rect 325626 499144 328034 499202
rect 328202 499144 330426 499202
rect 330594 499144 333002 499202
rect 333170 499144 335394 499202
rect 335562 499144 337786 499202
rect 337954 499144 340362 499202
rect 340530 499144 342754 499202
rect 342922 499144 345330 499202
rect 345498 499144 347722 499202
rect 347890 499144 350298 499202
rect 350466 499144 352690 499202
rect 352858 499144 355082 499202
rect 355250 499144 357658 499202
rect 357826 499144 360050 499202
rect 360218 499144 362626 499202
rect 362794 499144 365018 499202
rect 365186 499144 367594 499202
rect 367762 499144 369986 499202
rect 370154 499144 372378 499202
rect 372546 499144 374954 499202
rect 375122 499144 377346 499202
rect 377514 499144 379922 499202
rect 380090 499144 382314 499202
rect 382482 499144 384890 499202
rect 385058 499144 387282 499202
rect 387450 499144 389674 499202
rect 389842 499144 392250 499202
rect 392418 499144 394642 499202
rect 394810 499144 397218 499202
rect 397386 499144 399610 499202
rect 399778 499144 402186 499202
rect 402354 499144 404578 499202
rect 404746 499144 406970 499202
rect 407138 499144 409546 499202
rect 409714 499144 411938 499202
rect 412106 499144 414514 499202
rect 414682 499144 416906 499202
rect 417074 499144 419298 499202
rect 1768 856 419408 499144
rect 1768 800 2906 856
rect 3074 800 5298 856
rect 5466 800 7874 856
rect 8042 800 10266 856
rect 10434 800 12842 856
rect 13010 800 15234 856
rect 15402 800 17626 856
rect 17794 800 20202 856
rect 20370 800 22594 856
rect 22762 800 25170 856
rect 25338 800 27562 856
rect 27730 800 30138 856
rect 30306 800 32530 856
rect 32698 800 34922 856
rect 35090 800 37498 856
rect 37666 800 39890 856
rect 40058 800 42466 856
rect 42634 800 44858 856
rect 45026 800 47434 856
rect 47602 800 49826 856
rect 49994 800 52218 856
rect 52386 800 54794 856
rect 54962 800 57186 856
rect 57354 800 59762 856
rect 59930 800 62154 856
rect 62322 800 64730 856
rect 64898 800 67122 856
rect 67290 800 69514 856
rect 69682 800 72090 856
rect 72258 800 74482 856
rect 74650 800 77058 856
rect 77226 800 79450 856
rect 79618 800 82026 856
rect 82194 800 84418 856
rect 84586 800 86810 856
rect 86978 800 89386 856
rect 89554 800 91778 856
rect 91946 800 94354 856
rect 94522 800 96746 856
rect 96914 800 99322 856
rect 99490 800 101714 856
rect 101882 800 104106 856
rect 104274 800 106682 856
rect 106850 800 109074 856
rect 109242 800 111650 856
rect 111818 800 114042 856
rect 114210 800 116618 856
rect 116786 800 119010 856
rect 119178 800 121402 856
rect 121570 800 123978 856
rect 124146 800 126370 856
rect 126538 800 128946 856
rect 129114 800 131338 856
rect 131506 800 133914 856
rect 134082 800 136306 856
rect 136474 800 138698 856
rect 138866 800 141274 856
rect 141442 800 143666 856
rect 143834 800 146242 856
rect 146410 800 148634 856
rect 148802 800 151210 856
rect 151378 800 153602 856
rect 153770 800 155994 856
rect 156162 800 158570 856
rect 158738 800 160962 856
rect 161130 800 163538 856
rect 163706 800 165930 856
rect 166098 800 168506 856
rect 168674 800 170898 856
rect 171066 800 173290 856
rect 173458 800 175866 856
rect 176034 800 178258 856
rect 178426 800 180834 856
rect 181002 800 183226 856
rect 183394 800 185802 856
rect 185970 800 188194 856
rect 188362 800 190586 856
rect 190754 800 193162 856
rect 193330 800 195554 856
rect 195722 800 198130 856
rect 198298 800 200522 856
rect 200690 800 203098 856
rect 203266 800 205490 856
rect 205658 800 207882 856
rect 208050 800 210458 856
rect 210626 800 212850 856
rect 213018 800 215426 856
rect 215594 800 217818 856
rect 217986 800 220394 856
rect 220562 800 222786 856
rect 222954 800 225178 856
rect 225346 800 227754 856
rect 227922 800 230146 856
rect 230314 800 232722 856
rect 232890 800 235114 856
rect 235282 800 237690 856
rect 237858 800 240082 856
rect 240250 800 242474 856
rect 242642 800 245050 856
rect 245218 800 247442 856
rect 247610 800 250018 856
rect 250186 800 252410 856
rect 252578 800 254986 856
rect 255154 800 257378 856
rect 257546 800 259770 856
rect 259938 800 262346 856
rect 262514 800 264738 856
rect 264906 800 267314 856
rect 267482 800 269706 856
rect 269874 800 272282 856
rect 272450 800 274674 856
rect 274842 800 277066 856
rect 277234 800 279642 856
rect 279810 800 282034 856
rect 282202 800 284610 856
rect 284778 800 287002 856
rect 287170 800 289578 856
rect 289746 800 291970 856
rect 292138 800 294362 856
rect 294530 800 296938 856
rect 297106 800 299330 856
rect 299498 800 301906 856
rect 302074 800 304298 856
rect 304466 800 306874 856
rect 307042 800 309266 856
rect 309434 800 311658 856
rect 311826 800 314234 856
rect 314402 800 316626 856
rect 316794 800 319202 856
rect 319370 800 321594 856
rect 321762 800 324170 856
rect 324338 800 326562 856
rect 326730 800 328954 856
rect 329122 800 331530 856
rect 331698 800 333922 856
rect 334090 800 336498 856
rect 336666 800 338890 856
rect 339058 800 341466 856
rect 341634 800 343858 856
rect 344026 800 346250 856
rect 346418 800 348826 856
rect 348994 800 351218 856
rect 351386 800 353794 856
rect 353962 800 356186 856
rect 356354 800 358762 856
rect 358930 800 361154 856
rect 361322 800 363546 856
rect 363714 800 366122 856
rect 366290 800 368514 856
rect 368682 800 371090 856
rect 371258 800 373482 856
rect 373650 800 376058 856
rect 376226 800 378450 856
rect 378618 800 380842 856
rect 381010 800 383418 856
rect 383586 800 385810 856
rect 385978 800 388386 856
rect 388554 800 390778 856
rect 390946 800 393354 856
rect 393522 800 395746 856
rect 395914 800 398138 856
rect 398306 800 400714 856
rect 400882 800 403106 856
rect 403274 800 405682 856
rect 405850 800 408074 856
rect 408242 800 410650 856
rect 410818 800 413042 856
rect 413210 800 415434 856
rect 415602 800 418010 856
rect 418178 800 419408 856
<< metal3 >>
rect 0 497496 800 497616
rect 419200 495320 420000 495440
rect 0 493688 800 493808
rect 419200 491784 420000 491904
rect 0 490152 800 490272
rect 419200 487976 420000 488096
rect 0 486344 800 486464
rect 419200 484440 420000 484560
rect 0 482808 800 482928
rect 419200 480632 420000 480752
rect 0 479272 800 479392
rect 419200 477096 420000 477216
rect 0 475464 800 475584
rect 419200 473560 420000 473680
rect 0 471928 800 472048
rect 419200 469752 420000 469872
rect 0 468120 800 468240
rect 419200 466216 420000 466336
rect 0 464584 800 464704
rect 419200 462408 420000 462528
rect 0 460776 800 460896
rect 419200 458872 420000 458992
rect 0 457240 800 457360
rect 419200 455064 420000 455184
rect 0 453704 800 453824
rect 419200 451528 420000 451648
rect 0 449896 800 450016
rect 419200 447992 420000 448112
rect 0 446360 800 446480
rect 419200 444184 420000 444304
rect 0 442552 800 442672
rect 419200 440648 420000 440768
rect 0 439016 800 439136
rect 419200 436840 420000 436960
rect 0 435208 800 435328
rect 419200 433304 420000 433424
rect 0 431672 800 431792
rect 419200 429496 420000 429616
rect 0 428136 800 428256
rect 419200 425960 420000 426080
rect 0 424328 800 424448
rect 419200 422424 420000 422544
rect 0 420792 800 420912
rect 419200 418616 420000 418736
rect 0 416984 800 417104
rect 419200 415080 420000 415200
rect 0 413448 800 413568
rect 419200 411272 420000 411392
rect 0 409640 800 409760
rect 419200 407736 420000 407856
rect 0 406104 800 406224
rect 419200 403928 420000 404048
rect 0 402568 800 402688
rect 419200 400392 420000 400512
rect 0 398760 800 398880
rect 419200 396856 420000 396976
rect 0 395224 800 395344
rect 419200 393048 420000 393168
rect 0 391416 800 391536
rect 419200 389512 420000 389632
rect 0 387880 800 388000
rect 419200 385704 420000 385824
rect 0 384072 800 384192
rect 419200 382168 420000 382288
rect 0 380536 800 380656
rect 419200 378360 420000 378480
rect 0 377000 800 377120
rect 419200 374824 420000 374944
rect 0 373192 800 373312
rect 419200 371288 420000 371408
rect 0 369656 800 369776
rect 419200 367480 420000 367600
rect 0 365848 800 365968
rect 419200 363944 420000 364064
rect 0 362312 800 362432
rect 419200 360136 420000 360256
rect 0 358504 800 358624
rect 419200 356600 420000 356720
rect 0 354968 800 355088
rect 419200 352792 420000 352912
rect 0 351432 800 351552
rect 419200 349256 420000 349376
rect 0 347624 800 347744
rect 419200 345720 420000 345840
rect 0 344088 800 344208
rect 419200 341912 420000 342032
rect 0 340280 800 340400
rect 419200 338376 420000 338496
rect 0 336744 800 336864
rect 419200 334568 420000 334688
rect 0 332936 800 333056
rect 419200 331032 420000 331152
rect 0 329400 800 329520
rect 419200 327224 420000 327344
rect 0 325864 800 325984
rect 419200 323688 420000 323808
rect 0 322056 800 322176
rect 419200 320152 420000 320272
rect 0 318520 800 318640
rect 419200 316344 420000 316464
rect 0 314712 800 314832
rect 419200 312808 420000 312928
rect 0 311176 800 311296
rect 419200 309000 420000 309120
rect 0 307368 800 307488
rect 419200 305464 420000 305584
rect 0 303832 800 303952
rect 419200 301656 420000 301776
rect 0 300296 800 300416
rect 419200 298120 420000 298240
rect 0 296488 800 296608
rect 419200 294584 420000 294704
rect 0 292952 800 293072
rect 419200 290776 420000 290896
rect 0 289144 800 289264
rect 419200 287240 420000 287360
rect 0 285608 800 285728
rect 419200 283432 420000 283552
rect 0 281800 800 281920
rect 419200 279896 420000 280016
rect 0 278264 800 278384
rect 419200 276088 420000 276208
rect 0 274728 800 274848
rect 419200 272552 420000 272672
rect 0 270920 800 271040
rect 419200 269016 420000 269136
rect 0 267384 800 267504
rect 419200 265208 420000 265328
rect 0 263576 800 263696
rect 419200 261672 420000 261792
rect 0 260040 800 260160
rect 419200 257864 420000 257984
rect 0 256232 800 256352
rect 419200 254328 420000 254448
rect 0 252696 800 252816
rect 419200 250520 420000 250640
rect 0 249160 800 249280
rect 419200 246984 420000 247104
rect 0 245352 800 245472
rect 419200 243448 420000 243568
rect 0 241816 800 241936
rect 419200 239640 420000 239760
rect 0 238008 800 238128
rect 419200 236104 420000 236224
rect 0 234472 800 234592
rect 419200 232296 420000 232416
rect 0 230664 800 230784
rect 419200 228760 420000 228880
rect 0 227128 800 227248
rect 419200 224952 420000 225072
rect 0 223592 800 223712
rect 419200 221416 420000 221536
rect 0 219784 800 219904
rect 419200 217880 420000 218000
rect 0 216248 800 216368
rect 419200 214072 420000 214192
rect 0 212440 800 212560
rect 419200 210536 420000 210656
rect 0 208904 800 209024
rect 419200 206728 420000 206848
rect 0 205096 800 205216
rect 419200 203192 420000 203312
rect 0 201560 800 201680
rect 419200 199384 420000 199504
rect 0 198024 800 198144
rect 419200 195848 420000 195968
rect 0 194216 800 194336
rect 419200 192312 420000 192432
rect 0 190680 800 190800
rect 419200 188504 420000 188624
rect 0 186872 800 186992
rect 419200 184968 420000 185088
rect 0 183336 800 183456
rect 419200 181160 420000 181280
rect 0 179528 800 179648
rect 419200 177624 420000 177744
rect 0 175992 800 176112
rect 419200 173816 420000 173936
rect 0 172456 800 172576
rect 419200 170280 420000 170400
rect 0 168648 800 168768
rect 419200 166744 420000 166864
rect 0 165112 800 165232
rect 419200 162936 420000 163056
rect 0 161304 800 161424
rect 419200 159400 420000 159520
rect 0 157768 800 157888
rect 419200 155592 420000 155712
rect 0 153960 800 154080
rect 419200 152056 420000 152176
rect 0 150424 800 150544
rect 419200 148248 420000 148368
rect 0 146888 800 147008
rect 419200 144712 420000 144832
rect 0 143080 800 143200
rect 419200 141176 420000 141296
rect 0 139544 800 139664
rect 419200 137368 420000 137488
rect 0 135736 800 135856
rect 419200 133832 420000 133952
rect 0 132200 800 132320
rect 419200 130024 420000 130144
rect 0 128392 800 128512
rect 419200 126488 420000 126608
rect 0 124856 800 124976
rect 419200 122680 420000 122800
rect 0 121320 800 121440
rect 419200 119144 420000 119264
rect 0 117512 800 117632
rect 419200 115608 420000 115728
rect 0 113976 800 114096
rect 419200 111800 420000 111920
rect 0 110168 800 110288
rect 419200 108264 420000 108384
rect 0 106632 800 106752
rect 419200 104456 420000 104576
rect 0 102824 800 102944
rect 419200 100920 420000 101040
rect 0 99288 800 99408
rect 419200 97112 420000 97232
rect 0 95752 800 95872
rect 419200 93576 420000 93696
rect 0 91944 800 92064
rect 419200 90040 420000 90160
rect 0 88408 800 88528
rect 419200 86232 420000 86352
rect 0 84600 800 84720
rect 419200 82696 420000 82816
rect 0 81064 800 81184
rect 419200 78888 420000 79008
rect 0 77256 800 77376
rect 419200 75352 420000 75472
rect 0 73720 800 73840
rect 419200 71544 420000 71664
rect 0 70184 800 70304
rect 419200 68008 420000 68128
rect 0 66376 800 66496
rect 419200 64472 420000 64592
rect 0 62840 800 62960
rect 419200 60664 420000 60784
rect 0 59032 800 59152
rect 419200 57128 420000 57248
rect 0 55496 800 55616
rect 419200 53320 420000 53440
rect 0 51688 800 51808
rect 419200 49784 420000 49904
rect 0 48152 800 48272
rect 419200 45976 420000 46096
rect 0 44616 800 44736
rect 419200 42440 420000 42560
rect 0 40808 800 40928
rect 419200 38904 420000 39024
rect 0 37272 800 37392
rect 419200 35096 420000 35216
rect 0 33464 800 33584
rect 419200 31560 420000 31680
rect 0 29928 800 30048
rect 419200 27752 420000 27872
rect 0 26120 800 26240
rect 419200 24216 420000 24336
rect 0 22584 800 22704
rect 419200 20408 420000 20528
rect 0 19048 800 19168
rect 419200 16872 420000 16992
rect 0 15240 800 15360
rect 419200 13336 420000 13456
rect 0 11704 800 11824
rect 419200 9528 420000 9648
rect 0 7896 800 8016
rect 419200 5992 420000 6112
rect 0 4360 800 4480
rect 419200 2184 420000 2304
<< obsm3 >>
rect 800 497696 419200 497793
rect 880 497416 419200 497696
rect 800 495520 419200 497416
rect 800 495240 419120 495520
rect 800 493888 419200 495240
rect 880 493608 419200 493888
rect 800 491984 419200 493608
rect 800 491704 419120 491984
rect 800 490352 419200 491704
rect 880 490072 419200 490352
rect 800 488176 419200 490072
rect 800 487896 419120 488176
rect 800 486544 419200 487896
rect 880 486264 419200 486544
rect 800 484640 419200 486264
rect 800 484360 419120 484640
rect 800 483008 419200 484360
rect 880 482728 419200 483008
rect 800 480832 419200 482728
rect 800 480552 419120 480832
rect 800 479472 419200 480552
rect 880 479192 419200 479472
rect 800 477296 419200 479192
rect 800 477016 419120 477296
rect 800 475664 419200 477016
rect 880 475384 419200 475664
rect 800 473760 419200 475384
rect 800 473480 419120 473760
rect 800 472128 419200 473480
rect 880 471848 419200 472128
rect 800 469952 419200 471848
rect 800 469672 419120 469952
rect 800 468320 419200 469672
rect 880 468040 419200 468320
rect 800 466416 419200 468040
rect 800 466136 419120 466416
rect 800 464784 419200 466136
rect 880 464504 419200 464784
rect 800 462608 419200 464504
rect 800 462328 419120 462608
rect 800 460976 419200 462328
rect 880 460696 419200 460976
rect 800 459072 419200 460696
rect 800 458792 419120 459072
rect 800 457440 419200 458792
rect 880 457160 419200 457440
rect 800 455264 419200 457160
rect 800 454984 419120 455264
rect 800 453904 419200 454984
rect 880 453624 419200 453904
rect 800 451728 419200 453624
rect 800 451448 419120 451728
rect 800 450096 419200 451448
rect 880 449816 419200 450096
rect 800 448192 419200 449816
rect 800 447912 419120 448192
rect 800 446560 419200 447912
rect 880 446280 419200 446560
rect 800 444384 419200 446280
rect 800 444104 419120 444384
rect 800 442752 419200 444104
rect 880 442472 419200 442752
rect 800 440848 419200 442472
rect 800 440568 419120 440848
rect 800 439216 419200 440568
rect 880 438936 419200 439216
rect 800 437040 419200 438936
rect 800 436760 419120 437040
rect 800 435408 419200 436760
rect 880 435128 419200 435408
rect 800 433504 419200 435128
rect 800 433224 419120 433504
rect 800 431872 419200 433224
rect 880 431592 419200 431872
rect 800 429696 419200 431592
rect 800 429416 419120 429696
rect 800 428336 419200 429416
rect 880 428056 419200 428336
rect 800 426160 419200 428056
rect 800 425880 419120 426160
rect 800 424528 419200 425880
rect 880 424248 419200 424528
rect 800 422624 419200 424248
rect 800 422344 419120 422624
rect 800 420992 419200 422344
rect 880 420712 419200 420992
rect 800 418816 419200 420712
rect 800 418536 419120 418816
rect 800 417184 419200 418536
rect 880 416904 419200 417184
rect 800 415280 419200 416904
rect 800 415000 419120 415280
rect 800 413648 419200 415000
rect 880 413368 419200 413648
rect 800 411472 419200 413368
rect 800 411192 419120 411472
rect 800 409840 419200 411192
rect 880 409560 419200 409840
rect 800 407936 419200 409560
rect 800 407656 419120 407936
rect 800 406304 419200 407656
rect 880 406024 419200 406304
rect 800 404128 419200 406024
rect 800 403848 419120 404128
rect 800 402768 419200 403848
rect 880 402488 419200 402768
rect 800 400592 419200 402488
rect 800 400312 419120 400592
rect 800 398960 419200 400312
rect 880 398680 419200 398960
rect 800 397056 419200 398680
rect 800 396776 419120 397056
rect 800 395424 419200 396776
rect 880 395144 419200 395424
rect 800 393248 419200 395144
rect 800 392968 419120 393248
rect 800 391616 419200 392968
rect 880 391336 419200 391616
rect 800 389712 419200 391336
rect 800 389432 419120 389712
rect 800 388080 419200 389432
rect 880 387800 419200 388080
rect 800 385904 419200 387800
rect 800 385624 419120 385904
rect 800 384272 419200 385624
rect 880 383992 419200 384272
rect 800 382368 419200 383992
rect 800 382088 419120 382368
rect 800 380736 419200 382088
rect 880 380456 419200 380736
rect 800 378560 419200 380456
rect 800 378280 419120 378560
rect 800 377200 419200 378280
rect 880 376920 419200 377200
rect 800 375024 419200 376920
rect 800 374744 419120 375024
rect 800 373392 419200 374744
rect 880 373112 419200 373392
rect 800 371488 419200 373112
rect 800 371208 419120 371488
rect 800 369856 419200 371208
rect 880 369576 419200 369856
rect 800 367680 419200 369576
rect 800 367400 419120 367680
rect 800 366048 419200 367400
rect 880 365768 419200 366048
rect 800 364144 419200 365768
rect 800 363864 419120 364144
rect 800 362512 419200 363864
rect 880 362232 419200 362512
rect 800 360336 419200 362232
rect 800 360056 419120 360336
rect 800 358704 419200 360056
rect 880 358424 419200 358704
rect 800 356800 419200 358424
rect 800 356520 419120 356800
rect 800 355168 419200 356520
rect 880 354888 419200 355168
rect 800 352992 419200 354888
rect 800 352712 419120 352992
rect 800 351632 419200 352712
rect 880 351352 419200 351632
rect 800 349456 419200 351352
rect 800 349176 419120 349456
rect 800 347824 419200 349176
rect 880 347544 419200 347824
rect 800 345920 419200 347544
rect 800 345640 419120 345920
rect 800 344288 419200 345640
rect 880 344008 419200 344288
rect 800 342112 419200 344008
rect 800 341832 419120 342112
rect 800 340480 419200 341832
rect 880 340200 419200 340480
rect 800 338576 419200 340200
rect 800 338296 419120 338576
rect 800 336944 419200 338296
rect 880 336664 419200 336944
rect 800 334768 419200 336664
rect 800 334488 419120 334768
rect 800 333136 419200 334488
rect 880 332856 419200 333136
rect 800 331232 419200 332856
rect 800 330952 419120 331232
rect 800 329600 419200 330952
rect 880 329320 419200 329600
rect 800 327424 419200 329320
rect 800 327144 419120 327424
rect 800 326064 419200 327144
rect 880 325784 419200 326064
rect 800 323888 419200 325784
rect 800 323608 419120 323888
rect 800 322256 419200 323608
rect 880 321976 419200 322256
rect 800 320352 419200 321976
rect 800 320072 419120 320352
rect 800 318720 419200 320072
rect 880 318440 419200 318720
rect 800 316544 419200 318440
rect 800 316264 419120 316544
rect 800 314912 419200 316264
rect 880 314632 419200 314912
rect 800 313008 419200 314632
rect 800 312728 419120 313008
rect 800 311376 419200 312728
rect 880 311096 419200 311376
rect 800 309200 419200 311096
rect 800 308920 419120 309200
rect 800 307568 419200 308920
rect 880 307288 419200 307568
rect 800 305664 419200 307288
rect 800 305384 419120 305664
rect 800 304032 419200 305384
rect 880 303752 419200 304032
rect 800 301856 419200 303752
rect 800 301576 419120 301856
rect 800 300496 419200 301576
rect 880 300216 419200 300496
rect 800 298320 419200 300216
rect 800 298040 419120 298320
rect 800 296688 419200 298040
rect 880 296408 419200 296688
rect 800 294784 419200 296408
rect 800 294504 419120 294784
rect 800 293152 419200 294504
rect 880 292872 419200 293152
rect 800 290976 419200 292872
rect 800 290696 419120 290976
rect 800 289344 419200 290696
rect 880 289064 419200 289344
rect 800 287440 419200 289064
rect 800 287160 419120 287440
rect 800 285808 419200 287160
rect 880 285528 419200 285808
rect 800 283632 419200 285528
rect 800 283352 419120 283632
rect 800 282000 419200 283352
rect 880 281720 419200 282000
rect 800 280096 419200 281720
rect 800 279816 419120 280096
rect 800 278464 419200 279816
rect 880 278184 419200 278464
rect 800 276288 419200 278184
rect 800 276008 419120 276288
rect 800 274928 419200 276008
rect 880 274648 419200 274928
rect 800 272752 419200 274648
rect 800 272472 419120 272752
rect 800 271120 419200 272472
rect 880 270840 419200 271120
rect 800 269216 419200 270840
rect 800 268936 419120 269216
rect 800 267584 419200 268936
rect 880 267304 419200 267584
rect 800 265408 419200 267304
rect 800 265128 419120 265408
rect 800 263776 419200 265128
rect 880 263496 419200 263776
rect 800 261872 419200 263496
rect 800 261592 419120 261872
rect 800 260240 419200 261592
rect 880 259960 419200 260240
rect 800 258064 419200 259960
rect 800 257784 419120 258064
rect 800 256432 419200 257784
rect 880 256152 419200 256432
rect 800 254528 419200 256152
rect 800 254248 419120 254528
rect 800 252896 419200 254248
rect 880 252616 419200 252896
rect 800 250720 419200 252616
rect 800 250440 419120 250720
rect 800 249360 419200 250440
rect 880 249080 419200 249360
rect 800 247184 419200 249080
rect 800 246904 419120 247184
rect 800 245552 419200 246904
rect 880 245272 419200 245552
rect 800 243648 419200 245272
rect 800 243368 419120 243648
rect 800 242016 419200 243368
rect 880 241736 419200 242016
rect 800 239840 419200 241736
rect 800 239560 419120 239840
rect 800 238208 419200 239560
rect 880 237928 419200 238208
rect 800 236304 419200 237928
rect 800 236024 419120 236304
rect 800 234672 419200 236024
rect 880 234392 419200 234672
rect 800 232496 419200 234392
rect 800 232216 419120 232496
rect 800 230864 419200 232216
rect 880 230584 419200 230864
rect 800 228960 419200 230584
rect 800 228680 419120 228960
rect 800 227328 419200 228680
rect 880 227048 419200 227328
rect 800 225152 419200 227048
rect 800 224872 419120 225152
rect 800 223792 419200 224872
rect 880 223512 419200 223792
rect 800 221616 419200 223512
rect 800 221336 419120 221616
rect 800 219984 419200 221336
rect 880 219704 419200 219984
rect 800 218080 419200 219704
rect 800 217800 419120 218080
rect 800 216448 419200 217800
rect 880 216168 419200 216448
rect 800 214272 419200 216168
rect 800 213992 419120 214272
rect 800 212640 419200 213992
rect 880 212360 419200 212640
rect 800 210736 419200 212360
rect 800 210456 419120 210736
rect 800 209104 419200 210456
rect 880 208824 419200 209104
rect 800 206928 419200 208824
rect 800 206648 419120 206928
rect 800 205296 419200 206648
rect 880 205016 419200 205296
rect 800 203392 419200 205016
rect 800 203112 419120 203392
rect 800 201760 419200 203112
rect 880 201480 419200 201760
rect 800 199584 419200 201480
rect 800 199304 419120 199584
rect 800 198224 419200 199304
rect 880 197944 419200 198224
rect 800 196048 419200 197944
rect 800 195768 419120 196048
rect 800 194416 419200 195768
rect 880 194136 419200 194416
rect 800 192512 419200 194136
rect 800 192232 419120 192512
rect 800 190880 419200 192232
rect 880 190600 419200 190880
rect 800 188704 419200 190600
rect 800 188424 419120 188704
rect 800 187072 419200 188424
rect 880 186792 419200 187072
rect 800 185168 419200 186792
rect 800 184888 419120 185168
rect 800 183536 419200 184888
rect 880 183256 419200 183536
rect 800 181360 419200 183256
rect 800 181080 419120 181360
rect 800 179728 419200 181080
rect 880 179448 419200 179728
rect 800 177824 419200 179448
rect 800 177544 419120 177824
rect 800 176192 419200 177544
rect 880 175912 419200 176192
rect 800 174016 419200 175912
rect 800 173736 419120 174016
rect 800 172656 419200 173736
rect 880 172376 419200 172656
rect 800 170480 419200 172376
rect 800 170200 419120 170480
rect 800 168848 419200 170200
rect 880 168568 419200 168848
rect 800 166944 419200 168568
rect 800 166664 419120 166944
rect 800 165312 419200 166664
rect 880 165032 419200 165312
rect 800 163136 419200 165032
rect 800 162856 419120 163136
rect 800 161504 419200 162856
rect 880 161224 419200 161504
rect 800 159600 419200 161224
rect 800 159320 419120 159600
rect 800 157968 419200 159320
rect 880 157688 419200 157968
rect 800 155792 419200 157688
rect 800 155512 419120 155792
rect 800 154160 419200 155512
rect 880 153880 419200 154160
rect 800 152256 419200 153880
rect 800 151976 419120 152256
rect 800 150624 419200 151976
rect 880 150344 419200 150624
rect 800 148448 419200 150344
rect 800 148168 419120 148448
rect 800 147088 419200 148168
rect 880 146808 419200 147088
rect 800 144912 419200 146808
rect 800 144632 419120 144912
rect 800 143280 419200 144632
rect 880 143000 419200 143280
rect 800 141376 419200 143000
rect 800 141096 419120 141376
rect 800 139744 419200 141096
rect 880 139464 419200 139744
rect 800 137568 419200 139464
rect 800 137288 419120 137568
rect 800 135936 419200 137288
rect 880 135656 419200 135936
rect 800 134032 419200 135656
rect 800 133752 419120 134032
rect 800 132400 419200 133752
rect 880 132120 419200 132400
rect 800 130224 419200 132120
rect 800 129944 419120 130224
rect 800 128592 419200 129944
rect 880 128312 419200 128592
rect 800 126688 419200 128312
rect 800 126408 419120 126688
rect 800 125056 419200 126408
rect 880 124776 419200 125056
rect 800 122880 419200 124776
rect 800 122600 419120 122880
rect 800 121520 419200 122600
rect 880 121240 419200 121520
rect 800 119344 419200 121240
rect 800 119064 419120 119344
rect 800 117712 419200 119064
rect 880 117432 419200 117712
rect 800 115808 419200 117432
rect 800 115528 419120 115808
rect 800 114176 419200 115528
rect 880 113896 419200 114176
rect 800 112000 419200 113896
rect 800 111720 419120 112000
rect 800 110368 419200 111720
rect 880 110088 419200 110368
rect 800 108464 419200 110088
rect 800 108184 419120 108464
rect 800 106832 419200 108184
rect 880 106552 419200 106832
rect 800 104656 419200 106552
rect 800 104376 419120 104656
rect 800 103024 419200 104376
rect 880 102744 419200 103024
rect 800 101120 419200 102744
rect 800 100840 419120 101120
rect 800 99488 419200 100840
rect 880 99208 419200 99488
rect 800 97312 419200 99208
rect 800 97032 419120 97312
rect 800 95952 419200 97032
rect 880 95672 419200 95952
rect 800 93776 419200 95672
rect 800 93496 419120 93776
rect 800 92144 419200 93496
rect 880 91864 419200 92144
rect 800 90240 419200 91864
rect 800 89960 419120 90240
rect 800 88608 419200 89960
rect 880 88328 419200 88608
rect 800 86432 419200 88328
rect 800 86152 419120 86432
rect 800 84800 419200 86152
rect 880 84520 419200 84800
rect 800 82896 419200 84520
rect 800 82616 419120 82896
rect 800 81264 419200 82616
rect 880 80984 419200 81264
rect 800 79088 419200 80984
rect 800 78808 419120 79088
rect 800 77456 419200 78808
rect 880 77176 419200 77456
rect 800 75552 419200 77176
rect 800 75272 419120 75552
rect 800 73920 419200 75272
rect 880 73640 419200 73920
rect 800 71744 419200 73640
rect 800 71464 419120 71744
rect 800 70384 419200 71464
rect 880 70104 419200 70384
rect 800 68208 419200 70104
rect 800 67928 419120 68208
rect 800 66576 419200 67928
rect 880 66296 419200 66576
rect 800 64672 419200 66296
rect 800 64392 419120 64672
rect 800 63040 419200 64392
rect 880 62760 419200 63040
rect 800 60864 419200 62760
rect 800 60584 419120 60864
rect 800 59232 419200 60584
rect 880 58952 419200 59232
rect 800 57328 419200 58952
rect 800 57048 419120 57328
rect 800 55696 419200 57048
rect 880 55416 419200 55696
rect 800 53520 419200 55416
rect 800 53240 419120 53520
rect 800 51888 419200 53240
rect 880 51608 419200 51888
rect 800 49984 419200 51608
rect 800 49704 419120 49984
rect 800 48352 419200 49704
rect 880 48072 419200 48352
rect 800 46176 419200 48072
rect 800 45896 419120 46176
rect 800 44816 419200 45896
rect 880 44536 419200 44816
rect 800 42640 419200 44536
rect 800 42360 419120 42640
rect 800 41008 419200 42360
rect 880 40728 419200 41008
rect 800 39104 419200 40728
rect 800 38824 419120 39104
rect 800 37472 419200 38824
rect 880 37192 419200 37472
rect 800 35296 419200 37192
rect 800 35016 419120 35296
rect 800 33664 419200 35016
rect 880 33384 419200 33664
rect 800 31760 419200 33384
rect 800 31480 419120 31760
rect 800 30128 419200 31480
rect 880 29848 419200 30128
rect 800 27952 419200 29848
rect 800 27672 419120 27952
rect 800 26320 419200 27672
rect 880 26040 419200 26320
rect 800 24416 419200 26040
rect 800 24136 419120 24416
rect 800 22784 419200 24136
rect 880 22504 419200 22784
rect 800 20608 419200 22504
rect 800 20328 419120 20608
rect 800 19248 419200 20328
rect 880 18968 419200 19248
rect 800 17072 419200 18968
rect 800 16792 419120 17072
rect 800 15440 419200 16792
rect 880 15160 419200 15440
rect 800 13536 419200 15160
rect 800 13256 419120 13536
rect 800 11904 419200 13256
rect 880 11624 419200 11904
rect 800 9728 419200 11624
rect 800 9448 419120 9728
rect 800 8096 419200 9448
rect 880 7816 419200 8096
rect 800 6192 419200 7816
rect 800 5912 419120 6192
rect 800 4560 419200 5912
rect 880 4280 419200 4560
rect 800 2384 419200 4280
rect 800 2104 419120 2384
rect 800 851 419200 2104
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
<< obsm4 >>
rect 2451 2128 4128 497808
rect 4608 2128 19488 497808
rect 19968 2128 403888 497808
<< labels >>
rlabel metal2 s 21730 499200 21786 500000 6 io_in[0]
port 1 nsew default input
rlabel metal3 s 419200 203192 420000 203312 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 325514 499200 325570 500000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 329010 0 329066 800 6 io_in[12]
port 4 nsew default input
rlabel metal3 s 0 278264 800 278384 6 io_in[13]
port 5 nsew default input
rlabel metal3 s 0 102824 800 102944 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 46386 499200 46442 500000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 89442 0 89498 800 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 246578 499200 246634 500000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 393410 0 393466 800 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 177394 499200 177450 500000 6 io_in[19]
port 11 nsew default input
rlabel metal3 s 419200 130024 420000 130144 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 30194 0 30250 800 6 io_in[20]
port 13 nsew default input
rlabel metal3 s 0 212440 800 212560 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 82082 0 82138 800 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 318154 499200 318210 500000 6 io_in[23]
port 16 nsew default input
rlabel metal3 s 419200 13336 420000 13456 6 io_in[24]
port 17 nsew default input
rlabel metal3 s 0 161304 800 161424 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 47490 0 47546 800 6 io_in[26]
port 19 nsew default input
rlabel metal3 s 0 219784 800 219904 6 io_in[27]
port 20 nsew default input
rlabel metal3 s 419200 389512 420000 389632 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 96802 0 96858 800 6 io_in[29]
port 22 nsew default input
rlabel metal3 s 0 471928 800 472048 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 385866 0 385922 800 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 174818 499200 174874 500000 6 io_in[31]
port 25 nsew default input
rlabel metal3 s 0 62840 800 62960 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 194690 499200 194746 500000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 164882 499200 164938 500000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 203154 0 203210 800 6 io_in[35]
port 29 nsew default input
rlabel metal3 s 419200 400392 420000 400512 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 407026 499200 407082 500000 6 io_in[37]
port 31 nsew default input
rlabel metal3 s 419200 287240 420000 287360 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 163594 0 163650 800 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 64786 0 64842 800 6 io_in[5]
port 34 nsew default input
rlabel metal3 s 419200 484440 420000 484560 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 239034 499200 239090 500000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 36450 499200 36506 500000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 90914 499200 90970 500000 6 io_in[9]
port 38 nsew default input
rlabel metal3 s 419200 283432 420000 283552 6 io_oeb[0]
port 39 nsew default output
rlabel metal3 s 419200 440648 420000 440768 6 io_oeb[10]
port 40 nsew default output
rlabel metal3 s 419200 232296 420000 232416 6 io_oeb[11]
port 41 nsew default output
rlabel metal3 s 0 146888 800 147008 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 95698 499200 95754 500000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 79506 0 79562 800 6 io_oeb[14]
port 44 nsew default output
rlabel metal3 s 419200 68008 420000 68128 6 io_oeb[15]
port 45 nsew default output
rlabel metal3 s 0 121320 800 121440 6 io_oeb[16]
port 46 nsew default output
rlabel metal3 s 419200 224952 420000 225072 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 319258 0 319314 800 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 59818 0 59874 800 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 112994 499200 113050 500000 6 io_oeb[1]
port 50 nsew default output
rlabel metal3 s 419200 433304 420000 433424 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 300858 499200 300914 500000 6 io_oeb[21]
port 52 nsew default output
rlabel metal3 s 0 7896 800 8016 6 io_oeb[22]
port 53 nsew default output
rlabel metal3 s 0 55496 800 55616 6 io_oeb[23]
port 54 nsew default output
rlabel metal3 s 0 227128 800 227248 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 331586 0 331642 800 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 264794 0 264850 800 6 io_oeb[26]
port 57 nsew default output
rlabel metal3 s 419200 491784 420000 491904 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 379978 499200 380034 500000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 398194 0 398250 800 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 229282 499200 229338 500000 6 io_oeb[2]
port 61 nsew default output
rlabel metal3 s 0 216248 800 216368 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 240138 0 240194 800 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 34058 499200 34114 500000 6 io_oeb[32]
port 64 nsew default output
rlabel metal3 s 0 493688 800 493808 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 67178 0 67234 800 6 io_oeb[34]
port 66 nsew default output
rlabel metal3 s 0 245352 800 245472 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 14186 499200 14242 500000 6 io_oeb[36]
port 68 nsew default output
rlabel metal3 s 419200 301656 420000 301776 6 io_oeb[37]
port 69 nsew default output
rlabel metal3 s 0 124856 800 124976 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 399666 499200 399722 500000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 127898 499200 127954 500000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 419354 499200 419410 500000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 210514 0 210570 800 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 340418 499200 340474 500000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 86866 0 86922 800 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 103242 499200 103298 500000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 83370 499200 83426 500000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 109130 0 109186 800 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 306930 0 306986 800 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 321650 0 321706 800 6 io_out[13]
port 81 nsew default output
rlabel metal3 s 419200 272552 420000 272672 6 io_out[14]
port 82 nsew default output
rlabel metal3 s 419200 451528 420000 451648 6 io_out[15]
port 83 nsew default output
rlabel metal3 s 0 428136 800 428256 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 5354 0 5410 800 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 42522 0 42578 800 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 256330 499200 256386 500000 6 io_out[19]
port 87 nsew default output
rlabel metal3 s 0 110168 800 110288 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 247498 0 247554 800 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 49882 0 49938 800 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 104162 0 104218 800 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 358818 0 358874 800 6 io_out[23]
port 92 nsew default output
rlabel metal3 s 419200 312808 420000 312928 6 io_out[24]
port 93 nsew default output
rlabel metal3 s 0 369656 800 369776 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 84474 0 84530 800 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 105634 499200 105690 500000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 94410 0 94466 800 6 io_out[28]
port 97 nsew default output
rlabel metal3 s 0 249160 800 249280 6 io_out[29]
port 98 nsew default output
rlabel metal3 s 419200 469752 420000 469872 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 189722 499200 189778 500000 6 io_out[30]
port 100 nsew default output
rlabel metal3 s 419200 104456 420000 104576 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 266266 499200 266322 500000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 172426 499200 172482 500000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 71042 499200 71098 500000 6 io_out[34]
port 104 nsew default output
rlabel metal3 s 419200 126488 420000 126608 6 io_out[35]
port 105 nsew default output
rlabel metal3 s 0 296488 800 296608 6 io_out[36]
port 106 nsew default output
rlabel metal3 s 419200 462408 420000 462528 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 273626 499200 273682 500000 6 io_out[3]
port 108 nsew default output
rlabel metal3 s 419200 184968 420000 185088 6 io_out[4]
port 109 nsew default output
rlabel metal3 s 0 274728 800 274848 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 350354 499200 350410 500000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 111706 0 111762 800 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 245106 0 245162 800 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 48778 499200 48834 500000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 212906 0 212962 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal3 s 419200 93576 420000 93696 6 la_data_in[100]
port 116 nsew default input
rlabel metal3 s 419200 24216 420000 24336 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 130290 499200 130346 500000 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 372434 499200 372490 500000 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 281170 499200 281226 500000 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 343914 0 343970 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal3 s 0 208904 800 209024 6 la_data_in[106]
port 122 nsew default input
rlabel metal3 s 419200 155592 420000 155712 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 397274 499200 397330 500000 6 la_data_in[108]
port 124 nsew default input
rlabel metal3 s 0 179528 800 179648 6 la_data_in[109]
port 125 nsew default input
rlabel metal3 s 0 358504 800 358624 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 7930 0 7986 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal3 s 0 175992 800 176112 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 366178 0 366234 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 390834 0 390890 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 135258 499200 135314 500000 6 la_data_in[114]
port 131 nsew default input
rlabel metal3 s 0 186872 800 186992 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 313186 499200 313242 500000 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 282090 0 282146 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal3 s 0 497496 800 497616 6 la_data_in[11]
port 137 nsew default input
rlabel metal3 s 0 139544 800 139664 6 la_data_in[120]
port 138 nsew default input
rlabel metal3 s 0 402568 800 402688 6 la_data_in[121]
port 139 nsew default input
rlabel metal3 s 0 384072 800 384192 6 la_data_in[122]
port 140 nsew default input
rlabel metal3 s 419200 214072 420000 214192 6 la_data_in[123]
port 141 nsew default input
rlabel metal3 s 0 150424 800 150544 6 la_data_in[124]
port 142 nsew default input
rlabel metal3 s 419200 5992 420000 6112 6 la_data_in[125]
port 143 nsew default input
rlabel metal3 s 419200 385704 420000 385824 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 11794 499200 11850 500000 6 la_data_in[127]
port 145 nsew default input
rlabel metal3 s 419200 495320 420000 495440 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 162490 499200 162546 500000 6 la_data_in[15]
port 149 nsew default input
rlabel metal3 s 0 26120 800 26240 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 98274 499200 98330 500000 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 400770 0 400826 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 347778 499200 347834 500000 6 la_data_in[1]
port 154 nsew default input
rlabel metal3 s 419200 122680 420000 122800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 287058 0 287114 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal3 s 419200 455064 420000 455184 6 la_data_in[23]
port 158 nsew default input
rlabel metal3 s 419200 261672 420000 261792 6 la_data_in[24]
port 159 nsew default input
rlabel metal3 s 419200 334568 420000 334688 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 140226 499200 140282 500000 6 la_data_in[26]
port 161 nsew default input
rlabel metal3 s 0 303832 800 303952 6 la_data_in[27]
port 162 nsew default input
rlabel metal3 s 419200 119144 420000 119264 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 122930 499200 122986 500000 6 la_data_in[29]
port 164 nsew default input
rlabel metal3 s 0 340280 800 340400 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal3 s 419200 466216 420000 466336 6 la_data_in[31]
port 167 nsew default input
rlabel metal3 s 419200 217880 420000 218000 6 la_data_in[32]
port 168 nsew default input
rlabel metal3 s 0 70184 800 70304 6 la_data_in[33]
port 169 nsew default input
rlabel metal3 s 419200 378360 420000 378480 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 293498 499200 293554 500000 6 la_data_in[35]
port 171 nsew default input
rlabel metal3 s 0 398760 800 398880 6 la_data_in[36]
port 172 nsew default input
rlabel metal3 s 0 460776 800 460896 6 la_data_in[37]
port 173 nsew default input
rlabel metal3 s 419200 411272 420000 411392 6 la_data_in[38]
port 174 nsew default input
rlabel metal3 s 419200 356600 420000 356720 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal3 s 0 409640 800 409760 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 258906 499200 258962 500000 6 la_data_in[41]
port 178 nsew default input
rlabel metal3 s 0 51688 800 51808 6 la_data_in[42]
port 179 nsew default input
rlabel metal3 s 0 453704 800 453824 6 la_data_in[43]
port 180 nsew default input
rlabel metal3 s 419200 108264 420000 108384 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 263874 499200 263930 500000 6 la_data_in[45]
port 182 nsew default input
rlabel metal3 s 0 490152 800 490272 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 348882 0 348938 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 298466 499200 298522 500000 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 570 0 626 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal3 s 419200 367480 420000 367600 6 la_data_in[50]
port 188 nsew default input
rlabel metal3 s 0 190680 800 190800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal3 s 419200 254328 420000 254448 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 310794 499200 310850 500000 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 402242 499200 402298 500000 6 la_data_in[55]
port 193 nsew default input
rlabel metal3 s 419200 444184 420000 444304 6 la_data_in[56]
port 194 nsew default input
rlabel metal3 s 419200 458872 420000 458992 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 376114 0 376170 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 415490 0 415546 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 314290 0 314346 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal3 s 0 172456 800 172576 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 320546 499200 320602 500000 6 la_data_in[61]
port 200 nsew default input
rlabel metal3 s 419200 38904 420000 39024 6 la_data_in[62]
port 201 nsew default input
rlabel metal3 s 0 307368 800 307488 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 308218 499200 308274 500000 6 la_data_in[64]
port 203 nsew default input
rlabel metal3 s 0 81064 800 81184 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 279698 0 279754 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal3 s 419200 206728 420000 206848 6 la_data_in[67]
port 206 nsew default input
rlabel metal3 s 0 464584 800 464704 6 la_data_in[68]
port 207 nsew default input
rlabel metal3 s 0 377000 800 377120 6 la_data_in[69]
port 208 nsew default input
rlabel metal3 s 419200 477096 420000 477216 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 261298 499200 261354 500000 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 351274 0 351330 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal3 s 0 238008 800 238128 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 26514 499200 26570 500000 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 78402 499200 78458 500000 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal3 s 419200 177624 420000 177744 6 la_data_in[76]
port 216 nsew default input
rlabel metal3 s 419200 64472 420000 64592 6 la_data_in[77]
port 217 nsew default input
rlabel metal3 s 0 168648 800 168768 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 388442 0 388498 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal3 s 419200 298120 420000 298240 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 346306 0 346362 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal3 s 419200 9528 420000 9648 6 la_data_in[81]
port 222 nsew default input
rlabel metal3 s 419200 447992 420000 448112 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 192114 499200 192170 500000 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 20258 0 20314 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal3 s 0 431672 800 431792 6 la_data_in[86]
port 227 nsew default input
rlabel metal3 s 0 157768 800 157888 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 341522 0 341578 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 100666 499200 100722 500000 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 410706 0 410762 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 155130 499200 155186 500000 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 360106 499200 360162 500000 6 la_data_in[91]
port 233 nsew default input
rlabel metal3 s 0 143080 800 143200 6 la_data_in[92]
port 234 nsew default input
rlabel metal3 s 0 270920 800 271040 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 173346 0 173402 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 76010 499200 76066 500000 6 la_data_in[95]
port 237 nsew default input
rlabel metal3 s 419200 115608 420000 115728 6 la_data_in[96]
port 238 nsew default input
rlabel metal3 s 0 395224 800 395344 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 301962 0 302018 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal3 s 419200 309000 420000 309120 6 la_data_in[99]
port 241 nsew default input
rlabel metal3 s 0 289144 800 289264 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 207938 0 207994 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 395802 0 395858 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal3 s 419200 31560 420000 31680 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 22650 0 22706 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal3 s 419200 243448 420000 243568 6 la_data_out[104]
port 248 nsew default output
rlabel metal3 s 0 99288 800 99408 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal3 s 0 435208 800 435328 6 la_data_out[107]
port 251 nsew default output
rlabel metal3 s 0 420792 800 420912 6 la_data_out[108]
port 252 nsew default output
rlabel metal3 s 0 406104 800 406224 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 389730 499200 389786 500000 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 225234 0 225290 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 4434 499200 4490 500000 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal3 s 0 311176 800 311296 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 370042 499200 370098 500000 6 la_data_out[114]
port 259 nsew default output
rlabel metal3 s 419200 473560 420000 473680 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 299386 0 299442 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal3 s 419200 181160 420000 181280 6 la_data_out[117]
port 262 nsew default output
rlabel metal3 s 419200 239640 420000 239760 6 la_data_out[118]
port 263 nsew default output
rlabel metal3 s 0 66376 800 66496 6 la_data_out[119]
port 264 nsew default output
rlabel metal3 s 0 344088 800 344208 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 160098 499200 160154 500000 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 56322 499200 56378 500000 6 la_data_out[121]
port 267 nsew default output
rlabel metal3 s 0 153960 800 154080 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 288530 499200 288586 500000 6 la_data_out[124]
port 270 nsew default output
rlabel metal3 s 419200 111800 420000 111920 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 215482 0 215538 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 368570 0 368626 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 241610 499200 241666 500000 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 278594 499200 278650 500000 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 170954 0 171010 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 403162 0 403218 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 110602 499200 110658 500000 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 316682 0 316738 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal3 s 419200 374824 420000 374944 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 209410 499200 209466 500000 6 la_data_out[1]
port 282 nsew default output
rlabel metal3 s 419200 418616 420000 418736 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 115570 499200 115626 500000 6 la_data_out[21]
port 284 nsew default output
rlabel metal3 s 0 329400 800 329520 6 la_data_out[22]
port 285 nsew default output
rlabel metal3 s 419200 162936 420000 163056 6 la_data_out[23]
port 286 nsew default output
rlabel metal3 s 0 241816 800 241936 6 la_data_out[24]
port 287 nsew default output
rlabel metal3 s 419200 436840 420000 436960 6 la_data_out[25]
port 288 nsew default output
rlabel metal3 s 419200 290776 420000 290896 6 la_data_out[26]
port 289 nsew default output
rlabel metal3 s 0 332936 800 333056 6 la_data_out[27]
port 290 nsew default output
rlabel metal3 s 419200 199384 420000 199504 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal3 s 419200 195848 420000 195968 6 la_data_out[2]
port 293 nsew default output
rlabel metal3 s 0 336744 800 336864 6 la_data_out[30]
port 294 nsew default output
rlabel metal3 s 0 33464 800 33584 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 315762 499200 315818 500000 6 la_data_out[32]
port 296 nsew default output
rlabel metal3 s 419200 20408 420000 20528 6 la_data_out[33]
port 297 nsew default output
rlabel metal3 s 419200 133832 420000 133952 6 la_data_out[34]
port 298 nsew default output
rlabel metal3 s 419200 82696 420000 82816 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 222842 0 222898 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal3 s 419200 349256 420000 349376 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 43810 499200 43866 500000 6 la_data_out[38]
port 302 nsew default output
rlabel metal3 s 0 486344 800 486464 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 330482 499200 330538 500000 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 303250 499200 303306 500000 6 la_data_out[41]
port 306 nsew default output
rlabel metal3 s 419200 294584 420000 294704 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 145194 499200 145250 500000 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal3 s 0 205096 800 205216 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 211986 499200 212042 500000 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 414570 499200 414626 500000 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 61106 499200 61162 500000 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 220450 0 220506 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal3 s 0 77256 800 77376 6 la_data_out[4]
port 315 nsew default output
rlabel metal3 s 0 201560 800 201680 6 la_data_out[50]
port 316 nsew default output
rlabel metal3 s 0 446360 800 446480 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal3 s 419200 407736 420000 407856 6 la_data_out[53]
port 319 nsew default output
rlabel metal3 s 0 113976 800 114096 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 352746 499200 352802 500000 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 271234 499200 271290 500000 6 la_data_out[56]
port 322 nsew default output
rlabel metal3 s 419200 170280 420000 170400 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 198186 0 198242 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal3 s 0 117512 800 117632 6 la_data_out[59]
port 325 nsew default output
rlabel metal3 s 419200 382168 420000 382288 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 408130 0 408186 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 251362 499200 251418 500000 6 la_data_out[61]
port 328 nsew default output
rlabel metal3 s 419200 250520 420000 250640 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 323122 499200 323178 500000 6 la_data_out[64]
port 331 nsew default output
rlabel metal3 s 0 40808 800 40928 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 289634 0 289690 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 296994 0 297050 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 336554 0 336610 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 202050 499200 202106 500000 6 la_data_out[6]
port 337 nsew default output
rlabel metal3 s 0 4360 800 4480 6 la_data_out[70]
port 338 nsew default output
rlabel metal3 s 419200 257864 420000 257984 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 378506 0 378562 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal3 s 419200 42440 420000 42560 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 405738 0 405794 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 137834 499200 137890 500000 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 404634 499200 404690 500000 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 183282 0 183338 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 353850 0 353906 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 17682 0 17738 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal3 s 419200 141176 420000 141296 6 la_data_out[7]
port 348 nsew default output
rlabel metal3 s 0 91944 800 92064 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 272338 0 272394 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 337842 499200 337898 500000 6 la_data_out[83]
port 352 nsew default output
rlabel metal3 s 0 263576 800 263696 6 la_data_out[84]
port 353 nsew default output
rlabel metal3 s 419200 269016 420000 269136 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 277122 0 277178 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal3 s 0 387880 800 388000 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 309322 0 309378 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal3 s 0 22584 800 22704 6 la_data_out[89]
port 358 nsew default output
rlabel metal3 s 0 457240 800 457360 6 la_data_out[8]
port 359 nsew default output
rlabel metal3 s 0 479272 800 479392 6 la_data_out[90]
port 360 nsew default output
rlabel metal3 s 0 84600 800 84720 6 la_data_out[91]
port 361 nsew default output
rlabel metal3 s 419200 236104 420000 236224 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 147586 499200 147642 500000 6 la_data_out[93]
port 363 nsew default output
rlabel metal3 s 419200 228760 420000 228880 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 413098 0 413154 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 58714 499200 58770 500000 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 12898 0 12954 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 392306 499200 392362 500000 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 377402 499200 377458 500000 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 6826 499200 6882 500000 6 la_data_out[9]
port 370 nsew default output
rlabel metal3 s 0 380536 800 380656 6 la_oen[0]
port 371 nsew default input
rlabel metal3 s 419200 371288 420000 371408 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 207018 499200 207074 500000 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 153658 0 153714 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 165986 0 166042 800 6 la_oen[103]
port 375 nsew default input
rlabel metal3 s 419200 279896 420000 280016 6 la_oen[104]
port 376 nsew default input
rlabel metal3 s 419200 210536 420000 210656 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 15290 0 15346 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 190642 0 190698 800 6 la_oen[107]
port 379 nsew default input
rlabel metal3 s 419200 393048 420000 393168 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 184754 499200 184810 500000 6 la_oen[109]
port 381 nsew default input
rlabel metal3 s 419200 320152 420000 320272 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 187146 499200 187202 500000 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 295890 499200 295946 500000 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 292026 0 292082 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 200578 0 200634 800 6 la_oen[113]
port 386 nsew default input
rlabel metal3 s 0 449896 800 450016 6 la_oen[114]
port 387 nsew default input
rlabel metal3 s 0 59032 800 59152 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 132866 499200 132922 500000 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 226706 499200 226762 500000 6 la_oen[117]
port 390 nsew default input
rlabel metal3 s 419200 144712 420000 144832 6 la_oen[118]
port 391 nsew default input
rlabel metal3 s 0 183336 800 183456 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 108210 499200 108266 500000 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 283562 499200 283618 500000 6 la_oen[120]
port 394 nsew default input
rlabel metal3 s 0 88408 800 88528 6 la_oen[121]
port 395 nsew default input
rlabel metal3 s 419200 49784 420000 49904 6 la_oen[122]
port 396 nsew default input
rlabel metal3 s 0 11704 800 11824 6 la_oen[123]
port 397 nsew default input
rlabel metal3 s 419200 2184 420000 2304 6 la_oen[124]
port 398 nsew default input
rlabel metal3 s 419200 480632 420000 480752 6 la_oen[125]
port 399 nsew default input
rlabel metal3 s 419200 86232 420000 86352 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 62210 0 62266 800 6 la_oen[127]
port 401 nsew default input
rlabel metal3 s 0 198024 800 198144 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 342810 499200 342866 500000 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 361210 0 361266 800 6 la_oen[14]
port 404 nsew default input
rlabel metal3 s 419200 148248 420000 148368 6 la_oen[15]
port 405 nsew default input
rlabel metal3 s 419200 166744 420000 166864 6 la_oen[16]
port 406 nsew default input
rlabel metal3 s 419200 363944 420000 364064 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 244002 499200 244058 500000 6 la_oen[18]
port 408 nsew default input
rlabel metal3 s 0 95752 800 95872 6 la_oen[19]
port 409 nsew default input
rlabel metal3 s 0 292952 800 293072 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 193218 0 193274 800 6 la_oen[20]
port 411 nsew default input
rlabel metal3 s 419200 265208 420000 265328 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 236642 499200 236698 500000 6 la_oen[22]
port 413 nsew default input
rlabel metal3 s 419200 100920 420000 101040 6 la_oen[23]
port 414 nsew default input
rlabel metal3 s 0 373192 800 373312 6 la_oen[24]
port 415 nsew default input
rlabel metal3 s 419200 345720 420000 345840 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 188250 0 188306 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 124034 0 124090 800 6 la_oen[27]
port 418 nsew default input
rlabel metal3 s 419200 35096 420000 35216 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 227810 0 227866 800 6 la_oen[29]
port 420 nsew default input
rlabel metal3 s 419200 75352 420000 75472 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 230202 0 230258 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 304354 0 304410 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 2962 0 3018 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 380898 0 380954 800 6 la_oen[33]
port 425 nsew default input
rlabel metal3 s 419200 16872 420000 16992 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 88338 499200 88394 500000 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 53746 499200 53802 500000 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 9218 499200 9274 500000 6 la_oen[37]
port 429 nsew default input
rlabel metal3 s 0 354968 800 355088 6 la_oen[38]
port 430 nsew default input
rlabel metal3 s 0 256232 800 256352 6 la_oen[39]
port 431 nsew default input
rlabel metal3 s 419200 352792 420000 352912 6 la_oen[3]
port 432 nsew default input
rlabel metal3 s 419200 422424 420000 422544 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 367650 499200 367706 500000 6 la_oen[41]
port 434 nsew default input
rlabel metal3 s 419200 360136 420000 360256 6 la_oen[42]
port 435 nsew default input
rlabel metal3 s 0 475464 800 475584 6 la_oen[43]
port 436 nsew default input
rlabel metal3 s 419200 57128 420000 57248 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 355138 499200 355194 500000 6 la_oen[45]
port 438 nsew default input
rlabel metal3 s 419200 331032 420000 331152 6 la_oen[46]
port 439 nsew default input
rlabel metal3 s 419200 173816 420000 173936 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 219346 499200 219402 500000 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 248970 499200 249026 500000 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 150162 499200 150218 500000 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 345386 499200 345442 500000 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 205546 0 205602 800 6 la_oen[51]
port 445 nsew default input
rlabel metal3 s 419200 305464 420000 305584 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 73618 499200 73674 500000 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 409602 499200 409658 500000 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 66074 499200 66130 500000 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 305826 499200 305882 500000 6 la_oen[56]
port 450 nsew default input
rlabel metal3 s 0 413448 800 413568 6 la_oen[57]
port 451 nsew default input
rlabel metal3 s 0 223592 800 223712 6 la_oen[58]
port 452 nsew default input
rlabel metal3 s 419200 403928 420000 404048 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 80978 499200 81034 500000 6 la_oen[5]
port 454 nsew default input
rlabel metal3 s 0 416984 800 417104 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 199474 499200 199530 500000 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 237746 0 237802 800 6 la_oen[62]
port 457 nsew default input
rlabel metal3 s 419200 192312 420000 192432 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 333978 0 334034 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 101770 0 101826 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 375010 499200 375066 500000 6 la_oen[66]
port 461 nsew default input
rlabel metal3 s 0 314712 800 314832 6 la_oen[67]
port 462 nsew default input
rlabel metal3 s 0 285608 800 285728 6 la_oen[68]
port 463 nsew default input
rlabel metal3 s 419200 429496 420000 429616 6 la_oen[69]
port 464 nsew default input
rlabel metal3 s 0 135736 800 135856 6 la_oen[6]
port 465 nsew default input
rlabel metal3 s 0 424328 800 424448 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 290922 499200 290978 500000 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 362682 499200 362738 500000 6 la_oen[72]
port 468 nsew default input
rlabel metal3 s 0 442552 800 442672 6 la_oen[73]
port 469 nsew default input
rlabel metal3 s 419200 152056 420000 152176 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 129002 0 129058 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 185858 0 185914 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 93306 499200 93362 500000 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 216770 499200 216826 500000 6 la_oen[78]
port 474 nsew default input
rlabel metal3 s 419200 327224 420000 327344 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 63682 499200 63738 500000 6 la_oen[7]
port 476 nsew default input
rlabel metal3 s 0 439016 800 439136 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 16762 499200 16818 500000 6 la_oen[81]
port 478 nsew default input
rlabel metal3 s 419200 97112 420000 97232 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 253938 499200 253994 500000 6 la_oen[83]
port 480 nsew default input
rlabel metal3 s 0 106632 800 106752 6 la_oen[84]
port 481 nsew default input
rlabel metal3 s 419200 159400 420000 159520 6 la_oen[85]
port 482 nsew default input
rlabel metal3 s 419200 396856 420000 396976 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 411994 499200 412050 500000 6 la_oen[87]
port 484 nsew default input
rlabel metal3 s 419200 60664 420000 60784 6 la_oen[88]
port 485 nsew default input
rlabel metal3 s 0 347624 800 347744 6 la_oen[89]
port 486 nsew default input
rlabel metal3 s 419200 45976 420000 46096 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 167458 499200 167514 500000 6 la_oen[90]
port 488 nsew default input
rlabel metal3 s 419200 78888 420000 79008 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 91834 0 91890 800 6 la_oen[92]
port 490 nsew default input
rlabel metal3 s 0 234472 800 234592 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 333058 499200 333114 500000 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 373538 0 373594 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 276202 499200 276258 500000 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 363602 0 363658 800 6 la_oen[97]
port 495 nsew default input
rlabel metal3 s 419200 27752 420000 27872 6 la_oen[98]
port 496 nsew default input
rlabel metal3 s 0 322056 800 322176 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 294418 0 294474 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 161018 0 161074 800 6 vccd1
port 499 nsew default bidirectional
rlabel metal3 s 0 482808 800 482928 6 vccd2
port 500 nsew default bidirectional
rlabel metal2 s 169850 499200 169906 500000 6 vdda1
port 501 nsew default bidirectional
rlabel metal3 s 0 252696 800 252816 6 vdda2
port 502 nsew default bidirectional
rlabel metal3 s 419200 425960 420000 426080 6 vssa1
port 503 nsew default bidirectional
rlabel metal2 s 250074 0 250130 800 6 vssa2
port 504 nsew default bidirectional
rlabel metal2 s 99378 0 99434 800 6 vssd1
port 505 nsew default bidirectional
rlabel metal2 s 267370 0 267426 800 6 vssd2
port 506 nsew default bidirectional
rlabel metal2 s 39026 499200 39082 500000 6 wb_clk_i
port 507 nsew default input
rlabel metal2 s 1858 499200 1914 500000 6 wb_rst_i
port 508 nsew default input
rlabel metal2 s 224314 499200 224370 500000 6 wbs_ack_o
port 509 nsew default output
rlabel metal2 s 24122 499200 24178 500000 6 wbs_adr_i[0]
port 510 nsew default input
rlabel metal2 s 382370 499200 382426 500000 6 wbs_adr_i[10]
port 511 nsew default input
rlabel metal2 s 285954 499200 286010 500000 6 wbs_adr_i[11]
port 512 nsew default input
rlabel metal3 s 419200 137368 420000 137488 6 wbs_adr_i[12]
port 513 nsew default input
rlabel metal2 s 151266 0 151322 800 6 wbs_adr_i[13]
port 514 nsew default input
rlabel metal3 s 0 230664 800 230784 6 wbs_adr_i[14]
port 515 nsew default input
rlabel metal3 s 0 281800 800 281920 6 wbs_adr_i[15]
port 516 nsew default input
rlabel metal3 s 0 194216 800 194336 6 wbs_adr_i[16]
port 517 nsew default input
rlabel metal2 s 204442 499200 204498 500000 6 wbs_adr_i[17]
port 518 nsew default input
rlabel metal2 s 394698 499200 394754 500000 6 wbs_adr_i[18]
port 519 nsew default input
rlabel metal3 s 0 300296 800 300416 6 wbs_adr_i[19]
port 520 nsew default input
rlabel metal3 s 0 44616 800 44736 6 wbs_adr_i[1]
port 521 nsew default input
rlabel metal3 s 419200 53320 420000 53440 6 wbs_adr_i[20]
port 522 nsew default input
rlabel metal3 s 419200 341912 420000 342032 6 wbs_adr_i[21]
port 523 nsew default input
rlabel metal2 s 197082 499200 197138 500000 6 wbs_adr_i[22]
port 524 nsew default input
rlabel metal2 s 120538 499200 120594 500000 6 wbs_adr_i[23]
port 525 nsew default input
rlabel metal3 s 419200 338376 420000 338496 6 wbs_adr_i[24]
port 526 nsew default input
rlabel metal2 s 311714 0 311770 800 6 wbs_adr_i[25]
port 527 nsew default input
rlabel metal2 s 126426 0 126482 800 6 wbs_adr_i[26]
port 528 nsew default input
rlabel metal3 s 0 37272 800 37392 6 wbs_adr_i[27]
port 529 nsew default input
rlabel metal2 s 156050 0 156106 800 6 wbs_adr_i[28]
port 530 nsew default input
rlabel metal2 s 214378 499200 214434 500000 6 wbs_adr_i[29]
port 531 nsew default input
rlabel metal2 s 356242 0 356298 800 6 wbs_adr_i[2]
port 532 nsew default input
rlabel metal3 s 419200 188504 420000 188624 6 wbs_adr_i[30]
port 533 nsew default input
rlabel metal3 s 0 73720 800 73840 6 wbs_adr_i[31]
port 534 nsew default input
rlabel metal2 s 274730 0 274786 800 6 wbs_adr_i[3]
port 535 nsew default input
rlabel metal2 s 182178 499200 182234 500000 6 wbs_adr_i[4]
port 536 nsew default input
rlabel metal2 s 232778 0 232834 800 6 wbs_adr_i[5]
port 537 nsew default input
rlabel metal2 s 269762 0 269818 800 6 wbs_adr_i[6]
port 538 nsew default input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[7]
port 539 nsew default input
rlabel metal3 s 0 132200 800 132320 6 wbs_adr_i[8]
port 540 nsew default input
rlabel metal2 s 326618 0 326674 800 6 wbs_adr_i[9]
port 541 nsew default input
rlabel metal2 s 51354 499200 51410 500000 6 wbs_cyc_i
port 542 nsew default input
rlabel metal2 s 195610 0 195666 800 6 wbs_dat_i[0]
port 543 nsew default input
rlabel metal3 s 0 267384 800 267504 6 wbs_dat_i[10]
port 544 nsew default input
rlabel metal2 s 387338 499200 387394 500000 6 wbs_dat_i[11]
port 545 nsew default input
rlabel metal3 s 0 29928 800 30048 6 wbs_dat_i[12]
port 546 nsew default input
rlabel metal2 s 384946 499200 385002 500000 6 wbs_dat_i[13]
port 547 nsew default input
rlabel metal3 s 419200 487976 420000 488096 6 wbs_dat_i[14]
port 548 nsew default input
rlabel metal2 s 335450 499200 335506 500000 6 wbs_dat_i[15]
port 549 nsew default input
rlabel metal2 s 158626 0 158682 800 6 wbs_dat_i[16]
port 550 nsew default input
rlabel metal2 s 41418 499200 41474 500000 6 wbs_dat_i[17]
port 551 nsew default input
rlabel metal3 s 0 391416 800 391536 6 wbs_dat_i[18]
port 552 nsew default input
rlabel metal2 s 231674 499200 231730 500000 6 wbs_dat_i[19]
port 553 nsew default input
rlabel metal3 s 419200 316344 420000 316464 6 wbs_dat_i[1]
port 554 nsew default input
rlabel metal3 s 419200 323688 420000 323808 6 wbs_dat_i[20]
port 555 nsew default input
rlabel metal2 s 29090 499200 29146 500000 6 wbs_dat_i[21]
port 556 nsew default input
rlabel metal2 s 131394 0 131450 800 6 wbs_dat_i[22]
port 557 nsew default input
rlabel metal3 s 419200 71544 420000 71664 6 wbs_dat_i[23]
port 558 nsew default input
rlabel metal3 s 419200 90040 420000 90160 6 wbs_dat_i[24]
port 559 nsew default input
rlabel metal2 s 338946 0 339002 800 6 wbs_dat_i[25]
port 560 nsew default input
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_i[26]
port 561 nsew default input
rlabel metal3 s 419200 276088 420000 276208 6 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 255042 0 255098 800 6 wbs_dat_i[28]
port 563 nsew default input
rlabel metal2 s 178314 0 178370 800 6 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 257434 0 257490 800 6 wbs_dat_i[2]
port 565 nsew default input
rlabel metal3 s 0 365848 800 365968 6 wbs_dat_i[30]
port 566 nsew default input
rlabel metal2 s 371146 0 371202 800 6 wbs_dat_i[31]
port 567 nsew default input
rlabel metal2 s 234066 499200 234122 500000 6 wbs_dat_i[3]
port 568 nsew default input
rlabel metal2 s 116674 0 116730 800 6 wbs_dat_i[4]
port 569 nsew default input
rlabel metal2 s 157522 499200 157578 500000 6 wbs_dat_i[5]
port 570 nsew default input
rlabel metal2 s 357714 499200 357770 500000 6 wbs_dat_i[6]
port 571 nsew default input
rlabel metal3 s 0 318520 800 318640 6 wbs_dat_i[7]
port 572 nsew default input
rlabel metal2 s 179786 499200 179842 500000 6 wbs_dat_i[8]
port 573 nsew default input
rlabel metal2 s 383474 0 383530 800 6 wbs_dat_i[9]
port 574 nsew default input
rlabel metal3 s 0 260040 800 260160 6 wbs_dat_o[0]
port 575 nsew default output
rlabel metal2 s 418066 0 418122 800 6 wbs_dat_o[10]
port 576 nsew default output
rlabel metal2 s 217874 0 217930 800 6 wbs_dat_o[11]
port 577 nsew default output
rlabel metal3 s 0 165112 800 165232 6 wbs_dat_o[12]
port 578 nsew default output
rlabel metal2 s 31482 499200 31538 500000 6 wbs_dat_o[13]
port 579 nsew default output
rlabel metal2 s 416962 499200 417018 500000 6 wbs_dat_o[14]
port 580 nsew default output
rlabel metal2 s 242530 0 242586 800 6 wbs_dat_o[15]
port 581 nsew default output
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_o[16]
port 582 nsew default output
rlabel metal2 s 365074 499200 365130 500000 6 wbs_dat_o[17]
port 583 nsew default output
rlabel metal2 s 85946 499200 86002 500000 6 wbs_dat_o[18]
port 584 nsew default output
rlabel metal2 s 142802 499200 142858 500000 6 wbs_dat_o[19]
port 585 nsew default output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[1]
port 586 nsew default output
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_o[20]
port 587 nsew default output
rlabel metal2 s 119066 0 119122 800 6 wbs_dat_o[21]
port 588 nsew default output
rlabel metal2 s 284666 0 284722 800 6 wbs_dat_o[22]
port 589 nsew default output
rlabel metal2 s 324226 0 324282 800 6 wbs_dat_o[23]
port 590 nsew default output
rlabel metal3 s 0 351432 800 351552 6 wbs_dat_o[24]
port 591 nsew default output
rlabel metal2 s 117962 499200 118018 500000 6 wbs_dat_o[25]
port 592 nsew default output
rlabel metal3 s 0 15240 800 15360 6 wbs_dat_o[26]
port 593 nsew default output
rlabel metal3 s 0 362312 800 362432 6 wbs_dat_o[27]
port 594 nsew default output
rlabel metal3 s 419200 415080 420000 415200 6 wbs_dat_o[28]
port 595 nsew default output
rlabel metal2 s 152554 499200 152610 500000 6 wbs_dat_o[29]
port 596 nsew default output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[2]
port 597 nsew default output
rlabel metal3 s 0 128392 800 128512 6 wbs_dat_o[30]
port 598 nsew default output
rlabel metal2 s 19154 499200 19210 500000 6 wbs_dat_o[31]
port 599 nsew default output
rlabel metal2 s 125506 499200 125562 500000 6 wbs_dat_o[3]
port 600 nsew default output
rlabel metal2 s 328090 499200 328146 500000 6 wbs_dat_o[4]
port 601 nsew default output
rlabel metal2 s 268658 499200 268714 500000 6 wbs_dat_o[5]
port 602 nsew default output
rlabel metal2 s 68650 499200 68706 500000 6 wbs_dat_o[6]
port 603 nsew default output
rlabel metal2 s 259826 0 259882 800 6 wbs_dat_o[7]
port 604 nsew default output
rlabel metal2 s 235170 0 235226 800 6 wbs_dat_o[8]
port 605 nsew default output
rlabel metal3 s 0 468120 800 468240 6 wbs_dat_o[9]
port 606 nsew default output
rlabel metal3 s 0 325864 800 325984 6 wbs_sel_i[0]
port 607 nsew default input
rlabel metal3 s 419200 246984 420000 247104 6 wbs_sel_i[1]
port 608 nsew default input
rlabel metal2 s 77114 0 77170 800 6 wbs_sel_i[2]
port 609 nsew default input
rlabel metal2 s 221738 499200 221794 500000 6 wbs_sel_i[3]
port 610 nsew default input
rlabel metal3 s 419200 221416 420000 221536 6 wbs_stb_i
port 611 nsew default input
rlabel metal3 s 0 48152 800 48272 6 wbs_we_i
port 612 nsew default input
rlabel metal4 s 4208 2128 4528 497808 6 VPWR
port 613 nsew power input
rlabel metal4 s 19568 2128 19888 497808 6 VGND
port 614 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 420000 500000
string LEFview TRUE
<< end >>
